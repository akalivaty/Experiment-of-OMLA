

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  INV_X1 U558 ( .A(n600), .ZN(n653) );
  AND2_X2 U559 ( .A1(n527), .A2(G2105), .ZN(n869) );
  XNOR2_X1 U560 ( .A(n599), .B(KEYINPUT26), .ZN(n601) );
  NOR2_X1 U561 ( .A1(n679), .A2(G1966), .ZN(n671) );
  XNOR2_X1 U562 ( .A(n666), .B(KEYINPUT31), .ZN(n667) );
  NAND2_X1 U563 ( .A1(n597), .A2(G160), .ZN(n600) );
  NOR2_X1 U564 ( .A1(n533), .A2(n532), .ZN(G164) );
  NAND2_X1 U565 ( .A1(G40), .A2(G160), .ZN(n522) );
  NOR2_X4 U566 ( .A1(n527), .A2(G2105), .ZN(n874) );
  XNOR2_X2 U567 ( .A(KEYINPUT65), .B(G2104), .ZN(n527) );
  AND2_X1 U568 ( .A1(n723), .A2(n722), .ZN(n523) );
  XNOR2_X1 U569 ( .A(KEYINPUT94), .B(KEYINPUT30), .ZN(n660) );
  BUF_X1 U570 ( .A(n600), .Z(n680) );
  INV_X1 U571 ( .A(KEYINPUT98), .ZN(n695) );
  NAND2_X1 U572 ( .A1(n874), .A2(G101), .ZN(n538) );
  INV_X1 U573 ( .A(n529), .ZN(n877) );
  NOR2_X1 U574 ( .A1(G651), .A2(n580), .ZN(n791) );
  AND2_X1 U575 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U576 ( .A1(G126), .A2(n869), .ZN(n525) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n870) );
  NAND2_X1 U578 ( .A1(G114), .A2(n870), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U580 ( .A(KEYINPUT86), .B(n526), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n874), .A2(G102), .ZN(n531) );
  XOR2_X1 U582 ( .A(KEYINPUT17), .B(n528), .Z(n534) );
  INV_X1 U583 ( .A(n534), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n877), .A2(G138), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U586 ( .A1(G137), .A2(n534), .ZN(n536) );
  NAND2_X1 U587 ( .A1(G113), .A2(n870), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U589 ( .A(n537), .B(KEYINPUT66), .ZN(n540) );
  XNOR2_X1 U590 ( .A(KEYINPUT23), .B(n538), .ZN(n539) );
  NOR2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U592 ( .A1(n869), .A2(G125), .ZN(n541) );
  XNOR2_X2 U593 ( .A(KEYINPUT64), .B(n543), .ZN(G160) );
  INV_X1 U594 ( .A(G651), .ZN(n547) );
  NOR2_X1 U595 ( .A1(G543), .A2(n547), .ZN(n544) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n544), .Z(n790) );
  NAND2_X1 U597 ( .A1(G64), .A2(n790), .ZN(n546) );
  XOR2_X1 U598 ( .A(KEYINPUT0), .B(G543), .Z(n580) );
  NAND2_X1 U599 ( .A1(G52), .A2(n791), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n553) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n794) );
  NAND2_X1 U602 ( .A1(G90), .A2(n794), .ZN(n549) );
  NOR2_X1 U603 ( .A1(n580), .A2(n547), .ZN(n795) );
  NAND2_X1 U604 ( .A1(G77), .A2(n795), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U606 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  XNOR2_X1 U607 ( .A(KEYINPUT67), .B(n551), .ZN(n552) );
  NOR2_X1 U608 ( .A1(n553), .A2(n552), .ZN(G171) );
  INV_X1 U609 ( .A(G171), .ZN(G301) );
  NAND2_X1 U610 ( .A1(G63), .A2(n790), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G51), .A2(n791), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n557) );
  XOR2_X1 U613 ( .A(KEYINPUT6), .B(KEYINPUT75), .Z(n556) );
  XNOR2_X1 U614 ( .A(n557), .B(n556), .ZN(n565) );
  XNOR2_X1 U615 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n563) );
  NAND2_X1 U616 ( .A1(n794), .A2(G89), .ZN(n558) );
  XNOR2_X1 U617 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G76), .A2(n795), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT5), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n563), .B(n562), .ZN(n564) );
  NOR2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U623 ( .A(KEYINPUT7), .B(n566), .Z(n567) );
  XNOR2_X1 U624 ( .A(KEYINPUT76), .B(n567), .ZN(G168) );
  XOR2_X1 U625 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U626 ( .A1(G75), .A2(n795), .ZN(n569) );
  NAND2_X1 U627 ( .A1(G62), .A2(n790), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n794), .A2(G88), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT82), .B(n570), .Z(n571) );
  NOR2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n791), .A2(G50), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n574), .A2(n573), .ZN(G303) );
  NAND2_X1 U634 ( .A1(n791), .A2(G49), .ZN(n575) );
  XOR2_X1 U635 ( .A(KEYINPUT79), .B(n575), .Z(n577) );
  NAND2_X1 U636 ( .A1(G651), .A2(G74), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U638 ( .A(KEYINPUT80), .B(n578), .ZN(n579) );
  NOR2_X1 U639 ( .A1(n790), .A2(n579), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n580), .A2(G87), .ZN(n581) );
  NAND2_X1 U641 ( .A1(n582), .A2(n581), .ZN(G288) );
  NAND2_X1 U642 ( .A1(G86), .A2(n794), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G61), .A2(n790), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U645 ( .A1(G73), .A2(n795), .ZN(n585) );
  XNOR2_X1 U646 ( .A(n585), .B(KEYINPUT81), .ZN(n586) );
  XNOR2_X1 U647 ( .A(n586), .B(KEYINPUT2), .ZN(n587) );
  NOR2_X1 U648 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U649 ( .A1(n791), .A2(G48), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n590), .A2(n589), .ZN(G305) );
  INV_X1 U651 ( .A(G303), .ZN(G166) );
  NAND2_X1 U652 ( .A1(G85), .A2(n794), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G72), .A2(n795), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U655 ( .A1(G60), .A2(n790), .ZN(n594) );
  NAND2_X1 U656 ( .A1(G47), .A2(n791), .ZN(n593) );
  NAND2_X1 U657 ( .A1(n594), .A2(n593), .ZN(n595) );
  OR2_X1 U658 ( .A1(n596), .A2(n595), .ZN(G290) );
  NOR2_X1 U659 ( .A1(G164), .A2(G1384), .ZN(n703) );
  AND2_X1 U660 ( .A1(G40), .A2(n703), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n600), .A2(G8), .ZN(n598) );
  XOR2_X1 U662 ( .A(KEYINPUT90), .B(n598), .Z(n719) );
  INV_X1 U663 ( .A(n719), .ZN(n679) );
  NAND2_X1 U664 ( .A1(n653), .A2(G1996), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n680), .A2(G1341), .ZN(n615) );
  NAND2_X1 U666 ( .A1(n601), .A2(n615), .ZN(n602) );
  NAND2_X1 U667 ( .A1(n602), .A2(KEYINPUT92), .ZN(n614) );
  XNOR2_X1 U668 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n608) );
  NAND2_X1 U669 ( .A1(n794), .A2(G81), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G68), .A2(n795), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U673 ( .A(n606), .B(KEYINPUT13), .ZN(n607) );
  XNOR2_X1 U674 ( .A(n608), .B(n607), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n790), .A2(G56), .ZN(n609) );
  XNOR2_X1 U676 ( .A(n609), .B(KEYINPUT14), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G43), .A2(n791), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U679 ( .A1(n613), .A2(n612), .ZN(n971) );
  NAND2_X1 U680 ( .A1(n614), .A2(n971), .ZN(n619) );
  INV_X1 U681 ( .A(KEYINPUT26), .ZN(n616) );
  NOR2_X1 U682 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U683 ( .A1(KEYINPUT92), .A2(n617), .ZN(n618) );
  NOR2_X1 U684 ( .A1(n619), .A2(n618), .ZN(n629) );
  NAND2_X1 U685 ( .A1(G79), .A2(n795), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G54), .A2(n791), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U688 ( .A(KEYINPUT72), .B(n622), .ZN(n626) );
  NAND2_X1 U689 ( .A1(G92), .A2(n794), .ZN(n624) );
  NAND2_X1 U690 ( .A1(G66), .A2(n790), .ZN(n623) );
  NAND2_X1 U691 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U692 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U693 ( .A(KEYINPUT15), .B(n627), .Z(n955) );
  NOR2_X1 U694 ( .A1(n629), .A2(n955), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n628), .B(KEYINPUT93), .ZN(n635) );
  NAND2_X1 U696 ( .A1(n629), .A2(n955), .ZN(n633) );
  NOR2_X1 U697 ( .A1(n653), .A2(G1348), .ZN(n631) );
  NOR2_X1 U698 ( .A1(G2067), .A2(n680), .ZN(n630) );
  NOR2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n647) );
  NAND2_X1 U702 ( .A1(G65), .A2(n790), .ZN(n637) );
  NAND2_X1 U703 ( .A1(G53), .A2(n791), .ZN(n636) );
  NAND2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U705 ( .A(KEYINPUT68), .B(n638), .ZN(n642) );
  NAND2_X1 U706 ( .A1(G91), .A2(n794), .ZN(n640) );
  NAND2_X1 U707 ( .A1(G78), .A2(n795), .ZN(n639) );
  NAND2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n956) );
  NAND2_X1 U710 ( .A1(n653), .A2(G2072), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n643), .B(KEYINPUT27), .ZN(n645) );
  AND2_X1 U712 ( .A1(G1956), .A2(n680), .ZN(n644) );
  NOR2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U714 ( .A1(n956), .A2(n648), .ZN(n646) );
  NAND2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n651) );
  NOR2_X1 U716 ( .A1(n956), .A2(n648), .ZN(n649) );
  XOR2_X1 U717 ( .A(n649), .B(KEYINPUT28), .Z(n650) );
  NAND2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U719 ( .A(KEYINPUT29), .B(n652), .ZN(n658) );
  NAND2_X1 U720 ( .A1(G1961), .A2(n680), .ZN(n655) );
  XOR2_X1 U721 ( .A(KEYINPUT25), .B(G2078), .Z(n1008) );
  NAND2_X1 U722 ( .A1(n653), .A2(n1008), .ZN(n654) );
  NAND2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n663) );
  NOR2_X1 U724 ( .A1(G301), .A2(n663), .ZN(n656) );
  XOR2_X1 U725 ( .A(KEYINPUT91), .B(n656), .Z(n657) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n670) );
  NOR2_X1 U727 ( .A1(G2084), .A2(n680), .ZN(n673) );
  NOR2_X1 U728 ( .A1(n673), .A2(n671), .ZN(n659) );
  NAND2_X1 U729 ( .A1(G8), .A2(n659), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U731 ( .A1(G168), .A2(n662), .ZN(n665) );
  AND2_X1 U732 ( .A1(G301), .A2(n663), .ZN(n664) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n668) );
  INV_X1 U734 ( .A(KEYINPUT95), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n676) );
  NOR2_X1 U737 ( .A1(n671), .A2(n676), .ZN(n672) );
  XOR2_X1 U738 ( .A(KEYINPUT96), .B(n672), .Z(n675) );
  AND2_X1 U739 ( .A1(G8), .A2(n673), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n690) );
  INV_X1 U741 ( .A(n676), .ZN(n678) );
  AND2_X1 U742 ( .A1(G286), .A2(G8), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n687) );
  INV_X1 U744 ( .A(G8), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n679), .A2(G1971), .ZN(n682) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n680), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n683), .A2(G303), .ZN(n684) );
  OR2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  AND2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U751 ( .A(n688), .B(KEYINPUT32), .Z(n689) );
  NOR2_X1 U752 ( .A1(n690), .A2(n689), .ZN(n717) );
  INV_X1 U753 ( .A(n717), .ZN(n693) );
  NOR2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n720) );
  NOR2_X1 U755 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U756 ( .A1(n720), .A2(n691), .ZN(n967) );
  XOR2_X1 U757 ( .A(n967), .B(KEYINPUT97), .Z(n692) );
  NAND2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NAND2_X1 U760 ( .A1(n694), .A2(n966), .ZN(n696) );
  XNOR2_X1 U761 ( .A(n696), .B(n695), .ZN(n699) );
  XOR2_X1 U762 ( .A(KEYINPUT99), .B(G1981), .Z(n697) );
  XNOR2_X1 U763 ( .A(G305), .B(n697), .ZN(n721) );
  NOR2_X1 U764 ( .A1(n721), .A2(KEYINPUT33), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U766 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XOR2_X1 U767 ( .A(n700), .B(KEYINPUT24), .Z(n701) );
  NAND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n714) );
  NOR2_X1 U769 ( .A1(n703), .A2(n522), .ZN(n760) );
  NAND2_X1 U770 ( .A1(G140), .A2(n877), .ZN(n705) );
  NAND2_X1 U771 ( .A1(G104), .A2(n874), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U773 ( .A(KEYINPUT34), .B(n706), .ZN(n711) );
  NAND2_X1 U774 ( .A1(G128), .A2(n869), .ZN(n708) );
  NAND2_X1 U775 ( .A1(G116), .A2(n870), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U777 ( .A(KEYINPUT35), .B(n709), .Z(n710) );
  NOR2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U779 ( .A(KEYINPUT36), .B(n712), .ZN(n867) );
  XNOR2_X1 U780 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  NOR2_X1 U781 ( .A1(n867), .A2(n758), .ZN(n924) );
  NAND2_X1 U782 ( .A1(n760), .A2(n924), .ZN(n756) );
  AND2_X1 U783 ( .A1(n719), .A2(n756), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n728) );
  INV_X1 U785 ( .A(n756), .ZN(n726) );
  NAND2_X1 U786 ( .A1(G166), .A2(G8), .ZN(n715) );
  NOR2_X1 U787 ( .A1(G2090), .A2(n715), .ZN(n716) );
  NOR2_X1 U788 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U789 ( .A1(n719), .A2(n718), .ZN(n724) );
  NAND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n723) );
  INV_X1 U791 ( .A(n721), .ZN(n952) );
  AND2_X1 U792 ( .A1(n952), .A2(KEYINPUT33), .ZN(n722) );
  NOR2_X1 U793 ( .A1(n724), .A2(n523), .ZN(n725) );
  OR2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U795 ( .A1(n728), .A2(n727), .ZN(n749) );
  NAND2_X1 U796 ( .A1(G117), .A2(n870), .ZN(n730) );
  NAND2_X1 U797 ( .A1(G141), .A2(n877), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U799 ( .A1(n874), .A2(G105), .ZN(n731) );
  XOR2_X1 U800 ( .A(KEYINPUT38), .B(n731), .Z(n732) );
  NOR2_X1 U801 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U802 ( .A1(n869), .A2(G129), .ZN(n734) );
  NAND2_X1 U803 ( .A1(n735), .A2(n734), .ZN(n863) );
  NAND2_X1 U804 ( .A1(n863), .A2(G1996), .ZN(n745) );
  NAND2_X1 U805 ( .A1(n870), .A2(G107), .ZN(n736) );
  XOR2_X1 U806 ( .A(KEYINPUT87), .B(n736), .Z(n738) );
  NAND2_X1 U807 ( .A1(n869), .A2(G119), .ZN(n737) );
  NAND2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U809 ( .A(KEYINPUT88), .B(n739), .Z(n743) );
  NAND2_X1 U810 ( .A1(G131), .A2(n877), .ZN(n741) );
  NAND2_X1 U811 ( .A1(G95), .A2(n874), .ZN(n740) );
  AND2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U813 ( .A1(n743), .A2(n742), .ZN(n860) );
  NAND2_X1 U814 ( .A1(G1991), .A2(n860), .ZN(n744) );
  NAND2_X1 U815 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U816 ( .A(n746), .B(KEYINPUT89), .ZN(n750) );
  XOR2_X1 U817 ( .A(G1986), .B(G290), .Z(n961) );
  NAND2_X1 U818 ( .A1(n750), .A2(n961), .ZN(n747) );
  NAND2_X1 U819 ( .A1(n747), .A2(n760), .ZN(n748) );
  NAND2_X1 U820 ( .A1(n749), .A2(n748), .ZN(n763) );
  INV_X1 U821 ( .A(n750), .ZN(n930) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n751) );
  NOR2_X1 U823 ( .A1(G1991), .A2(n860), .ZN(n926) );
  NOR2_X1 U824 ( .A1(n751), .A2(n926), .ZN(n752) );
  NOR2_X1 U825 ( .A1(n930), .A2(n752), .ZN(n754) );
  NOR2_X1 U826 ( .A1(n863), .A2(G1996), .ZN(n753) );
  XNOR2_X1 U827 ( .A(n753), .B(KEYINPUT100), .ZN(n941) );
  NOR2_X1 U828 ( .A1(n754), .A2(n941), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n755), .B(KEYINPUT39), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U831 ( .A1(n867), .A2(n758), .ZN(n927) );
  NAND2_X1 U832 ( .A1(n759), .A2(n927), .ZN(n761) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U835 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U836 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U837 ( .A(G57), .ZN(G237) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U839 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n837) );
  NAND2_X1 U841 ( .A1(n837), .A2(G567), .ZN(n766) );
  XOR2_X1 U842 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  NAND2_X1 U843 ( .A1(n971), .A2(G860), .ZN(G153) );
  NAND2_X1 U844 ( .A1(G868), .A2(G301), .ZN(n768) );
  OR2_X1 U845 ( .A1(n955), .A2(G868), .ZN(n767) );
  NAND2_X1 U846 ( .A1(n768), .A2(n767), .ZN(G284) );
  XNOR2_X1 U847 ( .A(n956), .B(KEYINPUT69), .ZN(G299) );
  INV_X1 U848 ( .A(G868), .ZN(n775) );
  NOR2_X1 U849 ( .A1(G286), .A2(n775), .ZN(n769) );
  XOR2_X1 U850 ( .A(KEYINPUT77), .B(n769), .Z(n771) );
  NOR2_X1 U851 ( .A1(G868), .A2(G299), .ZN(n770) );
  NOR2_X1 U852 ( .A1(n771), .A2(n770), .ZN(G297) );
  INV_X1 U853 ( .A(G860), .ZN(n789) );
  NAND2_X1 U854 ( .A1(n789), .A2(G559), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n772), .A2(n955), .ZN(n773) );
  XNOR2_X1 U856 ( .A(n773), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U857 ( .A1(n955), .A2(G868), .ZN(n774) );
  NOR2_X1 U858 ( .A1(G559), .A2(n774), .ZN(n777) );
  AND2_X1 U859 ( .A1(n775), .A2(n971), .ZN(n776) );
  NOR2_X1 U860 ( .A1(n777), .A2(n776), .ZN(G282) );
  NAND2_X1 U861 ( .A1(n869), .A2(G123), .ZN(n778) );
  XNOR2_X1 U862 ( .A(n778), .B(KEYINPUT18), .ZN(n780) );
  NAND2_X1 U863 ( .A1(G135), .A2(n877), .ZN(n779) );
  NAND2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n784) );
  NAND2_X1 U865 ( .A1(G111), .A2(n870), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G99), .A2(n874), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U868 ( .A1(n784), .A2(n783), .ZN(n925) );
  XNOR2_X1 U869 ( .A(G2096), .B(n925), .ZN(n785) );
  XNOR2_X1 U870 ( .A(n785), .B(KEYINPUT78), .ZN(n787) );
  INV_X1 U871 ( .A(G2100), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G559), .A2(n955), .ZN(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(n971), .ZN(n807) );
  NAND2_X1 U875 ( .A1(n789), .A2(n807), .ZN(n800) );
  NAND2_X1 U876 ( .A1(G67), .A2(n790), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G55), .A2(n791), .ZN(n792) );
  NAND2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n799) );
  NAND2_X1 U879 ( .A1(G93), .A2(n794), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G80), .A2(n795), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U882 ( .A1(n799), .A2(n798), .ZN(n809) );
  XOR2_X1 U883 ( .A(n800), .B(n809), .Z(G145) );
  XNOR2_X1 U884 ( .A(G166), .B(n809), .ZN(n805) );
  XOR2_X1 U885 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n801) );
  XNOR2_X1 U886 ( .A(G305), .B(n801), .ZN(n802) );
  XNOR2_X1 U887 ( .A(n802), .B(G290), .ZN(n803) );
  XNOR2_X1 U888 ( .A(n803), .B(G299), .ZN(n804) );
  XNOR2_X1 U889 ( .A(n805), .B(n804), .ZN(n806) );
  XNOR2_X1 U890 ( .A(n806), .B(G288), .ZN(n887) );
  XNOR2_X1 U891 ( .A(n807), .B(n887), .ZN(n808) );
  NAND2_X1 U892 ( .A1(n808), .A2(G868), .ZN(n811) );
  OR2_X1 U893 ( .A1(G868), .A2(n809), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U895 ( .A1(G2084), .A2(G2078), .ZN(n813) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n812) );
  XNOR2_X1 U897 ( .A(n813), .B(n812), .ZN(n814) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n814), .ZN(n815) );
  XNOR2_X1 U899 ( .A(KEYINPUT21), .B(n815), .ZN(n816) );
  NAND2_X1 U900 ( .A1(n816), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U901 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U902 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n818) );
  NAND2_X1 U903 ( .A1(G132), .A2(G82), .ZN(n817) );
  XNOR2_X1 U904 ( .A(n818), .B(n817), .ZN(n819) );
  NOR2_X1 U905 ( .A1(n819), .A2(G218), .ZN(n820) );
  NAND2_X1 U906 ( .A1(G96), .A2(n820), .ZN(n921) );
  NAND2_X1 U907 ( .A1(n921), .A2(G2106), .ZN(n824) );
  NAND2_X1 U908 ( .A1(G69), .A2(G120), .ZN(n821) );
  NOR2_X1 U909 ( .A1(G237), .A2(n821), .ZN(n822) );
  NAND2_X1 U910 ( .A1(G108), .A2(n822), .ZN(n922) );
  NAND2_X1 U911 ( .A1(n922), .A2(G567), .ZN(n823) );
  NAND2_X1 U912 ( .A1(n824), .A2(n823), .ZN(n891) );
  NAND2_X1 U913 ( .A1(G483), .A2(G661), .ZN(n825) );
  NOR2_X1 U914 ( .A1(n891), .A2(n825), .ZN(n840) );
  NAND2_X1 U915 ( .A1(n840), .A2(G36), .ZN(G176) );
  XNOR2_X1 U916 ( .A(G2427), .B(G2443), .ZN(n835) );
  XOR2_X1 U917 ( .A(G2430), .B(KEYINPUT102), .Z(n827) );
  XNOR2_X1 U918 ( .A(G2454), .B(G2435), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U920 ( .A(G2438), .B(KEYINPUT101), .Z(n829) );
  XNOR2_X1 U921 ( .A(G1348), .B(G1341), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U923 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U924 ( .A(G2446), .B(G2451), .ZN(n832) );
  XNOR2_X1 U925 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U926 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U927 ( .A1(n836), .A2(G14), .ZN(n913) );
  XNOR2_X1 U928 ( .A(KEYINPUT103), .B(n913), .ZN(G401) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U931 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n840), .A2(n839), .ZN(G188) );
  NAND2_X1 U934 ( .A1(n869), .A2(G124), .ZN(n841) );
  XNOR2_X1 U935 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U936 ( .A1(G112), .A2(n870), .ZN(n842) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U938 ( .A1(G136), .A2(n877), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G100), .A2(n874), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U941 ( .A1(n847), .A2(n846), .ZN(G162) );
  XOR2_X1 U942 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n849) );
  XNOR2_X1 U943 ( .A(G162), .B(KEYINPUT109), .ZN(n848) );
  XNOR2_X1 U944 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U945 ( .A(n925), .B(n850), .ZN(n865) );
  NAND2_X1 U946 ( .A1(n870), .A2(G118), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT107), .B(n851), .Z(n853) );
  NAND2_X1 U948 ( .A1(n869), .A2(G130), .ZN(n852) );
  NAND2_X1 U949 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U950 ( .A(KEYINPUT108), .B(n854), .ZN(n859) );
  NAND2_X1 U951 ( .A1(G142), .A2(n877), .ZN(n856) );
  NAND2_X1 U952 ( .A1(G106), .A2(n874), .ZN(n855) );
  NAND2_X1 U953 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U954 ( .A(n857), .B(KEYINPUT45), .Z(n858) );
  NOR2_X1 U955 ( .A1(n859), .A2(n858), .ZN(n861) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U957 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U958 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U959 ( .A(n866), .B(G160), .ZN(n868) );
  XNOR2_X1 U960 ( .A(n868), .B(n867), .ZN(n882) );
  NAND2_X1 U961 ( .A1(G127), .A2(n869), .ZN(n872) );
  NAND2_X1 U962 ( .A1(G115), .A2(n870), .ZN(n871) );
  NAND2_X1 U963 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U964 ( .A(n873), .B(KEYINPUT47), .ZN(n876) );
  NAND2_X1 U965 ( .A1(G103), .A2(n874), .ZN(n875) );
  NAND2_X1 U966 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U967 ( .A1(n877), .A2(G139), .ZN(n878) );
  XOR2_X1 U968 ( .A(KEYINPUT110), .B(n878), .Z(n879) );
  NOR2_X1 U969 ( .A1(n880), .A2(n879), .ZN(n933) );
  XNOR2_X1 U970 ( .A(G164), .B(n933), .ZN(n881) );
  XNOR2_X1 U971 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U972 ( .A1(G37), .A2(n883), .ZN(n884) );
  XOR2_X1 U973 ( .A(KEYINPUT111), .B(n884), .Z(G395) );
  XNOR2_X1 U974 ( .A(G286), .B(KEYINPUT112), .ZN(n886) );
  XNOR2_X1 U975 ( .A(G171), .B(n971), .ZN(n885) );
  XNOR2_X1 U976 ( .A(n886), .B(n885), .ZN(n889) );
  XOR2_X1 U977 ( .A(n955), .B(n887), .Z(n888) );
  XNOR2_X1 U978 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U979 ( .A1(G37), .A2(n890), .ZN(G397) );
  INV_X1 U980 ( .A(n891), .ZN(G319) );
  XOR2_X1 U981 ( .A(G2474), .B(G1966), .Z(n893) );
  XNOR2_X1 U982 ( .A(G1996), .B(G1991), .ZN(n892) );
  XNOR2_X1 U983 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U984 ( .A(n894), .B(KEYINPUT105), .Z(n896) );
  XNOR2_X1 U985 ( .A(G1986), .B(G1961), .ZN(n895) );
  XNOR2_X1 U986 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U987 ( .A(G1971), .B(G1956), .Z(n898) );
  XNOR2_X1 U988 ( .A(G1981), .B(G1976), .ZN(n897) );
  XNOR2_X1 U989 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U990 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U991 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n901) );
  XNOR2_X1 U992 ( .A(n902), .B(n901), .ZN(G229) );
  XOR2_X1 U993 ( .A(G2096), .B(KEYINPUT43), .Z(n904) );
  XNOR2_X1 U994 ( .A(G2090), .B(KEYINPUT104), .ZN(n903) );
  XNOR2_X1 U995 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U996 ( .A(n905), .B(G2678), .Z(n907) );
  XNOR2_X1 U997 ( .A(G2067), .B(G2072), .ZN(n906) );
  XNOR2_X1 U998 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U999 ( .A(KEYINPUT42), .B(G2100), .Z(n909) );
  XNOR2_X1 U1000 ( .A(G2084), .B(G2078), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1002 ( .A(n911), .B(n910), .ZN(G227) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n912) );
  XOR2_X1 U1004 ( .A(KEYINPUT115), .B(n912), .Z(n920) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n913), .ZN(n914) );
  XOR2_X1 U1006 ( .A(KEYINPUT113), .B(n914), .Z(n917) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n915) );
  XNOR2_X1 U1008 ( .A(n915), .B(KEYINPUT49), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(KEYINPUT114), .B(n918), .ZN(n919) );
  NAND2_X1 U1011 ( .A1(n920), .A2(n919), .ZN(G225) );
  XOR2_X1 U1012 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1014 ( .A(G132), .ZN(G219) );
  INV_X1 U1015 ( .A(G120), .ZN(G236) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  INV_X1 U1017 ( .A(G82), .ZN(G220) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(G325) );
  INV_X1 U1020 ( .A(G325), .ZN(G261) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n932) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n946) );
  XOR2_X1 U1028 ( .A(G2072), .B(n933), .Z(n934) );
  XNOR2_X1 U1029 ( .A(KEYINPUT117), .B(n934), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(G164), .B(G2078), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(n935), .B(KEYINPUT118), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(n938), .B(KEYINPUT50), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(KEYINPUT119), .B(n939), .ZN(n944) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n942), .Z(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n950), .A2(G29), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT120), .B(n951), .ZN(n1031) );
  XNOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .ZN(n977) );
  XNOR2_X1 U1046 ( .A(G1966), .B(G168), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT57), .B(n954), .ZN(n975) );
  XNOR2_X1 U1049 ( .A(G1348), .B(n955), .ZN(n965) );
  XNOR2_X1 U1050 ( .A(n956), .B(G1956), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(G1971), .A2(G303), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(G1961), .B(KEYINPUT123), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(G301), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n969) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1060 ( .A(KEYINPUT124), .B(n970), .Z(n973) );
  XOR2_X1 U1061 ( .A(n971), .B(G1341), .Z(n972) );
  NOR2_X1 U1062 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1063 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1064 ( .A1(n977), .A2(n976), .ZN(n1005) );
  INV_X1 U1065 ( .A(G16), .ZN(n1003) );
  INV_X1 U1066 ( .A(G1341), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G19), .B(n978), .ZN(n982) );
  XNOR2_X1 U1068 ( .A(G1981), .B(G6), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G20), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1072 ( .A(KEYINPUT59), .B(G1348), .Z(n983) );
  XNOR2_X1 U1073 ( .A(G4), .B(n983), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1075 ( .A(KEYINPUT60), .B(n986), .Z(n988) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G21), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n998) );
  XNOR2_X1 U1078 ( .A(G1976), .B(KEYINPUT126), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n989), .B(G23), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(G1986), .B(KEYINPUT127), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(G24), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(G1971), .B(KEYINPUT125), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(G22), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n996), .B(KEYINPUT58), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G5), .B(G1961), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(KEYINPUT61), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1029) );
  XNOR2_X1 U1093 ( .A(G2067), .B(G26), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1996), .B(G32), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1008), .B(G27), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G33), .B(G2072), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT121), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(G28), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G25), .B(G1991), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(KEYINPUT53), .B(n1017), .Z(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT54), .B(G34), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(G2084), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(G35), .B(G2090), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(n1023), .B(KEYINPUT55), .ZN(n1025) );
  INV_X1 U1111 ( .A(G29), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(G11), .A2(n1026), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(KEYINPUT122), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

