//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT25), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(KEYINPUT23), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT66), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT24), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n213), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n211), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n212), .B1(new_n228), .B2(new_n219), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n224), .A2(new_n225), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(KEYINPUT68), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n210), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT65), .B(G176gat), .Z(new_n233));
  NOR2_X1   g032(.A1(new_n206), .A2(G169gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n209), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT64), .B1(new_n237), .B2(new_n212), .ZN(new_n238));
  INV_X1    g037(.A(new_n222), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT25), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n203), .B1(new_n232), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n210), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n221), .A2(new_n211), .A3(new_n226), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT68), .B1(new_n229), .B2(new_n230), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n241), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(KEYINPUT69), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT27), .B(G183gat), .ZN(new_n249));
  INV_X1    g048(.A(G190gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n251), .A2(KEYINPUT70), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(KEYINPUT70), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n204), .B1(new_n257), .B2(new_n208), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n212), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n248), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n265));
  INV_X1    g064(.A(G120gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(G113gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT71), .B(G120gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n268), .B2(G113gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n269), .A2(new_n271), .A3(KEYINPUT72), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(KEYINPUT71), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G120gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n276), .A3(G113gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n267), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G127gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(G134gat), .ZN(new_n281));
  INV_X1    g080(.A(G134gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G127gat), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n281), .A2(new_n283), .A3(KEYINPUT1), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n273), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n265), .B1(new_n272), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n261), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n242), .A2(new_n248), .A3(new_n260), .A4(new_n286), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G227gat), .ZN(new_n291));
  INV_X1    g090(.A(G233gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n202), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  AOI211_X1 g094(.A(KEYINPUT34), .B(new_n293), .C1(new_n288), .C2(new_n289), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n288), .A2(new_n293), .A3(new_n289), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT33), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G15gat), .B(G43gat), .Z(new_n302));
  XNOR2_X1  g101(.A(G71gat), .B(G99gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n298), .B(KEYINPUT32), .C1(new_n300), .C2(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n297), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n295), .ZN(new_n309));
  INV_X1    g108(.A(new_n296), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n305), .A2(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G78gat), .B(G106gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT80), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT31), .B(G50gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n317), .A3(new_n321), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n316), .B1(new_n328), .B2(KEYINPUT29), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n330));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(G141gat), .B(G148gat), .Z(new_n335));
  INV_X1    g134(.A(G155gat), .ZN(new_n336));
  INV_X1    g135(.A(G162gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(KEYINPUT77), .A3(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(KEYINPUT2), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(KEYINPUT76), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n331), .B1(new_n333), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n340), .ZN(new_n345));
  XNOR2_X1  g144(.A(G141gat), .B(G148gat), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n342), .B(new_n344), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(G228gat), .A2(G233gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n341), .A2(new_n347), .A3(new_n316), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n327), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n349), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G22gat), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n352), .B1(new_n325), .B2(new_n326), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT3), .B1(new_n358), .B2(KEYINPUT81), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(KEYINPUT81), .B2(new_n358), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n354), .B1(new_n360), .B2(new_n348), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n356), .B(new_n357), .C1(new_n361), .C2(new_n350), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n315), .B1(new_n362), .B2(KEYINPUT82), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(KEYINPUT81), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n316), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n358), .A2(KEYINPUT81), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n348), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n350), .B1(new_n367), .B2(new_n355), .ZN(new_n368));
  INV_X1    g167(.A(new_n356), .ZN(new_n369));
  OAI21_X1  g168(.A(G22gat), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n362), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n370), .B(new_n362), .C1(KEYINPUT82), .C2(new_n315), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n308), .A2(new_n311), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT0), .ZN(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g178(.A(KEYINPUT5), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n286), .A2(new_n348), .ZN(new_n383));
  INV_X1    g182(.A(new_n348), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT72), .B1(new_n269), .B2(new_n271), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n279), .A2(new_n284), .A3(new_n273), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n265), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n382), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT78), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n286), .B2(new_n348), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n286), .A2(new_n393), .A3(new_n351), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n387), .A2(new_n384), .A3(KEYINPUT4), .A4(new_n265), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n381), .A4(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n380), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n392), .A2(new_n395), .A3(new_n394), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(new_n382), .C1(new_n383), .C2(new_n388), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n398), .A2(new_n381), .B1(new_n400), .B2(KEYINPUT5), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n379), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n286), .A2(new_n348), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n384), .A3(new_n265), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n381), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n396), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n408));
  INV_X1    g207(.A(new_n379), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n396), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(new_n403), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n403), .B2(new_n412), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n242), .A2(new_n248), .A3(new_n260), .A4(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n232), .A2(new_n241), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n255), .A2(new_n259), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n419), .B(new_n416), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n327), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n352), .A2(new_n417), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n261), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n420), .A2(new_n421), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n417), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n328), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(G8gat), .B(G36gat), .Z(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT75), .ZN(new_n432));
  XOR2_X1   g231(.A(G64gat), .B(G92gat), .Z(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n415), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n430), .A2(new_n435), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n328), .B1(new_n418), .B2(new_n422), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n261), .A2(new_n425), .B1(new_n427), .B2(new_n417), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n328), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT30), .A3(new_n434), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n414), .A2(new_n438), .A3(new_n439), .A4(new_n443), .ZN(new_n444));
  NOR4_X1   g243(.A1(new_n397), .A2(new_n401), .A3(new_n403), .A4(new_n379), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n397), .A2(new_n401), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT6), .B1(new_n446), .B2(new_n409), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n447), .B2(new_n402), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n443), .B1(new_n436), .B2(new_n437), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT79), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n375), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n445), .B1(new_n413), .B2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n447), .A2(new_n454), .A3(new_n402), .ZN(new_n455));
  AOI211_X1 g254(.A(KEYINPUT35), .B(new_n449), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n375), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n444), .A2(new_n450), .A3(new_n374), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n434), .B1(new_n442), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n441), .B2(new_n327), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n423), .A2(new_n328), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT38), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n437), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n435), .B1(new_n430), .B2(KEYINPUT37), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n460), .B1(new_n424), .B2(new_n429), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT38), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n453), .A2(new_n465), .A3(new_n455), .A4(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n412), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n392), .A2(new_n395), .A3(new_n394), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n382), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n379), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT83), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n476), .A3(new_n379), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(new_n382), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n383), .A2(new_n388), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n472), .B1(new_n479), .B2(new_n381), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n475), .A2(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n470), .B1(new_n481), .B2(KEYINPUT40), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(new_n449), .C1(KEYINPUT40), .C2(new_n481), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n374), .B1(new_n469), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n459), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n308), .B2(new_n311), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n305), .A2(new_n307), .ZN(new_n489));
  INV_X1    g288(.A(new_n297), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n297), .A2(new_n305), .A3(new_n307), .ZN(new_n492));
  NOR2_X1   g291(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n458), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  INV_X1    g297(.A(G1gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(KEYINPUT16), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n498), .A2(new_n499), .ZN(new_n502));
  OAI21_X1  g301(.A(G8gat), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G8gat), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n500), .B(new_n504), .C1(new_n499), .C2(new_n498), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT14), .ZN(new_n508));
  INV_X1    g307(.A(G29gat), .ZN(new_n509));
  INV_X1    g308(.A(G36gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n511), .A2(new_n512), .B1(G29gat), .B2(G36gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n507), .B1(new_n513), .B2(KEYINPUT15), .ZN(new_n514));
  INV_X1    g313(.A(new_n512), .ZN(new_n515));
  NOR3_X1   g314(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n515), .A2(new_n516), .B1(new_n509), .B2(new_n510), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n517), .A2(new_n518), .A3(new_n507), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n520), .A2(KEYINPUT17), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  INV_X1    g322(.A(new_n521), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n507), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n523), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n506), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n503), .A2(new_n505), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n527), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT18), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n529), .A2(KEYINPUT18), .A3(new_n530), .A4(new_n533), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT11), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT85), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  XOR2_X1   g342(.A(G169gat), .B(G197gat), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n542), .B2(new_n543), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT12), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n531), .B(new_n532), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n530), .B(KEYINPUT13), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n537), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT86), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n556), .A2(new_n537), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT86), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n559), .A2(new_n560), .A3(new_n536), .A4(new_n553), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n536), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n549), .A3(new_n552), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT41), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT90), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(KEYINPUT8), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT91), .A3(KEYINPUT7), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(G85gat), .A3(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT91), .B1(new_n573), .B2(KEYINPUT7), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n572), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n580), .B(new_n572), .C1(new_n577), .C2(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n522), .B2(new_n528), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n566), .A2(KEYINPUT41), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n584), .ZN(new_n589));
  AOI211_X1 g388(.A(new_n586), .B(new_n588), .C1(new_n589), .C2(new_n532), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n583), .B(new_n582), .C1(new_n520), .C2(new_n521), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT92), .B1(new_n591), .B2(new_n587), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n585), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT93), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n595), .B(new_n585), .C1(new_n590), .C2(new_n592), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n597), .B2(new_n598), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n569), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G57gat), .B(G64gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G71gat), .ZN(new_n609));
  INV_X1    g408(.A(G78gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT9), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n608), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n612), .B(new_n611), .C1(new_n607), .C2(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n619), .B1(new_n618), .B2(new_n620), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n606), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n618), .A2(new_n620), .ZN(new_n625));
  INV_X1    g424(.A(new_n619), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n621), .A3(new_n605), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT88), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n624), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n624), .B2(new_n628), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n604), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n631), .A3(new_n603), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT21), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n506), .B1(new_n638), .B2(new_n618), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT89), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n634), .A2(new_n636), .A3(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n599), .ZN(new_n645));
  INV_X1    g444(.A(new_n598), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n584), .B1(new_n524), .B2(new_n527), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n586), .B1(new_n647), .B2(new_n588), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n591), .A2(KEYINPUT92), .A3(new_n587), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n595), .B1(new_n650), .B2(new_n585), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n645), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n568), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n602), .A2(new_n644), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n602), .A2(new_n644), .A3(new_n654), .A4(KEYINPUT94), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT95), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n583), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n582), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n579), .A2(new_n661), .A3(new_n581), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n618), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n618), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n584), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n660), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n666), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n665), .A2(new_n667), .A3(new_n671), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n672), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n659), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n497), .A2(new_n565), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n414), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(new_n499), .ZN(G1324gat));
  AND2_X1   g484(.A1(new_n497), .A2(new_n565), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n449), .A3(new_n682), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G8gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT42), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  MUX2_X1   g490(.A(new_n689), .B(KEYINPUT42), .S(new_n691), .Z(G1325gat));
  INV_X1    g491(.A(new_n494), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n308), .A2(new_n311), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n486), .B1(new_n491), .B2(new_n492), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT96), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT96), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n488), .A2(new_n495), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT97), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(KEYINPUT97), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n683), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n308), .A2(new_n311), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n683), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT98), .ZN(G1326gat));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n686), .A2(KEYINPUT99), .A3(new_n374), .A4(new_n682), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT99), .ZN(new_n712));
  INV_X1    g511(.A(new_n374), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n683), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n710), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n711), .A2(new_n710), .A3(new_n714), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT43), .B(G22gat), .Z(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(G1327gat));
  NAND2_X1  g521(.A1(new_n602), .A2(new_n654), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n469), .A2(new_n483), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n713), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n444), .A2(new_n450), .A3(new_n374), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n496), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n451), .A2(KEYINPUT35), .B1(new_n456), .B2(new_n375), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT44), .B(new_n723), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n644), .ZN(new_n730));
  INV_X1    g529(.A(new_n681), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n565), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n723), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n488), .A2(new_n697), .A3(new_n495), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n697), .B1(new_n488), .B2(new_n495), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n459), .A2(new_n484), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n738), .B2(new_n458), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n729), .B(new_n734), .C1(new_n739), .C2(KEYINPUT44), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n740), .A2(KEYINPUT102), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(KEYINPUT102), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G29gat), .B1(new_n743), .B2(new_n414), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n735), .A2(new_n732), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT101), .Z(new_n746));
  NAND3_X1  g545(.A1(new_n497), .A2(new_n565), .A3(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(G29gat), .A3(new_n414), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT45), .Z(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n749), .ZN(G1328gat));
  INV_X1    g549(.A(new_n449), .ZN(new_n751));
  OAI21_X1  g550(.A(G36gat), .B1(new_n743), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n747), .A2(G36gat), .A3(new_n751), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1329gat));
  NOR2_X1   g554(.A1(new_n706), .A2(G43gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n747), .A2(KEYINPUT103), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT103), .B1(new_n747), .B2(new_n757), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G43gat), .B1(new_n740), .B2(new_n699), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n703), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n741), .A2(new_n763), .A3(new_n742), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n764), .A2(G43gat), .B1(new_n759), .B2(new_n758), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g565(.A1(new_n713), .A2(G50gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n747), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n747), .A2(KEYINPUT105), .A3(new_n767), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT106), .B1(new_n740), .B2(new_n713), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G50gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n740), .A2(KEYINPUT106), .A3(new_n713), .ZN(new_n774));
  OAI221_X1 g573(.A(KEYINPUT48), .B1(new_n770), .B2(new_n771), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n768), .B(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n741), .A2(new_n374), .A3(new_n742), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(G50gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n775), .B1(new_n779), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g579(.A1(new_n659), .A2(new_n565), .A3(new_n731), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT107), .Z(new_n782));
  NAND2_X1  g581(.A1(new_n738), .A2(new_n458), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n414), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT108), .B(G57gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1332gat));
  INV_X1    g586(.A(new_n784), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT109), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n790), .B(new_n792), .ZN(G1333gat));
  OAI21_X1  g592(.A(new_n609), .B1(new_n784), .B2(new_n706), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n763), .A2(G71gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g596(.A1(new_n784), .A2(new_n713), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(new_n610), .ZN(G1335gat));
  NAND2_X1  g598(.A1(new_n733), .A2(new_n730), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT110), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n681), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n729), .B(new_n802), .C1(new_n739), .C2(KEYINPUT44), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n414), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n725), .A2(new_n726), .B1(new_n696), .B2(new_n698), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n723), .B(new_n801), .C1(new_n805), .C2(new_n728), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n783), .A2(KEYINPUT51), .A3(new_n723), .A4(new_n801), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n414), .A2(G85gat), .A3(new_n731), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n804), .B1(new_n811), .B2(new_n812), .ZN(G1336gat));
  OAI21_X1  g612(.A(G92gat), .B1(new_n803), .B2(new_n751), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n808), .A2(KEYINPUT112), .A3(new_n809), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n806), .A2(new_n816), .A3(new_n807), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n751), .A2(G92gat), .A3(new_n731), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT111), .Z(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT52), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n814), .B(new_n823), .C1(new_n811), .C2(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1337gat));
  OAI21_X1  g624(.A(G99gat), .B1(new_n803), .B2(new_n703), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n706), .A2(G99gat), .A3(new_n731), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n811), .B2(new_n827), .ZN(G1338gat));
  NOR3_X1   g627(.A1(new_n713), .A2(new_n731), .A3(G106gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n815), .A2(new_n817), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G106gat), .B1(new_n803), .B2(new_n713), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT53), .ZN(new_n833));
  INV_X1    g632(.A(new_n809), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT51), .B1(new_n739), .B2(new_n801), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n831), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n833), .A2(KEYINPUT113), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n837), .B1(new_n830), .B2(new_n831), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n831), .A2(new_n836), .A3(new_n837), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(G1339gat));
  NAND4_X1  g643(.A1(new_n657), .A2(new_n733), .A3(new_n658), .A4(new_n731), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n671), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n668), .A2(new_n669), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n672), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n668), .B2(new_n669), .ZN(new_n851));
  XNOR2_X1  g650(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n679), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(KEYINPUT55), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n680), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT116), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n857), .A3(new_n680), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n850), .A2(new_n853), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n565), .A2(new_n856), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n554), .A2(new_n555), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n529), .A2(new_n533), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(G229gat), .A3(G233gat), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n864), .A2(new_n866), .B1(new_n546), .B2(new_n550), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n558), .B2(new_n561), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n863), .B1(new_n868), .B2(new_n681), .ZN(new_n869));
  INV_X1    g668(.A(new_n867), .ZN(new_n870));
  AND4_X1   g669(.A1(new_n863), .A2(new_n562), .A3(new_n681), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n862), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n735), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n858), .A3(new_n861), .ZN(new_n874));
  INV_X1    g673(.A(new_n868), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n874), .A2(new_n735), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n644), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT118), .B1(new_n847), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n845), .B(KEYINPUT114), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n868), .A2(new_n681), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT117), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n868), .A2(new_n863), .A3(new_n681), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n723), .B1(new_n884), .B2(new_n862), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n874), .A2(new_n735), .A3(new_n875), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n730), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n879), .A2(new_n880), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n414), .A2(new_n449), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n878), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n375), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n733), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n892), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g692(.A1(new_n891), .A2(new_n731), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n268), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n266), .B2(new_n894), .ZN(G1341gat));
  NOR2_X1   g695(.A1(new_n891), .A2(new_n730), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(new_n280), .ZN(G1342gat));
  INV_X1    g697(.A(new_n375), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n735), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n890), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G134gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n901), .B2(G134gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n890), .A2(KEYINPUT119), .A3(new_n282), .A4(new_n900), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n904), .A2(KEYINPUT56), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT56), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(G1343gat));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n713), .B1(new_n701), .B2(new_n702), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n878), .A2(new_n888), .A3(new_n910), .A4(new_n889), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(G141gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n565), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n909), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n699), .A2(new_n889), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n699), .A2(KEYINPUT120), .A3(new_n889), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n878), .A2(new_n374), .A3(new_n888), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n565), .A2(new_n680), .A3(new_n854), .A4(new_n861), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n723), .B1(new_n925), .B2(new_n881), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n730), .B1(new_n886), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n879), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n713), .A2(new_n923), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n921), .B1(new_n924), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n913), .B1(new_n931), .B2(new_n565), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n911), .A2(G141gat), .A3(new_n733), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n916), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT58), .B1(new_n933), .B2(KEYINPUT121), .ZN(new_n935));
  AOI211_X1 g734(.A(new_n733), .B(new_n921), .C1(new_n924), .C2(new_n930), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n935), .B(new_n914), .C1(new_n936), .C2(new_n913), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(G1344gat));
  INV_X1    g737(.A(G148gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n912), .A2(new_n939), .A3(new_n681), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT59), .B(new_n939), .C1(new_n931), .C2(new_n681), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n921), .B(KEYINPUT122), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n845), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n845), .A2(new_n945), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n927), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n923), .A3(new_n374), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n943), .A2(new_n944), .A3(new_n681), .A4(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n942), .B1(new_n950), .B2(G148gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n940), .B1(new_n941), .B2(new_n951), .ZN(G1345gat));
  INV_X1    g751(.A(new_n931), .ZN(new_n953));
  OAI21_X1  g752(.A(G155gat), .B1(new_n953), .B2(new_n730), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n912), .A2(new_n336), .A3(new_n644), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1346gat));
  OAI21_X1  g755(.A(G162gat), .B1(new_n953), .B2(new_n735), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n912), .A2(new_n337), .A3(new_n723), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n899), .A2(new_n751), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n878), .A2(new_n888), .A3(new_n414), .A4(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n565), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n964), .A3(G169gat), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n964), .B1(new_n963), .B2(G169gat), .ZN(new_n967));
  OAI22_X1  g766(.A1(new_n966), .A2(new_n967), .B1(G169gat), .B2(new_n963), .ZN(G1348gat));
  NOR2_X1   g767(.A1(new_n961), .A2(new_n731), .ZN(new_n969));
  MUX2_X1   g768(.A(G176gat), .B(new_n233), .S(new_n969), .Z(G1349gat));
  NAND3_X1  g769(.A1(new_n962), .A2(new_n249), .A3(new_n644), .ZN(new_n971));
  OAI21_X1  g770(.A(G183gat), .B1(new_n961), .B2(new_n730), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(KEYINPUT125), .A3(new_n972), .ZN(new_n973));
  XOR2_X1   g772(.A(KEYINPUT126), .B(KEYINPUT60), .Z(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n973), .B(new_n975), .ZN(G1350gat));
  NAND2_X1  g775(.A1(new_n962), .A2(new_n723), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(new_n978), .A3(G190gat), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n978), .B1(new_n977), .B2(G190gat), .ZN(new_n981));
  OAI22_X1  g780(.A1(new_n980), .A2(new_n981), .B1(G190gat), .B2(new_n977), .ZN(G1351gat));
  NAND2_X1  g781(.A1(new_n910), .A2(new_n449), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n878), .A2(new_n414), .A3(new_n888), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(G197gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(new_n988), .A3(new_n565), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n944), .A2(new_n949), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n763), .A2(new_n448), .A3(new_n751), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n990), .A2(new_n565), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n992), .B2(new_n988), .ZN(G1352gat));
  NAND3_X1  g792(.A1(new_n990), .A2(new_n681), .A3(new_n991), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(G204gat), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n731), .A2(G204gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT62), .B1(new_n987), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n998));
  INV_X1    g797(.A(new_n996), .ZN(new_n999));
  NOR4_X1   g798(.A1(new_n985), .A2(new_n998), .A3(new_n986), .A4(new_n999), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n995), .B1(new_n997), .B2(new_n1000), .ZN(G1353gat));
  NAND3_X1  g800(.A1(new_n987), .A2(new_n319), .A3(new_n644), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n944), .A2(new_n644), .A3(new_n949), .A4(new_n991), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(G1354gat));
  NAND3_X1  g805(.A1(new_n987), .A2(new_n320), .A3(new_n723), .ZN(new_n1007));
  AND3_X1   g806(.A1(new_n990), .A2(new_n723), .A3(new_n991), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1007), .B1(new_n1008), .B2(new_n320), .ZN(G1355gat));
endmodule


