//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT78), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT37), .ZN(new_n206));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT67), .B(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT27), .B(G183gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT28), .A3(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT27), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n209), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n212), .B1(new_n218), .B2(KEYINPUT28), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR3_X1   g022(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G169gat), .A3(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n220), .A2(KEYINPUT24), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT66), .B(G183gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(new_n209), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n233), .A2(new_n222), .ZN(new_n247));
  NOR2_X1   g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(new_n239), .B2(new_n241), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n227), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n227), .B2(new_n251), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n208), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n227), .A2(new_n251), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n208), .A2(KEYINPUT29), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G211gat), .A2(G218gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT22), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(G197gat), .A2(G204gat), .ZN(new_n263));
  AND2_X1   g062(.A1(G197gat), .A2(G204gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G211gat), .B(G218gat), .Z(new_n266));
  INV_X1    g065(.A(KEYINPUT74), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G197gat), .ZN(new_n269));
  INV_X1    g068(.A(G204gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n271), .A2(new_n272), .B1(new_n261), .B2(new_n260), .ZN(new_n273));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT74), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n266), .B1(new_n265), .B2(KEYINPUT73), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n268), .A2(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT77), .B1(new_n259), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT77), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n267), .B1(new_n265), .B2(new_n266), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(KEYINPUT74), .A3(new_n274), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n274), .B1(new_n273), .B2(new_n277), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n265), .A2(KEYINPUT73), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g085(.A(new_n281), .B(new_n286), .C1(new_n255), .C2(new_n258), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n206), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n207), .B1(new_n227), .B2(new_n251), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n216), .B1(new_n243), .B2(KEYINPUT27), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(new_n209), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n225), .B1(new_n292), .B2(new_n212), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n239), .A2(new_n241), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n222), .B(new_n233), .C1(new_n294), .C2(new_n248), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n295), .A2(new_n246), .B1(new_n238), .B2(new_n244), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT75), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n227), .A2(new_n251), .A3(new_n252), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n207), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n289), .B1(new_n301), .B2(KEYINPUT76), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n303), .A3(new_n207), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n279), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n205), .B1(new_n288), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(KEYINPUT76), .ZN(new_n307));
  INV_X1    g106(.A(new_n289), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n286), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n297), .A2(new_n299), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n311), .A2(new_n208), .B1(new_n256), .B2(new_n257), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n281), .B1(new_n312), .B2(new_n286), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n259), .A2(KEYINPUT77), .A3(new_n279), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n206), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT38), .B1(new_n306), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT38), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n286), .B1(new_n302), .B2(new_n304), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n206), .B1(new_n259), .B2(new_n286), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT90), .B1(new_n306), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n205), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n310), .A2(new_n315), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G225gat), .A2(G233gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n327));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT2), .ZN(new_n329));
  OR2_X1    g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT79), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT80), .B(G162gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(G155gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G155gat), .B(G162gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n330), .A3(new_n331), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n345));
  INV_X1    g144(.A(G127gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G134gat), .ZN(new_n347));
  INV_X1    g146(.A(G134gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G127gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT68), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G113gat), .B(G120gat), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n351), .B(new_n352), .C1(KEYINPUT1), .C2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G120gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G113gat), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G120gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G127gat), .B(G134gat), .ZN(new_n361));
  AND2_X1   g160(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n362));
  NOR2_X1   g161(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n360), .A2(new_n361), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n354), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n338), .B(new_n368), .C1(new_n341), .C2(new_n343), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n345), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT81), .B1(new_n344), .B2(KEYINPUT3), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n326), .B(new_n327), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n344), .A2(new_n367), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT4), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n354), .A2(new_n366), .ZN(new_n376));
  AND2_X1   g175(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n378));
  OAI21_X1  g177(.A(G155gat), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT2), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n330), .A2(new_n331), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n333), .A2(new_n334), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n336), .B1(new_n342), .B2(KEYINPUT79), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n380), .A2(new_n383), .B1(new_n384), .B2(new_n332), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT82), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n376), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT82), .B1(new_n344), .B2(new_n367), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n375), .B1(new_n389), .B2(KEYINPUT4), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n369), .A2(new_n367), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n385), .B2(new_n368), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n394), .A3(new_n345), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n388), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n374), .A2(KEYINPUT4), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n395), .A2(new_n397), .A3(new_n326), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n344), .A2(new_n367), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n387), .A2(new_n388), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n326), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n327), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n391), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n404), .A3(new_n409), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n373), .A2(new_n390), .B1(new_n399), .B2(new_n403), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(new_n409), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT6), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n325), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT37), .B1(new_n313), .B2(new_n314), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n324), .B1(new_n419), .B2(new_n310), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n309), .A2(new_n279), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT38), .B1(new_n421), .B2(new_n320), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n317), .A2(new_n323), .A3(new_n418), .A4(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G78gat), .B(G106gat), .Z(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT85), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G22gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT3), .B1(new_n279), .B2(new_n298), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT86), .B1(new_n432), .B2(new_n385), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n282), .A2(new_n283), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n284), .A2(new_n285), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT29), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n434), .B(new_n344), .C1(new_n437), .C2(KEYINPUT3), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n369), .A2(new_n298), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n286), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G228gat), .ZN(new_n442));
  INV_X1    g241(.A(G233gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n273), .A2(new_n274), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n282), .B2(new_n283), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n368), .B1(new_n447), .B2(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n344), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n439), .B2(new_n286), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n431), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n430), .B(new_n451), .C1(new_n441), .C2(new_n444), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n429), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n444), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n344), .B1(new_n437), .B2(KEYINPUT3), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n457), .A2(KEYINPUT86), .B1(new_n286), .B2(new_n439), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n458), .B2(new_n438), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n430), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n452), .A3(new_n431), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n428), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n387), .A2(new_n388), .A3(new_n326), .A4(new_n400), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT89), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n390), .A2(new_n395), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT39), .B(new_n466), .C1(new_n467), .C2(new_n326), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n326), .B1(new_n390), .B2(new_n395), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n410), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n468), .A2(KEYINPUT40), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT40), .B1(new_n468), .B2(new_n471), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n472), .A2(new_n473), .A3(new_n416), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n310), .A2(KEYINPUT30), .A3(new_n315), .A4(new_n324), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n280), .A2(new_n287), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n205), .B1(new_n476), .B2(new_n305), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n309), .A2(new_n286), .B1(new_n313), .B2(new_n314), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT30), .B1(new_n479), .B2(new_n324), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n425), .A2(new_n464), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n256), .A2(new_n376), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n227), .A2(new_n251), .A3(new_n367), .ZN(new_n485));
  NAND2_X1  g284(.A1(G227gat), .A2(G233gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT64), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT32), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G71gat), .B(G99gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT72), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G15gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G43gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n484), .A2(new_n485), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n486), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT34), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n487), .A2(KEYINPUT34), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT32), .B(new_n488), .C1(new_n495), .C2(new_n490), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n497), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n497), .A2(new_n503), .B1(new_n502), .B2(new_n500), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n483), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(KEYINPUT36), .A3(new_n504), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n412), .B1(new_n415), .B2(new_n409), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n391), .A2(new_n404), .A3(new_n409), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT84), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT84), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n411), .A2(new_n514), .A3(new_n412), .A4(new_n413), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n417), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n325), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n516), .A2(new_n518), .A3(new_n475), .A4(new_n477), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n455), .A2(KEYINPUT87), .A3(new_n462), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT87), .B1(new_n455), .B2(new_n462), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n510), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n504), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n463), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT35), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n478), .A2(new_n480), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT91), .B(KEYINPUT35), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n414), .B2(new_n417), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n482), .A2(new_n523), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n533));
  NAND2_X1  g332(.A1(G29gat), .A2(G36gat), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT94), .B1(G29gat), .B2(G36gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(G43gat), .B(G50gat), .ZN(new_n536));
  OAI221_X1 g335(.A(new_n534), .B1(KEYINPUT14), .B2(new_n535), .C1(new_n536), .C2(KEYINPUT15), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n536), .A2(KEYINPUT15), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(KEYINPUT14), .ZN(new_n539));
  NOR3_X1   g338(.A1(KEYINPUT94), .A2(G29gat), .A3(G36gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT15), .B(new_n536), .C1(new_n537), .C2(new_n541), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G8gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT16), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(G1gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(G1gat), .B2(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI221_X1 g351(.A(new_n548), .B1(new_n549), .B2(new_n545), .C1(G1gat), .C2(new_n546), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n544), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n542), .A2(new_n543), .B1(new_n553), .B2(new_n552), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n558), .B(KEYINPUT13), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n533), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(KEYINPUT96), .B(new_n559), .C1(new_n555), .C2(new_n556), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n544), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n554), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n542), .A2(KEYINPUT17), .A3(new_n543), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n556), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n558), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n568), .A2(KEYINPUT18), .A3(new_n558), .A4(new_n569), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n563), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G197gat), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT11), .B(G169gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT92), .B(KEYINPUT12), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n574), .A2(KEYINPUT93), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n574), .B2(KEYINPUT93), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n532), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT98), .ZN(new_n588));
  NAND2_X1  g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT97), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G57gat), .B(G64gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT99), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT9), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT100), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n591), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G71gat), .ZN(new_n598));
  INV_X1    g397(.A(G78gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n592), .B1(new_n589), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n346), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n346), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n586), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  INV_X1    g413(.A(new_n586), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n554), .B1(new_n604), .B2(KEYINPUT21), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT101), .Z(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n620));
  INV_X1    g419(.A(G155gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n613), .A2(new_n616), .A3(new_n623), .A4(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G85gat), .A2(G92gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g431(.A1(G99gat), .A2(G106gat), .ZN(new_n633));
  INV_X1    g432(.A(G85gat), .ZN(new_n634));
  INV_X1    g433(.A(G92gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(KEYINPUT8), .A2(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G99gat), .B(G106gat), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(new_n640), .A3(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n543), .B2(new_n542), .ZN(new_n643));
  AND3_X1   g442(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT103), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n565), .A2(new_n567), .A3(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G190gat), .B(G218gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  INV_X1    g453(.A(new_n648), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n643), .A2(new_n647), .A3(new_n644), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n654), .B(new_n650), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n653), .A2(KEYINPUT105), .A3(new_n657), .A4(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n661), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n654), .B1(new_n649), .B2(new_n650), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n668), .A3(new_n657), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n649), .A2(KEYINPUT104), .A3(new_n654), .A4(new_n650), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n660), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n593), .A2(new_n596), .ZN(new_n673));
  INV_X1    g472(.A(new_n591), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n675), .A2(new_n602), .A3(new_n641), .A4(new_n639), .ZN(new_n676));
  INV_X1    g475(.A(new_n641), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n640), .B1(new_n632), .B2(new_n636), .ZN(new_n678));
  OAI22_X1  g477(.A1(new_n597), .A2(new_n603), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G230gat), .A2(G233gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT10), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n676), .A2(new_n684), .A3(new_n679), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n641), .A4(new_n639), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n681), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n691), .B(new_n692), .Z(new_n693));
  AOI21_X1  g492(.A(new_n682), .B1(new_n685), .B2(new_n686), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT106), .ZN(new_n695));
  AND4_X1   g494(.A1(new_n683), .A2(new_n690), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n693), .B1(new_n688), .B2(new_n683), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n629), .A2(new_n672), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n585), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n516), .B(KEYINPUT107), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g504(.A1(new_n701), .A2(new_n528), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n545), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT108), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT16), .B(G8gat), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT42), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(G1325gat));
  INV_X1    g511(.A(new_n510), .ZN(new_n713));
  OAI21_X1  g512(.A(G15gat), .B1(new_n701), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n524), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n701), .B2(new_n715), .ZN(G1326gat));
  INV_X1    g515(.A(new_n522), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT43), .B(G22gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  NAND3_X1  g519(.A1(new_n629), .A2(new_n672), .A3(new_n698), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n585), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n723), .A2(G29gat), .A3(new_n703), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT45), .Z(new_n725));
  INV_X1    g524(.A(new_n672), .ZN(new_n726));
  AND4_X1   g525(.A1(new_n317), .A2(new_n323), .A3(new_n418), .A4(new_n424), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n481), .A2(new_n464), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n523), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n527), .A2(new_n531), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n532), .B2(new_n726), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n628), .A2(new_n584), .A3(new_n699), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT110), .B1(new_n737), .B2(new_n703), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G29gat), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n737), .A2(KEYINPUT110), .A3(new_n703), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n725), .B1(new_n739), .B2(new_n740), .ZN(G1328gat));
  NOR3_X1   g540(.A1(new_n723), .A2(G36gat), .A3(new_n528), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT46), .ZN(new_n743));
  OAI21_X1  g542(.A(G36gat), .B1(new_n737), .B2(new_n528), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1329gat));
  INV_X1    g544(.A(G43gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n723), .B2(new_n524), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n713), .A2(new_n746), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n737), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g550(.A(new_n723), .ZN(new_n752));
  AOI211_X1 g551(.A(G50gat), .B(new_n717), .C1(new_n752), .C2(KEYINPUT111), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G50gat), .B1(new_n737), .B2(new_n464), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(KEYINPUT48), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n735), .A2(new_n522), .A3(new_n736), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n753), .A2(new_n754), .B1(G50gat), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(KEYINPUT48), .B2(new_n759), .ZN(G1331gat));
  NAND2_X1  g559(.A1(new_n729), .A2(new_n730), .ZN(new_n761));
  NOR4_X1   g560(.A1(new_n629), .A2(new_n672), .A3(new_n583), .A4(new_n698), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n702), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g565(.A1(new_n528), .A2(KEYINPUT112), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n528), .A2(KEYINPUT112), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  AND2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n771), .B2(new_n772), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n763), .B2(new_n713), .ZN(new_n776));
  INV_X1    g575(.A(new_n524), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n598), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n763), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n717), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(new_n599), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n628), .A2(new_n583), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n698), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n735), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n703), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788));
  AOI211_X1 g587(.A(new_n788), .B(KEYINPUT51), .C1(new_n731), .C2(new_n783), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n761), .A2(new_n672), .A3(new_n783), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT114), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n532), .A2(new_n726), .A3(new_n784), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n761), .A2(KEYINPUT51), .A3(new_n672), .A4(new_n783), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n702), .A2(new_n634), .A3(new_n699), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n787), .B1(new_n800), .B2(new_n801), .ZN(G1336gat));
  XNOR2_X1  g601(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n735), .A2(new_n769), .A3(new_n785), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(G92gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n769), .A2(new_n635), .A3(new_n699), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n791), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n808), .B2(new_n796), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT115), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n528), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n732), .A2(new_n734), .A3(new_n812), .A4(new_n785), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G92gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n809), .B2(KEYINPUT115), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT52), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n807), .A2(new_n816), .ZN(G1337gat));
  OAI21_X1  g616(.A(G99gat), .B1(new_n786), .B2(new_n713), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n698), .A2(new_n524), .A3(G99gat), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n800), .B2(new_n819), .ZN(G1338gat));
  NAND4_X1  g619(.A1(new_n732), .A2(new_n734), .A3(new_n522), .A4(new_n785), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G106gat), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n808), .A2(new_n796), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n464), .A2(new_n698), .A3(G106gat), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n796), .B(KEYINPUT113), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n788), .B1(new_n794), .B2(KEYINPUT51), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n790), .A2(KEYINPUT114), .A3(new_n791), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n825), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n732), .A2(new_n734), .A3(new_n463), .A4(new_n785), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G106gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n832), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n824), .B1(new_n793), .B2(new_n799), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n834), .B2(G106gat), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT117), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n827), .B1(new_n838), .B2(new_n841), .ZN(G1339gat));
  NAND3_X1  g641(.A1(new_n685), .A2(new_n686), .A3(new_n682), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n690), .A2(new_n844), .A3(new_n695), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n693), .B1(new_n694), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n847), .A3(KEYINPUT55), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n845), .A2(new_n847), .A3(KEYINPUT118), .A4(KEYINPUT55), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n696), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  INV_X1    g652(.A(new_n845), .ZN(new_n854));
  INV_X1    g653(.A(new_n847), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n583), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n557), .A2(new_n560), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT119), .Z(new_n859));
  AOI21_X1  g658(.A(new_n558), .B1(new_n568), .B2(new_n569), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n578), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n563), .A2(new_n572), .A3(new_n573), .A4(new_n580), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n699), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n672), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  AND4_X1   g664(.A1(new_n672), .A2(new_n852), .A3(new_n863), .A4(new_n856), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n629), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n726), .A2(new_n584), .A3(new_n628), .A4(new_n698), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n703), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n525), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n769), .ZN(new_n871));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n583), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n522), .B1(new_n867), .B2(new_n868), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n769), .A2(new_n524), .A3(new_n703), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n584), .A2(new_n357), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(G1340gat));
  AOI21_X1  g676(.A(G120gat), .B1(new_n871), .B2(new_n699), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n698), .A2(new_n355), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n875), .B2(new_n879), .ZN(G1341gat));
  INV_X1    g679(.A(new_n875), .ZN(new_n881));
  OAI21_X1  g680(.A(G127gat), .B1(new_n881), .B2(new_n629), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n871), .A2(new_n346), .A3(new_n628), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1342gat));
  NAND2_X1  g683(.A1(new_n672), .A2(new_n528), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n870), .A2(G134gat), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(KEYINPUT120), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n672), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT56), .B1(new_n892), .B2(G134gat), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n890), .B(new_n891), .C1(new_n893), .C2(new_n886), .ZN(G1343gat));
  NOR2_X1   g693(.A1(new_n510), .A2(new_n464), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n584), .A2(G141gat), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n869), .A2(new_n770), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n770), .A2(new_n713), .A3(new_n702), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n464), .B1(new_n867), .B2(new_n868), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n868), .ZN(new_n904));
  XNOR2_X1  g703(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n845), .B2(new_n847), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n581), .A2(new_n582), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n852), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n672), .B1(new_n909), .B2(new_n864), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n629), .B1(new_n910), .B2(new_n866), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n904), .B1(new_n911), .B2(KEYINPUT122), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n672), .A2(new_n852), .A3(new_n863), .A4(new_n856), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n852), .A2(new_n908), .B1(new_n863), .B2(new_n699), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n672), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n629), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n717), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n903), .B(new_n583), .C1(new_n918), .C2(new_n902), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n899), .B1(new_n919), .B2(G141gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(G1344gat));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n903), .B1(new_n918), .B2(new_n902), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n923), .B(G148gat), .C1(new_n924), .C2(new_n698), .ZN(new_n925));
  INV_X1    g724(.A(G148gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n717), .B1(new_n911), .B2(new_n868), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT124), .B1(new_n927), .B2(KEYINPUT57), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n904), .B1(new_n915), .B2(new_n629), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n929), .B(new_n902), .C1(new_n930), .C2(new_n717), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n901), .A2(KEYINPUT57), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n900), .A2(new_n698), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n926), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n925), .B1(new_n923), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n869), .A2(new_n895), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(new_n769), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n926), .A3(new_n699), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(G1345gat));
  OAI21_X1  g739(.A(G155gat), .B1(new_n924), .B2(new_n629), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n621), .A3(new_n628), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n941), .A2(KEYINPUT125), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1346gat));
  OAI21_X1  g746(.A(new_n340), .B1(new_n924), .B2(new_n726), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n885), .A2(new_n340), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n937), .B2(new_n949), .ZN(G1347gat));
  AOI21_X1  g749(.A(new_n702), .B1(new_n867), .B2(new_n868), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(new_n525), .A3(new_n769), .ZN(new_n952));
  AOI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n583), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n702), .A2(new_n528), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n873), .A2(new_n777), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n584), .A2(new_n229), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1348gat));
  NAND3_X1  g756(.A1(new_n952), .A2(new_n230), .A3(new_n699), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n955), .A2(new_n699), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n230), .ZN(G1349gat));
  AND2_X1   g759(.A1(new_n628), .A2(new_n211), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n952), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n955), .A2(new_n628), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n243), .B2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT60), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n963), .A2(new_n243), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT60), .B1(new_n967), .B2(new_n962), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n210), .A3(new_n672), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n672), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G190gat), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(G1351gat));
  AND2_X1   g774(.A1(new_n769), .A2(new_n895), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n951), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n269), .B1(new_n977), .B2(new_n584), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n954), .A2(new_n713), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n933), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n583), .A2(G197gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g784(.A(KEYINPUT126), .B(new_n978), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1352gat));
  NAND4_X1  g786(.A1(new_n951), .A2(new_n270), .A3(new_n699), .A4(new_n976), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n989), .A2(KEYINPUT62), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT62), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(G204gat), .B1(new_n981), .B2(new_n698), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1353gat));
  OR3_X1    g794(.A1(new_n977), .A2(G211gat), .A3(new_n629), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n933), .A2(new_n628), .A3(new_n980), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n997), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT63), .B1(new_n997), .B2(G211gat), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(G1354gat));
  OAI21_X1  g799(.A(G218gat), .B1(new_n981), .B2(new_n726), .ZN(new_n1001));
  OR2_X1    g800(.A1(new_n726), .A2(G218gat), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1001), .B1(new_n977), .B2(new_n1002), .ZN(G1355gat));
endmodule


