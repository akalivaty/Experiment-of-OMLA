//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n445, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  OR4_X1    g030(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(new_n460), .B2(new_n461), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AND4_X1   g047(.A1(G137), .A2(new_n470), .A3(new_n472), .A4(new_n464), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT69), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n468), .A2(new_n473), .A3(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n465), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n470), .A2(new_n472), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n464), .ZN(new_n487));
  AND2_X1   g062(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n464), .A2(KEYINPUT71), .A3(KEYINPUT4), .A4(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(new_n465), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n464), .B2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(G2104), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n491), .A2(new_n495), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT72), .Z(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n504), .A2(new_n505), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n510), .A2(new_n517), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(new_n508), .A2(G51), .ZN(new_n524));
  AND3_X1   g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(G89), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n524), .B1(KEYINPUT7), .B2(new_n525), .C1(new_n519), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n514), .A2(G63), .ZN(new_n528));
  NAND3_X1  g103(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n516), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G168));
  XNOR2_X1  g107(.A(KEYINPUT75), .B(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n518), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n519), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT74), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n538), .B2(G651), .ZN(G171));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n519), .A2(new_n540), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  AOI22_X1  g126(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n516), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n520), .A2(G91), .ZN(new_n554));
  OAI211_X1 g129(.A(G53), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(G299));
  INV_X1    g132(.A(G171), .ZN(G301));
  NAND2_X1  g133(.A1(new_n531), .A2(KEYINPUT76), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n527), .A2(KEYINPUT76), .A3(new_n530), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(G286));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  INV_X1    g137(.A(G49), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n534), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n508), .A2(KEYINPUT77), .A3(G49), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n520), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n570));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n519), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n514), .A2(new_n518), .A3(KEYINPUT78), .A4(G86), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n511), .A2(new_n513), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n508), .B2(G48), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n574), .A2(new_n579), .ZN(G305));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  XNOR2_X1  g156(.A(KEYINPUT79), .B(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n519), .A2(new_n581), .B1(new_n534), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n516), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND3_X1  g162(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n519), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(G54), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n516), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n599), .B2(G171), .ZN(G284));
  OAI21_X1  g176(.A(new_n600), .B1(new_n599), .B2(G171), .ZN(G321));
  NAND2_X1  g177(.A1(G299), .A2(new_n599), .ZN(new_n603));
  INV_X1    g178(.A(G286), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n599), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n599), .ZN(G280));
  INV_X1    g181(.A(new_n598), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g188(.A1(new_n469), .A2(G2105), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n465), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT13), .Z(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G2100), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n617), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n478), .A2(G123), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n481), .A2(G135), .ZN(new_n622));
  NOR2_X1   g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  OAI211_X1 g201(.A(new_n620), .B(new_n626), .C1(new_n618), .C2(G2100), .ZN(G156));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT15), .B(G2435), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT83), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n634), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT82), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n638), .A2(new_n641), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n629), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  AOI21_X1  g220(.A(KEYINPUT84), .B1(new_n645), .B2(new_n628), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n647));
  NOR4_X1   g222(.A1(new_n642), .A2(new_n643), .A3(new_n647), .A4(new_n629), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n644), .B(G14), .C1(new_n646), .C2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT85), .Z(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT86), .Z(new_n657));
  INV_X1    g232(.A(new_n654), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n655), .B(KEYINPUT17), .Z(new_n659));
  OAI21_X1  g234(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n654), .A2(new_n655), .A3(new_n651), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n659), .A3(new_n651), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT87), .B(G2096), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  AND3_X1   g251(.A1(new_n671), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(KEYINPUT89), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(new_n670), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT90), .Z(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n680), .B2(KEYINPUT20), .ZN(new_n681));
  OAI221_X1 g256(.A(new_n681), .B1(KEYINPUT20), .B2(new_n680), .C1(new_n675), .C2(new_n671), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G35), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G162), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT29), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G2090), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT31), .B(G11), .Z(new_n696));
  INV_X1    g271(.A(KEYINPUT24), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n691), .B1(new_n697), .B2(G34), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT101), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(G34), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(KEYINPUT101), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G160), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n691), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT102), .B(G2084), .Z(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT30), .B(G28), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(new_n691), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n625), .B2(new_n691), .ZN(new_n709));
  NOR4_X1   g284(.A1(new_n695), .A2(new_n696), .A3(new_n706), .A4(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G21), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G168), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G27), .A2(G29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G164), .B2(G29), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G2078), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n478), .A2(G129), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n614), .A2(G105), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n481), .A2(G141), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND4_X1  g298(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G29), .B2(G32), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n727), .A2(new_n728), .B1(new_n704), .B2(new_n705), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G19), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n545), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT98), .B(G1341), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n718), .B(new_n730), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n711), .A2(G20), .ZN(new_n737));
  INV_X1    g312(.A(G299), .ZN(new_n738));
  OAI211_X1 g313(.A(KEYINPUT23), .B(new_n737), .C1(new_n738), .C2(new_n711), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(KEYINPUT23), .B2(new_n737), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1956), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n710), .A2(new_n715), .A3(new_n736), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n733), .A2(new_n735), .ZN(new_n743));
  OR2_X1    g318(.A1(G29), .A2(G33), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(new_n464), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n614), .A2(G103), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G139), .ZN(new_n750));
  INV_X1    g325(.A(new_n481), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(KEYINPUT100), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(KEYINPUT100), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n744), .B1(new_n755), .B2(new_n691), .ZN(new_n756));
  INV_X1    g331(.A(G2072), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NAND2_X1  g334(.A1(G171), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G5), .B2(G16), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n759), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n691), .A2(G26), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n478), .A2(G128), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n481), .A2(G140), .ZN(new_n766));
  OR3_X1    g341(.A1(KEYINPUT99), .A2(G104), .A3(G2105), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n464), .A2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(KEYINPUT99), .B1(G104), .B2(G2105), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n767), .A2(new_n768), .A3(G2104), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n765), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n764), .B1(new_n772), .B2(new_n691), .ZN(new_n773));
  MUX2_X1   g348(.A(new_n764), .B(new_n773), .S(KEYINPUT28), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2067), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n756), .B2(new_n757), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n607), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G4), .B2(G16), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT97), .B(G1348), .Z(new_n779));
  AOI21_X1  g354(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n763), .B(new_n780), .C1(G2067), .C2(new_n774), .ZN(new_n781));
  OR3_X1    g356(.A1(new_n742), .A2(new_n743), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n691), .A2(G25), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n481), .A2(G131), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT92), .ZN(new_n785));
  OR2_X1    g360(.A1(G95), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT93), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n478), .A2(G119), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n785), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n783), .B1(new_n792), .B2(new_n691), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT35), .B(G1991), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n711), .A2(G24), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n586), .B2(new_n711), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G1986), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT96), .B1(new_n801), .B2(G16), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n801), .A2(KEYINPUT96), .A3(G16), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n802), .B(new_n803), .C1(G166), .C2(new_n711), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n711), .A2(G6), .ZN(new_n807));
  INV_X1    g382(.A(G305), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n711), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT32), .B(G1981), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n711), .A2(G23), .ZN(new_n812));
  INV_X1    g387(.A(G288), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n711), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1976), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n806), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n795), .B(new_n800), .C1(new_n818), .C2(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n798), .A2(G1986), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n819), .A2(new_n824), .A3(new_n820), .A4(new_n821), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n782), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n778), .A2(new_n779), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n827), .ZN(G150));
  NAND2_X1  g404(.A1(new_n508), .A2(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OAI221_X1 g407(.A(new_n830), .B1(new_n519), .B2(new_n831), .C1(new_n832), .C2(new_n516), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n607), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n545), .A2(new_n833), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n545), .A2(new_n833), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n837), .B(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n835), .B1(new_n842), .B2(G860), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT103), .ZN(G145));
  XNOR2_X1  g419(.A(new_n485), .B(KEYINPUT104), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n625), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G160), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n478), .A2(G130), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n481), .A2(G142), .ZN(new_n849));
  NOR2_X1   g424(.A1(G106), .A2(G2105), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n616), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n792), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n755), .A2(G164), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n502), .B(new_n746), .C1(new_n753), .C2(new_n754), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n771), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n771), .A3(new_n857), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n725), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n862), .A2(new_n858), .A3(new_n724), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n855), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n724), .B1(new_n862), .B2(new_n858), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(new_n725), .A3(new_n860), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n854), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n847), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(G37), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g446(.A(KEYINPUT105), .B(new_n855), .C1(new_n861), .C2(new_n863), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n871), .A2(new_n867), .A3(new_n847), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g450(.A(new_n610), .B(new_n840), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n598), .B1(new_n878), .B2(new_n738), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n738), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n598), .A2(KEYINPUT106), .A3(G299), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n885), .A3(new_n881), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n877), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n880), .A2(KEYINPUT107), .A3(new_n881), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n876), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT109), .ZN(new_n894));
  NAND2_X1  g469(.A1(G288), .A2(new_n586), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(G288), .A2(new_n586), .ZN(new_n897));
  OAI21_X1  g472(.A(G166), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(G303), .A3(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G305), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n808), .A3(new_n900), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n894), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n894), .A3(new_n903), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT42), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n909), .A3(new_n904), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n893), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n908), .B2(new_n904), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n905), .A2(KEYINPUT42), .A3(new_n906), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n892), .A4(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n915), .A3(new_n892), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT110), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n893), .B(KEYINPUT111), .C1(new_n910), .C2(new_n907), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n913), .A2(new_n917), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(G868), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n833), .A2(new_n599), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT115), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n880), .A2(KEYINPUT107), .A3(new_n881), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT107), .B1(new_n880), .B2(new_n881), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G286), .A2(G171), .ZN(new_n930));
  INV_X1    g505(.A(new_n840), .ZN(new_n931));
  NOR2_X1   g506(.A1(G171), .A2(new_n531), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G301), .B1(new_n559), .B2(new_n560), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n840), .B1(new_n935), .B2(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n926), .B1(new_n929), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n889), .A2(new_n890), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n939), .A2(KEYINPUT115), .A3(new_n936), .A4(new_n934), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n941));
  INV_X1    g516(.A(new_n883), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n880), .A2(new_n881), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(KEYINPUT114), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n936), .A2(KEYINPUT112), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT112), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n943), .A2(KEYINPUT114), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n938), .B(new_n940), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n902), .A2(new_n903), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n902), .A2(KEYINPUT113), .A3(new_n903), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n882), .B1(new_n945), .B2(new_n946), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n884), .A2(new_n886), .B1(new_n934), .B2(new_n936), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n958), .B2(new_n950), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n955), .A2(new_n959), .A3(KEYINPUT43), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n953), .B(new_n952), .C1(new_n956), .C2(new_n957), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT43), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT44), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n955), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n959), .B2(new_n961), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(G397));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n502), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G125), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n467), .B1(new_n480), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G2105), .ZN(new_n976));
  INV_X1    g551(.A(new_n475), .ZN(new_n977));
  INV_X1    g552(.A(new_n473), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .A4(G40), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n973), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT116), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n982), .A2(G1986), .A3(G290), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n984));
  XNOR2_X1  g559(.A(new_n983), .B(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n792), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n794), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n724), .B(G1996), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n771), .B(G2067), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n986), .A2(new_n794), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n985), .B1(new_n981), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n982), .B2(G1996), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n981), .B1(new_n724), .B2(new_n990), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n981), .A2(KEYINPUT46), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT47), .Z(new_n1001));
  NAND2_X1  g576(.A1(new_n987), .A2(new_n991), .ZN(new_n1002));
  INV_X1    g577(.A(G2067), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n772), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n982), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n994), .A2(new_n1001), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(G305), .B2(G1981), .ZN(new_n1008));
  INV_X1    g583(.A(G1981), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n574), .A2(KEYINPUT118), .A3(new_n1009), .A4(new_n579), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n579), .B1(new_n571), .B2(new_n519), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1008), .A2(new_n1010), .B1(G1981), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT49), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n979), .A2(new_n971), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1011), .A2(G1981), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT119), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1012), .A2(new_n1022), .A3(KEYINPUT49), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1013), .B(new_n1016), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1016), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n813), .A2(G1976), .ZN(new_n1028));
  OR3_X1    g603(.A1(new_n1026), .A2(new_n1028), .A3(KEYINPUT52), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G303), .A2(G8), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n1032));
  XNOR2_X1  g607(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g609(.A(G40), .ZN(new_n1035));
  NOR4_X1   g610(.A1(new_n468), .A2(new_n475), .A3(new_n1035), .A4(new_n473), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n502), .A2(new_n1037), .A3(new_n970), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1039), .A2(G2090), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT45), .B1(new_n502), .B2(new_n970), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n979), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n805), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1015), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1033), .A2(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1030), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1024), .A2(new_n1025), .A3(new_n813), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1017), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1016), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(KEYINPUT120), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1041), .B2(new_n979), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1043), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n714), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(G2084), .B2(new_n1039), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AND4_X1   g634(.A1(new_n1059), .A2(new_n1024), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n604), .B1(new_n1033), .B2(new_n1046), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT63), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NOR4_X1   g639(.A1(new_n1030), .A2(new_n1061), .A3(new_n1064), .A4(new_n1058), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1048), .B(new_n1051), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n973), .A2(new_n1036), .A3(new_n1043), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT121), .ZN(new_n1069));
  INV_X1    g644(.A(G1956), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1039), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1042), .A2(new_n1072), .A3(new_n1043), .A4(new_n1067), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(G299), .B(KEYINPUT57), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1348), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1039), .A2(new_n1077), .B1(new_n1003), .B2(new_n1014), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n598), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  XNOR2_X1  g655(.A(G299), .B(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(new_n1069), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n973), .A2(new_n1036), .A3(new_n998), .A4(new_n1043), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT58), .B(G1341), .Z(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n979), .B2(new_n971), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT122), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1089), .A3(new_n1086), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1090), .A3(new_n545), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT59), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1088), .A2(new_n1090), .A3(new_n1093), .A4(new_n545), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1078), .B1(KEYINPUT60), .B2(new_n607), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(new_n598), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1078), .A2(KEYINPUT60), .A3(new_n607), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1095), .A2(new_n1098), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1076), .A2(KEYINPUT61), .A3(new_n1082), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1076), .A2(KEYINPUT123), .A3(new_n1082), .A4(KEYINPUT61), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1083), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT124), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1039), .A2(G2084), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n531), .B(new_n1112), .C1(new_n1055), .C2(new_n714), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT125), .B(KEYINPUT51), .C1(new_n1113), .C2(new_n1015), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1056), .B(G168), .C1(G2084), .C2(new_n1039), .ZN(new_n1115));
  OR2_X1    g690(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1116));
  NAND2_X1  g691(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1115), .A2(G8), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1057), .A2(G8), .A3(new_n531), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1114), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(G171), .B(KEYINPUT54), .ZN(new_n1121));
  INV_X1    g696(.A(G2078), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1042), .A2(new_n1122), .A3(new_n1043), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT126), .B(KEYINPUT53), .Z(new_n1124));
  AOI22_X1  g699(.A1(new_n1123), .A2(new_n1124), .B1(new_n759), .B2(new_n1039), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1121), .B(new_n1125), .C1(new_n1126), .C2(new_n1123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(KEYINPUT53), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1055), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1121), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1120), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n1083), .C1(new_n1104), .C2(new_n1109), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1111), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1120), .A2(KEYINPUT62), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1120), .A2(KEYINPUT62), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(G171), .A3(new_n1129), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1033), .A2(new_n1046), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1047), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1030), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1066), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n993), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n586), .B(G1986), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n982), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1006), .B1(new_n1143), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g722(.A1(new_n958), .A2(new_n950), .ZN(new_n1149));
  INV_X1    g723(.A(G37), .ZN(new_n1150));
  NAND3_X1  g724(.A1(new_n1149), .A2(new_n961), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g725(.A1(new_n1151), .A2(KEYINPUT43), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n955), .A2(new_n959), .A3(new_n965), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n649), .A2(G319), .ZN(new_n1155));
  AOI211_X1 g729(.A(G227), .B(new_n1155), .C1(new_n869), .C2(new_n873), .ZN(new_n1156));
  AND3_X1   g730(.A1(new_n1154), .A2(new_n689), .A3(new_n1156), .ZN(G308));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n689), .A3(new_n1156), .ZN(G225));
endmodule


