

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U326 ( .A(n305), .B(n304), .ZN(n313) );
  XNOR2_X1 U327 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n365) );
  XNOR2_X1 U328 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U329 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n393) );
  XNOR2_X1 U330 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U331 ( .A(n394), .B(n393), .ZN(n573) );
  XNOR2_X1 U332 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U333 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n295) );
  XNOR2_X1 U335 ( .A(G71GAT), .B(G78GAT), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U337 ( .A(G57GAT), .B(n296), .Z(n332) );
  XOR2_X1 U338 ( .A(G204GAT), .B(KEYINPUT76), .Z(n318) );
  XNOR2_X1 U339 ( .A(n318), .B(G64GAT), .ZN(n298) );
  XOR2_X1 U340 ( .A(G120GAT), .B(G148GAT), .Z(n400) );
  XNOR2_X1 U341 ( .A(G176GAT), .B(n400), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n332), .B(n299), .ZN(n305) );
  XOR2_X1 U344 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n301) );
  XNOR2_X1 U345 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n300) );
  XOR2_X1 U346 ( .A(n301), .B(n300), .Z(n303) );
  NAND2_X1 U347 ( .A1(G230GAT), .A2(G233GAT), .ZN(n302) );
  XOR2_X1 U348 ( .A(KEYINPUT74), .B(G92GAT), .Z(n307) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .ZN(n306) );
  XNOR2_X1 U350 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U351 ( .A(G106GAT), .B(n308), .Z(n375) );
  XOR2_X1 U352 ( .A(KEYINPUT77), .B(KEYINPUT72), .Z(n310) );
  XNOR2_X1 U353 ( .A(KEYINPUT78), .B(KEYINPUT75), .ZN(n309) );
  XNOR2_X1 U354 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U355 ( .A(n375), .B(n311), .ZN(n312) );
  XNOR2_X1 U356 ( .A(n313), .B(n312), .ZN(n387) );
  XNOR2_X1 U357 ( .A(KEYINPUT41), .B(n387), .ZN(n546) );
  INV_X1 U358 ( .A(n546), .ZN(n531) );
  XOR2_X1 U359 ( .A(G92GAT), .B(G218GAT), .Z(n315) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n327) );
  XOR2_X1 U362 ( .A(G64GAT), .B(KEYINPUT82), .Z(n317) );
  XNOR2_X1 U363 ( .A(G8GAT), .B(G211GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n336) );
  XOR2_X1 U365 ( .A(n318), .B(n336), .Z(n320) );
  NAND2_X1 U366 ( .A1(G226GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U368 ( .A(n321), .B(KEYINPUT96), .Z(n325) );
  XOR2_X1 U369 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n323) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n418) );
  XNOR2_X1 U372 ( .A(G183GAT), .B(n418), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U375 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n329) );
  XNOR2_X1 U376 ( .A(KEYINPUT17), .B(G176GAT), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U378 ( .A(G169GAT), .B(n330), .ZN(n450) );
  XNOR2_X1 U379 ( .A(n331), .B(n450), .ZN(n514) );
  XOR2_X1 U380 ( .A(KEYINPUT14), .B(KEYINPUT83), .Z(n334) );
  XNOR2_X1 U381 ( .A(G1GAT), .B(KEYINPUT84), .ZN(n333) );
  XNOR2_X1 U382 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U383 ( .A(n332), .B(n335), .ZN(n344) );
  XOR2_X1 U384 ( .A(G22GAT), .B(G155GAT), .Z(n423) );
  XOR2_X1 U385 ( .A(n336), .B(n423), .Z(n338) );
  NAND2_X1 U386 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U388 ( .A(n339), .B(KEYINPUT12), .Z(n342) );
  XNOR2_X1 U389 ( .A(G15GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U390 ( .A(n340), .B(G127GAT), .ZN(n442) );
  XNOR2_X1 U391 ( .A(n442), .B(KEYINPUT15), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U393 ( .A(n344), .B(n343), .ZN(n551) );
  XNOR2_X1 U394 ( .A(KEYINPUT108), .B(n551), .ZN(n564) );
  XNOR2_X1 U395 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n345), .B(G29GAT), .ZN(n347) );
  INV_X1 U397 ( .A(KEYINPUT8), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n349) );
  XNOR2_X1 U399 ( .A(G43GAT), .B(G50GAT), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n379) );
  XNOR2_X1 U401 ( .A(G141GAT), .B(G113GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n350), .B(G1GAT), .ZN(n395) );
  XNOR2_X1 U403 ( .A(n379), .B(n395), .ZN(n352) );
  XOR2_X1 U404 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n358) );
  XOR2_X1 U406 ( .A(KEYINPUT29), .B(G8GAT), .Z(n354) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(G15GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G197GAT), .Z(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n360) );
  NAND2_X1 U412 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U414 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n362) );
  XNOR2_X1 U415 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n364), .B(n363), .ZN(n383) );
  INV_X1 U418 ( .A(n383), .ZN(n544) );
  NAND2_X1 U419 ( .A1(n544), .A2(n546), .ZN(n366) );
  NOR2_X1 U420 ( .A1(n564), .A2(n367), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n368), .B(KEYINPUT110), .ZN(n380) );
  XOR2_X1 U422 ( .A(G218GAT), .B(G162GAT), .Z(n424) );
  XOR2_X1 U423 ( .A(n424), .B(KEYINPUT79), .Z(n370) );
  NAND2_X1 U424 ( .A1(G232GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U426 ( .A(KEYINPUT80), .B(KEYINPUT9), .Z(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(n374), .B(n373), .Z(n377) );
  XOR2_X1 U430 ( .A(G190GAT), .B(G134GAT), .Z(n438) );
  XNOR2_X1 U431 ( .A(n438), .B(n375), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n384) );
  NAND2_X1 U434 ( .A1(n380), .A2(n384), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n381), .B(KEYINPUT111), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n382), .B(KEYINPUT47), .ZN(n390) );
  XOR2_X1 U437 ( .A(KEYINPUT70), .B(n383), .Z(n523) );
  INV_X1 U438 ( .A(n384), .ZN(n555) );
  XNOR2_X1 U439 ( .A(n555), .B(KEYINPUT81), .ZN(n567) );
  XNOR2_X1 U440 ( .A(KEYINPUT36), .B(n567), .ZN(n585) );
  INV_X1 U441 ( .A(n551), .ZN(n582) );
  NOR2_X1 U442 ( .A1(n585), .A2(n582), .ZN(n385) );
  XOR2_X1 U443 ( .A(KEYINPUT45), .B(n385), .Z(n386) );
  NOR2_X1 U444 ( .A1(n523), .A2(n386), .ZN(n388) );
  NAND2_X1 U445 ( .A1(n388), .A2(n387), .ZN(n389) );
  NAND2_X1 U446 ( .A1(n390), .A2(n389), .ZN(n392) );
  XNOR2_X1 U447 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n524) );
  NAND2_X1 U449 ( .A1(n514), .A2(n524), .ZN(n394) );
  XOR2_X1 U450 ( .A(KEYINPUT0), .B(KEYINPUT86), .Z(n437) );
  XOR2_X1 U451 ( .A(n437), .B(n395), .Z(n397) );
  NAND2_X1 U452 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n405) );
  XOR2_X1 U454 ( .A(G85GAT), .B(G155GAT), .Z(n399) );
  XNOR2_X1 U455 ( .A(G127GAT), .B(G134GAT), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U457 ( .A(n401), .B(n400), .Z(n403) );
  XNOR2_X1 U458 ( .A(G29GAT), .B(G162GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n413) );
  XOR2_X1 U461 ( .A(KEYINPUT95), .B(G57GAT), .Z(n411) );
  XNOR2_X1 U462 ( .A(KEYINPUT94), .B(KEYINPUT3), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n406), .B(KEYINPUT2), .ZN(n420) );
  XOR2_X1 U464 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U465 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n420), .B(n409), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n574) );
  INV_X1 U470 ( .A(n574), .ZN(n489) );
  XOR2_X1 U471 ( .A(G204GAT), .B(G211GAT), .Z(n415) );
  XNOR2_X1 U472 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n432) );
  XOR2_X1 U474 ( .A(G148GAT), .B(G78GAT), .Z(n417) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U477 ( .A(n419), .B(n418), .Z(n422) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(n420), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n428) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U483 ( .A(n428), .B(n427), .Z(n430) );
  XNOR2_X1 U484 ( .A(G50GAT), .B(G106GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U486 ( .A(n432), .B(n431), .Z(n463) );
  NAND2_X1 U487 ( .A1(n489), .A2(n463), .ZN(n433) );
  OR2_X1 U488 ( .A1(n573), .A2(n433), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n434), .B(KEYINPUT55), .ZN(n452) );
  XOR2_X1 U490 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n436) );
  XNOR2_X1 U491 ( .A(KEYINPUT89), .B(KEYINPUT87), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n449) );
  XOR2_X1 U493 ( .A(G71GAT), .B(n437), .Z(n440) );
  XNOR2_X1 U494 ( .A(G113GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n441), .B(G99GAT), .Z(n447) );
  XOR2_X1 U497 ( .A(n442), .B(G120GAT), .Z(n444) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n516) );
  NAND2_X1 U504 ( .A1(n452), .A2(n516), .ZN(n566) );
  NOR2_X1 U505 ( .A1(n531), .A2(n566), .ZN(n455) );
  XNOR2_X1 U506 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n453) );
  XNOR2_X1 U507 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n473) );
  NAND2_X1 U508 ( .A1(n387), .A2(n523), .ZN(n487) );
  NAND2_X1 U509 ( .A1(n516), .A2(n514), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n463), .A2(n456), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT25), .ZN(n460) );
  XOR2_X1 U512 ( .A(KEYINPUT27), .B(n514), .Z(n462) );
  NOR2_X1 U513 ( .A1(n516), .A2(n463), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n458), .B(KEYINPUT26), .ZN(n575) );
  INV_X1 U515 ( .A(n575), .ZN(n543) );
  NOR2_X1 U516 ( .A1(n462), .A2(n543), .ZN(n459) );
  NOR2_X1 U517 ( .A1(n460), .A2(n459), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n574), .A2(n461), .ZN(n468) );
  XNOR2_X1 U519 ( .A(KEYINPUT90), .B(n516), .ZN(n466) );
  NOR2_X1 U520 ( .A1(n489), .A2(n462), .ZN(n525) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT64), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT28), .ZN(n529) );
  NAND2_X1 U523 ( .A1(n525), .A2(n529), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n483) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(KEYINPUT85), .Z(n470) );
  NAND2_X1 U527 ( .A1(n551), .A2(n567), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n471) );
  OR2_X1 U529 ( .A1(n483), .A2(n471), .ZN(n501) );
  NOR2_X1 U530 ( .A1(n487), .A2(n501), .ZN(n479) );
  NAND2_X1 U531 ( .A1(n574), .A2(n479), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(G1324GAT) );
  XOR2_X1 U533 ( .A(G8GAT), .B(KEYINPUT97), .Z(n475) );
  NAND2_X1 U534 ( .A1(n479), .A2(n514), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U537 ( .A1(n479), .A2(n516), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(n478), .ZN(G1326GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n481) );
  INV_X1 U541 ( .A(n529), .ZN(n520) );
  NAND2_X1 U542 ( .A1(n479), .A2(n520), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n551), .A2(n483), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(KEYINPUT101), .ZN(n485) );
  NOR2_X1 U547 ( .A1(n585), .A2(n485), .ZN(n486) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n486), .ZN(n510) );
  NOR2_X1 U549 ( .A1(n510), .A2(n487), .ZN(n488) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(n488), .Z(n497) );
  NOR2_X1 U551 ( .A1(n497), .A2(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  INV_X1 U554 ( .A(n514), .ZN(n492) );
  NOR2_X1 U555 ( .A1(n492), .A2(n497), .ZN(n493) );
  XOR2_X1 U556 ( .A(KEYINPUT102), .B(n493), .Z(n494) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  INV_X1 U558 ( .A(n516), .ZN(n526) );
  NOR2_X1 U559 ( .A1(n526), .A2(n497), .ZN(n495) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(n495), .Z(n496) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT103), .ZN(n499) );
  NOR2_X1 U563 ( .A1(n529), .A2(n497), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  NAND2_X1 U567 ( .A1(n546), .A2(n383), .ZN(n511) );
  NOR2_X1 U568 ( .A1(n511), .A2(n501), .ZN(n506) );
  NAND2_X1 U569 ( .A1(n574), .A2(n506), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n514), .A2(n506), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n516), .A2(n506), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n508) );
  NAND2_X1 U576 ( .A1(n506), .A2(n520), .ZN(n507) );
  XNOR2_X1 U577 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U578 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  NOR2_X1 U579 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(KEYINPUT106), .ZN(n519) );
  NAND2_X1 U581 ( .A1(n574), .A2(n519), .ZN(n513) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n514), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n515), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U585 ( .A(G99GAT), .B(KEYINPUT107), .Z(n518) );
  NAND2_X1 U586 ( .A1(n519), .A2(n516), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n518), .B(n517), .ZN(G1338GAT) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1339GAT) );
  INV_X1 U591 ( .A(n523), .ZN(n559) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n542) );
  NOR2_X1 U593 ( .A1(n526), .A2(n542), .ZN(n527) );
  XOR2_X1 U594 ( .A(KEYINPUT113), .B(n527), .Z(n528) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n538) );
  NOR2_X1 U596 ( .A1(n559), .A2(n538), .ZN(n530) );
  XOR2_X1 U597 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  NOR2_X1 U598 ( .A1(n531), .A2(n538), .ZN(n533) );
  XNOR2_X1 U599 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  INV_X1 U602 ( .A(n538), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n564), .A2(n535), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  NOR2_X1 U606 ( .A1(n567), .A2(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U609 ( .A(G134GAT), .B(n541), .Z(G1343GAT) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n544), .A2(n556), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n550) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U615 ( .A1(n556), .A2(n546), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n553) );
  NAND2_X1 U619 ( .A1(n556), .A2(n551), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(G162GAT), .B(KEYINPUT119), .Z(n558) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1347GAT) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n566), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  INV_X1 U629 ( .A(n566), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n578) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n584) );
  NOR2_X1 U641 ( .A1(n383), .A2(n584), .ZN(n577) );
  XOR2_X1 U642 ( .A(n578), .B(n577), .Z(G1352GAT) );
  NOR2_X1 U643 ( .A1(n387), .A2(n584), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G218GAT), .B(n588), .Z(G1355GAT) );
endmodule

