

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756;

  XNOR2_X1 U377 ( .A(n439), .B(n363), .ZN(n562) );
  INV_X1 U378 ( .A(G953), .ZN(n747) );
  NOR2_X1 U379 ( .A1(n579), .A2(n691), .ZN(n581) );
  NAND2_X1 U380 ( .A1(n562), .A2(n601), .ZN(n675) );
  OR2_X1 U381 ( .A1(n425), .A2(n424), .ZN(n665) );
  NOR2_X1 U382 ( .A1(n732), .A2(KEYINPUT2), .ZN(n648) );
  XNOR2_X1 U383 ( .A(n447), .B(KEYINPUT45), .ZN(n629) );
  NAND2_X1 U384 ( .A1(n559), .A2(n558), .ZN(n402) );
  NOR2_X1 U385 ( .A1(n567), .A2(KEYINPUT85), .ZN(n446) );
  XNOR2_X1 U386 ( .A(n392), .B(n565), .ZN(n568) );
  XNOR2_X1 U387 ( .A(n581), .B(n580), .ZN(n754) );
  NOR2_X1 U388 ( .A1(n544), .A2(n525), .ZN(n534) );
  XNOR2_X1 U389 ( .A(n619), .B(KEYINPUT38), .ZN(n672) );
  XNOR2_X1 U390 ( .A(n358), .B(n456), .ZN(n686) );
  NOR2_X2 U391 ( .A1(n394), .A2(n502), .ZN(n503) );
  OR2_X2 U392 ( .A1(n568), .A2(n566), .ZN(n567) );
  XNOR2_X1 U393 ( .A(G146), .B(G125), .ZN(n475) );
  NOR2_X1 U394 ( .A1(n659), .A2(n576), .ZN(n585) );
  OR2_X1 U395 ( .A1(n488), .A2(G902), .ZN(n439) );
  NAND2_X1 U396 ( .A1(n754), .A2(n753), .ZN(n374) );
  INV_X1 U397 ( .A(KEYINPUT47), .ZN(n450) );
  NOR2_X1 U398 ( .A1(G900), .A2(n571), .ZN(n572) );
  XNOR2_X1 U399 ( .A(n455), .B(KEYINPUT102), .ZN(n571) );
  OR2_X1 U400 ( .A1(n686), .A2(n570), .ZN(n455) );
  NOR2_X1 U401 ( .A1(G953), .A2(G237), .ZN(n507) );
  XNOR2_X1 U402 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n494) );
  XNOR2_X1 U403 ( .A(G122), .B(G140), .ZN(n459) );
  XOR2_X1 U404 ( .A(G131), .B(G104), .Z(n462) );
  XNOR2_X1 U405 ( .A(G143), .B(G113), .ZN(n461) );
  XNOR2_X1 U406 ( .A(G140), .B(G137), .ZN(n526) );
  XNOR2_X1 U407 ( .A(n388), .B(n504), .ZN(n403) );
  XNOR2_X1 U408 ( .A(G134), .B(G131), .ZN(n504) );
  NAND2_X1 U409 ( .A1(n416), .A2(n445), .ZN(n447) );
  XNOR2_X1 U410 ( .A(n387), .B(n448), .ZN(n386) );
  INV_X1 U411 ( .A(KEYINPUT18), .ZN(n448) );
  XNOR2_X1 U412 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n387) );
  XNOR2_X1 U413 ( .A(n453), .B(n452), .ZN(n451) );
  INV_X1 U414 ( .A(KEYINPUT28), .ZN(n452) );
  NAND2_X1 U415 ( .A1(n381), .A2(n665), .ZN(n453) );
  XNOR2_X1 U416 ( .A(n440), .B(G478), .ZN(n554) );
  OR2_X1 U417 ( .A1(n638), .A2(G902), .ZN(n440) );
  NAND2_X1 U418 ( .A1(n513), .A2(n428), .ZN(n427) );
  XNOR2_X1 U419 ( .A(n422), .B(n420), .ZN(n511) );
  XNOR2_X1 U420 ( .A(n421), .B(G101), .ZN(n420) );
  XNOR2_X1 U421 ( .A(n423), .B(n473), .ZN(n422) );
  INV_X1 U422 ( .A(G119), .ZN(n421) );
  XNOR2_X1 U423 ( .A(G128), .B(G119), .ZN(n515) );
  XNOR2_X1 U424 ( .A(G110), .B(KEYINPUT93), .ZN(n516) );
  XNOR2_X1 U425 ( .A(n403), .B(n526), .ZN(n742) );
  XNOR2_X1 U426 ( .A(n397), .B(n561), .ZN(n690) );
  NOR2_X1 U427 ( .A1(n596), .A2(n597), .ZN(n616) );
  XNOR2_X1 U428 ( .A(n616), .B(KEYINPUT110), .ZN(n435) );
  XNOR2_X1 U429 ( .A(n503), .B(KEYINPUT22), .ZN(n537) );
  XNOR2_X1 U430 ( .A(n480), .B(n479), .ZN(n481) );
  INV_X1 U431 ( .A(KEYINPUT74), .ZN(n479) );
  NAND2_X1 U432 ( .A1(n665), .A2(n673), .ZN(n582) );
  NAND2_X1 U433 ( .A1(n725), .A2(n366), .ZN(n405) );
  NOR2_X1 U434 ( .A1(n407), .A2(n729), .ZN(n406) );
  NOR2_X1 U435 ( .A1(n364), .A2(G210), .ZN(n407) );
  XNOR2_X1 U436 ( .A(G146), .B(G137), .ZN(n505) );
  XOR2_X1 U437 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n506) );
  XNOR2_X1 U438 ( .A(KEYINPUT3), .B(G113), .ZN(n423) );
  XNOR2_X1 U439 ( .A(n372), .B(KEYINPUT48), .ZN(n633) );
  AND2_X1 U440 ( .A1(n376), .A2(n614), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n374), .B(n369), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n577), .B(n454), .ZN(n381) );
  INV_X1 U443 ( .A(KEYINPUT68), .ZN(n454) );
  OR2_X1 U444 ( .A1(G902), .A2(G237), .ZN(n483) );
  XNOR2_X1 U445 ( .A(G902), .B(KEYINPUT15), .ZN(n623) );
  INV_X1 U446 ( .A(KEYINPUT105), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n469), .B(KEYINPUT69), .ZN(n456) );
  XNOR2_X1 U448 ( .A(n436), .B(n491), .ZN(n493) );
  XNOR2_X1 U449 ( .A(G107), .B(G122), .ZN(n491) );
  XNOR2_X1 U450 ( .A(n437), .B(KEYINPUT9), .ZN(n436) );
  XNOR2_X1 U451 ( .A(KEYINPUT7), .B(KEYINPUT97), .ZN(n437) );
  XNOR2_X1 U452 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U453 ( .A(n460), .B(n457), .ZN(n464) );
  XNOR2_X1 U454 ( .A(n417), .B(n731), .ZN(n639) );
  XNOR2_X1 U455 ( .A(n589), .B(n365), .ZN(n615) );
  XNOR2_X1 U456 ( .A(n378), .B(n377), .ZN(n590) );
  INV_X1 U457 ( .A(KEYINPUT106), .ZN(n377) );
  NAND2_X1 U458 ( .A1(n451), .A2(n379), .ZN(n378) );
  XNOR2_X1 U459 ( .A(n606), .B(n380), .ZN(n379) );
  NOR2_X1 U460 ( .A1(n554), .A2(n562), .ZN(n595) );
  BUF_X1 U461 ( .A(n552), .Z(n606) );
  NAND2_X1 U462 ( .A1(n426), .A2(n429), .ZN(n425) );
  NAND2_X1 U463 ( .A1(G472), .A2(G902), .ZN(n429) );
  XNOR2_X1 U464 ( .A(n474), .B(n511), .ZN(n731) );
  XNOR2_X1 U465 ( .A(n530), .B(n472), .ZN(n474) );
  XNOR2_X1 U466 ( .A(KEYINPUT16), .B(G122), .ZN(n472) );
  XNOR2_X1 U467 ( .A(n383), .B(n384), .ZN(n727) );
  XNOR2_X1 U468 ( .A(n742), .B(n531), .ZN(n643) );
  XNOR2_X1 U469 ( .A(G146), .B(G101), .ZN(n528) );
  XNOR2_X1 U470 ( .A(n432), .B(n430), .ZN(n753) );
  XNOR2_X1 U471 ( .A(n431), .B(KEYINPUT107), .ZN(n430) );
  NAND2_X1 U472 ( .A1(n615), .A2(n595), .ZN(n432) );
  INV_X1 U473 ( .A(KEYINPUT40), .ZN(n431) );
  XNOR2_X1 U474 ( .A(n434), .B(KEYINPUT36), .ZN(n600) );
  NAND2_X1 U475 ( .A1(n435), .A2(n599), .ZN(n434) );
  XNOR2_X1 U476 ( .A(KEYINPUT71), .B(KEYINPUT35), .ZN(n565) );
  XNOR2_X1 U477 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n538) );
  NAND2_X1 U478 ( .A1(n537), .A2(n536), .ZN(n539) );
  NOR2_X1 U479 ( .A1(n603), .A2(n601), .ZN(n717) );
  XNOR2_X1 U480 ( .A(n595), .B(n438), .ZN(n714) );
  INV_X1 U481 ( .A(KEYINPUT101), .ZN(n438) );
  INV_X1 U482 ( .A(KEYINPUT60), .ZN(n410) );
  NOR2_X1 U483 ( .A1(n408), .A2(n404), .ZN(n642) );
  NOR2_X1 U484 ( .A1(n725), .A2(n364), .ZN(n408) );
  NAND2_X1 U485 ( .A1(n405), .A2(n406), .ZN(n404) );
  AND2_X1 U486 ( .A1(n547), .A2(KEYINPUT100), .ZN(n355) );
  XOR2_X1 U487 ( .A(n517), .B(n516), .Z(n356) );
  XOR2_X1 U488 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n357) );
  XOR2_X1 U489 ( .A(KEYINPUT91), .B(KEYINPUT14), .Z(n358) );
  NOR2_X1 U490 ( .A1(n470), .A2(n686), .ZN(n359) );
  OR2_X1 U491 ( .A1(n394), .A2(n653), .ZN(n360) );
  AND2_X1 U492 ( .A1(n651), .A2(n650), .ZN(n361) );
  AND2_X1 U493 ( .A1(n569), .A2(n568), .ZN(n362) );
  XOR2_X1 U494 ( .A(n490), .B(n489), .Z(n363) );
  XNOR2_X1 U495 ( .A(n641), .B(n640), .ZN(n364) );
  XNOR2_X1 U496 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n365) );
  AND2_X1 U497 ( .A1(n364), .A2(G210), .ZN(n366) );
  INV_X1 U498 ( .A(G902), .ZN(n428) );
  XOR2_X1 U499 ( .A(n700), .B(KEYINPUT62), .Z(n367) );
  XOR2_X1 U500 ( .A(n467), .B(n466), .Z(n368) );
  XNOR2_X1 U501 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n369) );
  NOR2_X1 U502 ( .A1(G952), .A2(n747), .ZN(n729) );
  INV_X1 U503 ( .A(n729), .ZN(n409) );
  XOR2_X1 U504 ( .A(KEYINPUT63), .B(n702), .Z(n370) );
  NAND2_X1 U505 ( .A1(n371), .A2(n560), .ZN(n397) );
  NAND2_X1 U506 ( .A1(n390), .A2(n389), .ZN(n371) );
  NOR2_X1 U507 ( .A1(n446), .A2(n362), .ZN(n445) );
  NAND2_X1 U508 ( .A1(n375), .A2(n373), .ZN(n372) );
  NAND2_X1 U509 ( .A1(n594), .A2(n449), .ZN(n376) );
  NAND2_X1 U510 ( .A1(n714), .A2(n381), .ZN(n596) );
  XNOR2_X2 U511 ( .A(n382), .B(n524), .ZN(n658) );
  NOR2_X1 U512 ( .A1(n727), .A2(G902), .ZN(n382) );
  XNOR2_X1 U513 ( .A(n356), .B(n741), .ZN(n383) );
  XNOR2_X1 U514 ( .A(n518), .B(n520), .ZN(n384) );
  XNOR2_X1 U515 ( .A(n478), .B(n385), .ZN(n393) );
  XNOR2_X1 U516 ( .A(n386), .B(n475), .ZN(n385) );
  XNOR2_X1 U517 ( .A(n393), .B(n388), .ZN(n417) );
  XNOR2_X2 U518 ( .A(n496), .B(KEYINPUT4), .ZN(n388) );
  NAND2_X1 U519 ( .A1(n548), .A2(n355), .ZN(n389) );
  NAND2_X1 U520 ( .A1(n391), .A2(n442), .ZN(n390) );
  NAND2_X1 U521 ( .A1(n548), .A2(n547), .ZN(n391) );
  NAND2_X1 U522 ( .A1(n564), .A2(n563), .ZN(n392) );
  XNOR2_X2 U523 ( .A(n441), .B(G143), .ZN(n496) );
  NOR2_X1 U524 ( .A1(n394), .A2(n663), .ZN(n550) );
  NOR2_X1 U525 ( .A1(n690), .A2(n394), .ZN(n396) );
  XNOR2_X2 U526 ( .A(n484), .B(KEYINPUT0), .ZN(n394) );
  NAND2_X1 U527 ( .A1(n395), .A2(n752), .ZN(n443) );
  NAND2_X1 U528 ( .A1(n534), .A2(n654), .ZN(n395) );
  XNOR2_X1 U529 ( .A(n395), .B(G110), .ZN(G12) );
  XNOR2_X1 U530 ( .A(n396), .B(KEYINPUT34), .ZN(n564) );
  NAND2_X1 U531 ( .A1(n567), .A2(KEYINPUT85), .ZN(n398) );
  NAND2_X1 U532 ( .A1(n399), .A2(n398), .ZN(n401) );
  INV_X1 U533 ( .A(n402), .ZN(n399) );
  NAND2_X1 U534 ( .A1(n401), .A2(n400), .ZN(n416) );
  NAND2_X1 U535 ( .A1(n402), .A2(KEYINPUT85), .ZN(n400) );
  XNOR2_X1 U536 ( .A(n512), .B(n403), .ZN(n700) );
  AND2_X4 U537 ( .A1(n635), .A2(n651), .ZN(n725) );
  NAND2_X1 U538 ( .A1(n548), .A2(n547), .ZN(n666) );
  XNOR2_X1 U539 ( .A(n411), .B(n410), .ZN(G60) );
  NAND2_X1 U540 ( .A1(n415), .A2(n409), .ZN(n411) );
  XNOR2_X1 U541 ( .A(n412), .B(n370), .ZN(G57) );
  NAND2_X1 U542 ( .A1(n414), .A2(n409), .ZN(n412) );
  XNOR2_X1 U543 ( .A(n413), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U544 ( .A1(n418), .A2(n409), .ZN(n413) );
  XNOR2_X1 U545 ( .A(n701), .B(n367), .ZN(n414) );
  XNOR2_X1 U546 ( .A(n636), .B(n368), .ZN(n415) );
  XNOR2_X2 U547 ( .A(n539), .B(n538), .ZN(n752) );
  NAND2_X1 U548 ( .A1(n628), .A2(n627), .ZN(n635) );
  XNOR2_X1 U549 ( .A(n637), .B(n419), .ZN(n418) );
  INV_X1 U550 ( .A(n638), .ZN(n419) );
  NAND2_X1 U551 ( .A1(n700), .A2(G472), .ZN(n426) );
  NOR2_X1 U552 ( .A1(n700), .A2(n427), .ZN(n424) );
  NOR2_X2 U553 ( .A1(n676), .A2(n675), .ZN(n578) );
  XNOR2_X2 U554 ( .A(n433), .B(KEYINPUT108), .ZN(n676) );
  NAND2_X1 U555 ( .A1(n672), .A2(n673), .ZN(n433) );
  XNOR2_X2 U556 ( .A(G128), .B(KEYINPUT64), .ZN(n441) );
  INV_X1 U557 ( .A(KEYINPUT100), .ZN(n442) );
  XNOR2_X2 U558 ( .A(n552), .B(n533), .ZN(n548) );
  NAND2_X1 U559 ( .A1(n443), .A2(KEYINPUT44), .ZN(n541) );
  NOR2_X1 U560 ( .A1(n443), .A2(KEYINPUT44), .ZN(n569) );
  NAND2_X1 U561 ( .A1(n444), .A2(n359), .ZN(n484) );
  NAND2_X1 U562 ( .A1(n590), .A2(n444), .ZN(n591) );
  XNOR2_X2 U563 ( .A(n598), .B(KEYINPUT19), .ZN(n444) );
  XNOR2_X1 U564 ( .A(n592), .B(n450), .ZN(n449) );
  AND2_X1 U565 ( .A1(n507), .A2(G214), .ZN(n457) );
  XNOR2_X1 U566 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n458) );
  INV_X1 U567 ( .A(KEYINPUT80), .ZN(n647) );
  INV_X1 U568 ( .A(n658), .ZN(n586) );
  XNOR2_X1 U569 ( .A(n511), .B(n510), .ZN(n512) );
  INV_X1 U570 ( .A(n598), .ZN(n599) );
  NOR2_X1 U571 ( .A1(n600), .A2(n654), .ZN(n720) );
  XNOR2_X1 U572 ( .A(KEYINPUT124), .B(KEYINPUT67), .ZN(n467) );
  XNOR2_X1 U573 ( .A(KEYINPUT10), .B(n475), .ZN(n741) );
  XNOR2_X1 U574 ( .A(n357), .B(n459), .ZN(n460) );
  XNOR2_X1 U575 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U576 ( .A(n741), .B(n465), .ZN(n488) );
  XNOR2_X1 U577 ( .A(n488), .B(KEYINPUT59), .ZN(n466) );
  XNOR2_X1 U578 ( .A(KEYINPUT92), .B(G898), .ZN(n734) );
  NOR2_X1 U579 ( .A1(n747), .A2(n734), .ZN(n730) );
  NAND2_X1 U580 ( .A1(n730), .A2(G902), .ZN(n468) );
  NAND2_X1 U581 ( .A1(G952), .A2(n747), .ZN(n573) );
  AND2_X1 U582 ( .A1(n468), .A2(n573), .ZN(n470) );
  NAND2_X1 U583 ( .A1(G237), .A2(G234), .ZN(n469) );
  XNOR2_X1 U584 ( .A(G110), .B(G107), .ZN(n471) );
  XNOR2_X1 U585 ( .A(n471), .B(G104), .ZN(n530) );
  INV_X1 U586 ( .A(G116), .ZN(n473) );
  XOR2_X1 U587 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n477) );
  NAND2_X1 U588 ( .A1(G224), .A2(n747), .ZN(n476) );
  XNOR2_X1 U589 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U590 ( .A1(n639), .A2(n623), .ZN(n482) );
  NAND2_X1 U591 ( .A1(G210), .A2(n483), .ZN(n480) );
  XNOR2_X2 U592 ( .A(n482), .B(n481), .ZN(n608) );
  NAND2_X1 U593 ( .A1(G214), .A2(n483), .ZN(n673) );
  NAND2_X2 U594 ( .A1(n608), .A2(n673), .ZN(n598) );
  NAND2_X1 U595 ( .A1(n623), .A2(G234), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n485), .B(KEYINPUT94), .ZN(n486) );
  XNOR2_X1 U597 ( .A(KEYINPUT20), .B(n486), .ZN(n521) );
  NAND2_X1 U598 ( .A1(n521), .A2(G221), .ZN(n487) );
  XNOR2_X1 U599 ( .A(n487), .B(KEYINPUT21), .ZN(n659) );
  XNOR2_X1 U600 ( .A(KEYINPUT13), .B(KEYINPUT96), .ZN(n490) );
  INV_X1 U601 ( .A(G475), .ZN(n489) );
  XNOR2_X1 U602 ( .A(G134), .B(G116), .ZN(n492) );
  XNOR2_X1 U603 ( .A(n493), .B(n492), .ZN(n500) );
  NAND2_X1 U604 ( .A1(n747), .A2(G234), .ZN(n495) );
  XNOR2_X1 U605 ( .A(n495), .B(n494), .ZN(n519) );
  NAND2_X1 U606 ( .A1(G217), .A2(n519), .ZN(n498) );
  INV_X1 U607 ( .A(n496), .ZN(n497) );
  XNOR2_X1 U608 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U609 ( .A(n500), .B(n499), .ZN(n638) );
  INV_X1 U610 ( .A(n554), .ZN(n601) );
  NOR2_X1 U611 ( .A1(n659), .A2(n675), .ZN(n501) );
  XOR2_X1 U612 ( .A(KEYINPUT98), .B(n501), .Z(n502) );
  INV_X1 U613 ( .A(n537), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n506), .B(n505), .ZN(n509) );
  NAND2_X1 U615 ( .A1(n507), .A2(G210), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U617 ( .A(G472), .ZN(n513) );
  INV_X1 U618 ( .A(n665), .ZN(n663) );
  INV_X1 U619 ( .A(n526), .ZN(n514) );
  XNOR2_X1 U620 ( .A(n515), .B(n514), .ZN(n518) );
  XOR2_X1 U621 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n517) );
  NAND2_X1 U622 ( .A1(G221), .A2(n519), .ZN(n520) );
  XOR2_X1 U623 ( .A(KEYINPUT25), .B(KEYINPUT70), .Z(n523) );
  NAND2_X1 U624 ( .A1(G217), .A2(n521), .ZN(n522) );
  XNOR2_X1 U625 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U626 ( .A1(n663), .A2(n658), .ZN(n525) );
  NAND2_X1 U627 ( .A1(n747), .A2(G227), .ZN(n527) );
  XNOR2_X1 U628 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U629 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U630 ( .A1(n643), .A2(n428), .ZN(n532) );
  XNOR2_X2 U631 ( .A(n532), .B(G469), .ZN(n552) );
  XNOR2_X1 U632 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n533) );
  INV_X1 U633 ( .A(n548), .ZN(n654) );
  XNOR2_X1 U634 ( .A(n665), .B(KEYINPUT6), .ZN(n597) );
  NAND2_X1 U635 ( .A1(n597), .A2(n658), .ZN(n535) );
  NOR2_X1 U636 ( .A1(n654), .A2(n535), .ZN(n536) );
  INV_X1 U637 ( .A(KEYINPUT65), .ZN(n540) );
  XNOR2_X1 U638 ( .A(n541), .B(n540), .ZN(n559) );
  NAND2_X1 U639 ( .A1(n597), .A2(n586), .ZN(n542) );
  OR2_X1 U640 ( .A1(n542), .A2(n548), .ZN(n543) );
  NOR2_X1 U641 ( .A1(n544), .A2(n543), .ZN(n546) );
  INV_X1 U642 ( .A(KEYINPUT99), .ZN(n545) );
  XNOR2_X1 U643 ( .A(n546), .B(n545), .ZN(n755) );
  OR2_X1 U644 ( .A1(n658), .A2(n659), .ZN(n653) );
  INV_X1 U645 ( .A(n653), .ZN(n547) );
  INV_X1 U646 ( .A(n666), .ZN(n549) );
  NAND2_X1 U647 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U648 ( .A(n551), .B(KEYINPUT31), .ZN(n718) );
  NOR2_X1 U649 ( .A1(n665), .A2(n360), .ZN(n553) );
  AND2_X1 U650 ( .A1(n553), .A2(n606), .ZN(n707) );
  OR2_X1 U651 ( .A1(n718), .A2(n707), .ZN(n556) );
  INV_X1 U652 ( .A(n562), .ZN(n603) );
  NOR2_X1 U653 ( .A1(n595), .A2(n717), .ZN(n677) );
  XOR2_X1 U654 ( .A(KEYINPUT77), .B(n677), .Z(n593) );
  INV_X1 U655 ( .A(n593), .ZN(n555) );
  AND2_X1 U656 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U657 ( .A1(n755), .A2(n557), .ZN(n558) );
  INV_X1 U658 ( .A(n597), .ZN(n560) );
  INV_X1 U659 ( .A(KEYINPUT33), .ZN(n561) );
  NOR2_X1 U660 ( .A1(n562), .A2(n601), .ZN(n563) );
  INV_X1 U661 ( .A(KEYINPUT44), .ZN(n566) );
  NAND2_X1 U662 ( .A1(G953), .A2(G902), .ZN(n570) );
  XOR2_X1 U663 ( .A(KEYINPUT103), .B(n572), .Z(n575) );
  NOR2_X1 U664 ( .A1(n686), .A2(n573), .ZN(n574) );
  NOR2_X1 U665 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n658), .A2(n585), .ZN(n577) );
  INV_X1 U667 ( .A(n590), .ZN(n579) );
  INV_X1 U668 ( .A(n608), .ZN(n619) );
  XNOR2_X1 U669 ( .A(n578), .B(KEYINPUT41), .ZN(n691) );
  XNOR2_X1 U670 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n580) );
  XOR2_X1 U671 ( .A(KEYINPUT104), .B(KEYINPUT30), .Z(n583) );
  XNOR2_X1 U672 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U673 ( .A1(n585), .A2(n584), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n586), .ZN(n587) );
  NOR2_X1 U675 ( .A1(n605), .A2(n587), .ZN(n588) );
  NAND2_X1 U676 ( .A1(n672), .A2(n588), .ZN(n589) );
  XNOR2_X2 U677 ( .A(n591), .B(KEYINPUT73), .ZN(n592) );
  NAND2_X1 U678 ( .A1(n592), .A2(n593), .ZN(n594) );
  NOR2_X1 U679 ( .A1(n658), .A2(n601), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n607) );
  AND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n712) );
  XNOR2_X1 U684 ( .A(n712), .B(KEYINPUT78), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n677), .A2(KEYINPUT47), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U687 ( .A(KEYINPUT76), .B(n612), .ZN(n613) );
  NOR2_X1 U688 ( .A1(n720), .A2(n613), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n717), .A2(n615), .ZN(n722) );
  AND2_X1 U690 ( .A1(n616), .A2(n673), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n617), .A2(n654), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(KEYINPUT43), .ZN(n620) );
  AND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n723) );
  INV_X1 U694 ( .A(n723), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n722), .A2(n621), .ZN(n622) );
  NOR2_X2 U696 ( .A1(n633), .A2(n622), .ZN(n746) );
  INV_X1 U697 ( .A(n623), .ZN(n626) );
  AND2_X1 U698 ( .A1(n746), .A2(n626), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n629), .A2(n624), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n625), .B(KEYINPUT82), .ZN(n628) );
  NAND2_X1 U701 ( .A1(KEYINPUT2), .A2(n626), .ZN(n627) );
  BUF_X2 U702 ( .A(n629), .Z(n732) );
  NAND2_X1 U703 ( .A1(KEYINPUT2), .A2(n722), .ZN(n630) );
  XOR2_X1 U704 ( .A(KEYINPUT75), .B(n630), .Z(n631) );
  OR2_X1 U705 ( .A1(n631), .A2(n723), .ZN(n632) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n732), .A2(n634), .ZN(n651) );
  NAND2_X1 U708 ( .A1(n725), .A2(G475), .ZN(n636) );
  NAND2_X1 U709 ( .A1(G478), .A2(n725), .ZN(n637) );
  XOR2_X1 U710 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n641) );
  XNOR2_X1 U711 ( .A(n639), .B(KEYINPUT86), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n642), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U713 ( .A(n568), .B(G122), .ZN(G24) );
  NAND2_X1 U714 ( .A1(n725), .A2(G469), .ZN(n645) );
  XNOR2_X1 U715 ( .A(n643), .B(n458), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X1 U717 ( .A1(n646), .A2(n729), .ZN(G54) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n746), .A2(KEYINPUT2), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n649), .B(KEYINPUT81), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n652), .A2(n361), .ZN(n695) );
  NAND2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n656) );
  XOR2_X1 U723 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U725 ( .A(KEYINPUT117), .B(n657), .ZN(n662) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U727 ( .A(KEYINPUT49), .B(n660), .Z(n661) );
  NAND2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n668) );
  NAND2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U731 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U732 ( .A(n669), .B(KEYINPUT51), .ZN(n670) );
  XNOR2_X1 U733 ( .A(KEYINPUT119), .B(n670), .ZN(n671) );
  NOR2_X1 U734 ( .A1(n691), .A2(n671), .ZN(n683) );
  NOR2_X1 U735 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U736 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U737 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U738 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U739 ( .A1(n680), .A2(n690), .ZN(n681) );
  XNOR2_X1 U740 ( .A(n681), .B(KEYINPUT120), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U742 ( .A(n684), .B(KEYINPUT121), .Z(n685) );
  XNOR2_X1 U743 ( .A(KEYINPUT52), .B(n685), .ZN(n689) );
  INV_X1 U744 ( .A(n686), .ZN(n687) );
  NAND2_X1 U745 ( .A1(n687), .A2(G952), .ZN(n688) );
  NOR2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n693) );
  NOR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U749 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U750 ( .A(n696), .B(KEYINPUT122), .ZN(n697) );
  OR2_X2 U751 ( .A1(n697), .A2(G953), .ZN(n699) );
  XNOR2_X1 U752 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(G75) );
  NAND2_X1 U754 ( .A1(G472), .A2(n725), .ZN(n701) );
  XOR2_X1 U755 ( .A(KEYINPUT87), .B(KEYINPUT111), .Z(n702) );
  NAND2_X1 U756 ( .A1(n714), .A2(n707), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(G104), .ZN(G6) );
  XOR2_X1 U758 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n705) );
  XNOR2_X1 U759 ( .A(G107), .B(KEYINPUT26), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  XOR2_X1 U761 ( .A(KEYINPUT27), .B(n706), .Z(n709) );
  NAND2_X1 U762 ( .A1(n707), .A2(n717), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n709), .B(n708), .ZN(G9) );
  XOR2_X1 U764 ( .A(G128), .B(KEYINPUT29), .Z(n711) );
  NAND2_X1 U765 ( .A1(n717), .A2(n592), .ZN(n710) );
  XNOR2_X1 U766 ( .A(n711), .B(n710), .ZN(G30) );
  XNOR2_X1 U767 ( .A(G143), .B(n712), .ZN(G45) );
  NAND2_X1 U768 ( .A1(n592), .A2(n714), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n713), .B(G146), .ZN(G48) );
  XOR2_X1 U770 ( .A(G113), .B(KEYINPUT115), .Z(n716) );
  NAND2_X1 U771 ( .A1(n718), .A2(n714), .ZN(n715) );
  XNOR2_X1 U772 ( .A(n716), .B(n715), .ZN(G15) );
  NAND2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n719), .B(G116), .ZN(G18) );
  XNOR2_X1 U775 ( .A(n720), .B(G125), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n721), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U777 ( .A(G134), .B(n722), .ZN(G36) );
  XOR2_X1 U778 ( .A(G140), .B(n723), .Z(n724) );
  XNOR2_X1 U779 ( .A(KEYINPUT116), .B(n724), .ZN(G42) );
  NAND2_X1 U780 ( .A1(G217), .A2(n725), .ZN(n726) );
  XNOR2_X1 U781 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U782 ( .A1(n729), .A2(n728), .ZN(G66) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n740) );
  NAND2_X1 U784 ( .A1(n732), .A2(n747), .ZN(n738) );
  NAND2_X1 U785 ( .A1(G953), .A2(G224), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n733), .B(KEYINPUT61), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U788 ( .A(n736), .B(KEYINPUT126), .ZN(n737) );
  NAND2_X1 U789 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(G69) );
  XNOR2_X1 U791 ( .A(n742), .B(n741), .ZN(n745) );
  XOR2_X1 U792 ( .A(G227), .B(n745), .Z(n743) );
  NAND2_X1 U793 ( .A1(G900), .A2(n743), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(G953), .ZN(n750) );
  XNOR2_X1 U795 ( .A(n746), .B(n745), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n750), .A2(n749), .ZN(G72) );
  XOR2_X1 U798 ( .A(G119), .B(KEYINPUT127), .Z(n751) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(G21) );
  XNOR2_X1 U800 ( .A(G131), .B(n753), .ZN(G33) );
  XNOR2_X1 U801 ( .A(n754), .B(G137), .ZN(G39) );
  XOR2_X1 U802 ( .A(G101), .B(n755), .Z(n756) );
  XNOR2_X1 U803 ( .A(KEYINPUT112), .B(n756), .ZN(G3) );
endmodule

