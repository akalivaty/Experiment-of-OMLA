//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n212), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n211), .B(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n229), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G107), .B(G116), .Z(new_n235));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n237), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT68), .ZN(new_n246));
  AND2_X1   g0046(.A1(KEYINPUT67), .A2(G45), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT67), .A2(G45), .ZN(new_n248));
  NOR3_X1   g0048(.A1(new_n247), .A2(new_n248), .A3(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n246), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  OR2_X1    g0053(.A1(KEYINPUT67), .A2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT67), .A2(G45), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(KEYINPUT68), .A3(new_n251), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G226), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n259), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT69), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(G1698), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n276), .B1(new_n277), .B2(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n262), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n266), .A2(new_n267), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n269), .A2(G190), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n208), .B1(new_n212), .B2(new_n270), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n209), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G58), .A2(G68), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n209), .B1(new_n293), .B2(new_n238), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n286), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT70), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n263), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n209), .A2(G1), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(G50), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n299), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n295), .B(new_n303), .C1(G50), .C2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n283), .A2(new_n284), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n268), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n285), .B(new_n306), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n269), .A2(new_n283), .A3(new_n284), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G200), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n285), .A4(new_n306), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n318), .A2(new_n320), .A3(new_n305), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n271), .A2(new_n273), .A3(G226), .A4(G1698), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n279), .A2(G1698), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(new_n271), .A3(new_n273), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G87), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT77), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT77), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(G33), .A3(G87), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n324), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT78), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n324), .A2(new_n326), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n262), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n262), .A2(G232), .A3(new_n264), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n259), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n309), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n278), .A2(new_n325), .B1(new_n328), .B2(new_n330), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n334), .B1(new_n341), .B2(new_n324), .ZN(new_n342));
  INV_X1    g0142(.A(new_n335), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n282), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI211_X1 g0144(.A(G190), .B(new_n337), .C1(new_n253), .C2(new_n258), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT80), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT80), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  INV_X1    g0148(.A(new_n258), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT68), .B1(new_n257), .B2(new_n251), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(new_n338), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n347), .B1(new_n336), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n340), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n304), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n287), .A2(new_n301), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n354), .A2(new_n287), .B1(new_n300), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n286), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT7), .B1(new_n274), .B2(new_n209), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  AOI211_X1 g0160(.A(new_n360), .B(G20), .C1(new_n271), .C2(new_n273), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G58), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n240), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n364), .B2(new_n293), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n290), .A2(G159), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n358), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT76), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n274), .A2(new_n371), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n360), .B1(new_n278), .B2(G20), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(G20), .B1(new_n271), .B2(new_n273), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n371), .B1(new_n375), .B2(KEYINPUT7), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n365), .A2(new_n366), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n369), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n357), .B1(new_n370), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n353), .A2(new_n381), .A3(KEYINPUT17), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT17), .B1(new_n353), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G169), .B1(new_n336), .B2(new_n339), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n337), .B1(new_n253), .B2(new_n258), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n344), .A2(G179), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n373), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n378), .B1(new_n390), .B2(G68), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n286), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n367), .A2(KEYINPUT16), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(KEYINPUT76), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(new_n372), .A3(new_n373), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n395), .B2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n356), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n388), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n388), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT79), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n388), .A2(new_n397), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT18), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT79), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n388), .A2(new_n397), .A3(new_n398), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n384), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n319), .A2(KEYINPUT75), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  INV_X1    g0209(.A(G232), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G1698), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(G226), .B2(G1698), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n409), .B1(new_n412), .B2(new_n274), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n253), .A2(new_n258), .B1(new_n413), .B2(new_n282), .ZN(new_n414));
  INV_X1    g0214(.A(G238), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT72), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n265), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n416), .B2(new_n265), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n414), .B2(new_n418), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n408), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT14), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(KEYINPUT73), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT73), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n414), .A2(new_n426), .A3(new_n418), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(KEYINPUT13), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n420), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(G179), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n408), .C1(new_n420), .C2(new_n422), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n424), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n304), .A2(G68), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT12), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n240), .A2(G20), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n437), .B1(new_n288), .B2(new_n277), .C1(new_n291), .C2(new_n238), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n286), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT11), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT11), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n441), .A3(new_n286), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n300), .A2(G68), .A3(new_n302), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n436), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT74), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n436), .A2(new_n443), .A3(KEYINPUT74), .A4(new_n444), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n433), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n428), .A2(G190), .A3(new_n429), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n448), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n420), .A2(new_n422), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n451), .B(new_n452), .C1(new_n309), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n287), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT15), .B(G87), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n458), .A2(new_n288), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n358), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n300), .A2(G77), .A3(new_n302), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n304), .A2(G77), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G244), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n265), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n253), .B2(new_n258), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n280), .A2(new_n415), .B1(new_n203), .B2(new_n278), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT71), .ZN(new_n469));
  INV_X1    g0269(.A(G1698), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n278), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(new_n410), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n275), .A2(KEYINPUT71), .A3(G232), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n467), .B1(new_n474), .B2(new_n262), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n464), .B1(G200), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n348), .B2(new_n475), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n475), .A2(G179), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n319), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(new_n464), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NOR4_X1   g0281(.A1(new_n323), .A2(new_n407), .A3(new_n455), .A4(new_n481), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n486), .A2(G264), .A3(new_n262), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n271), .A2(new_n273), .A3(G257), .A4(G1698), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n271), .A2(new_n273), .A3(G250), .A4(new_n470), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G294), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT93), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n262), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT93), .A4(new_n490), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n484), .A2(new_n250), .A3(G1), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n483), .A2(new_n496), .A3(new_n262), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n319), .ZN(new_n499));
  INV_X1    g0299(.A(new_n497), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n500), .B(new_n487), .C1(new_n493), .C2(new_n494), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n317), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  INV_X1    g0305(.A(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n288), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n209), .B2(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n278), .A2(new_n209), .A3(G87), .ZN(new_n512));
  XOR2_X1   g0312(.A(KEYINPUT89), .B(KEYINPUT22), .Z(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n512), .A2(KEYINPUT89), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n505), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n512), .A2(new_n513), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(KEYINPUT24), .A3(new_n516), .A4(new_n511), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n286), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n354), .A2(KEYINPUT90), .A3(KEYINPUT25), .A4(new_n203), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT90), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n298), .A2(new_n203), .A3(new_n299), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT25), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT91), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n524), .A2(new_n527), .A3(new_n525), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n524), .B2(new_n525), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n522), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT92), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n263), .A2(G33), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n300), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n531), .B1(new_n530), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n521), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n504), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  XNOR2_X1  g0340(.A(KEYINPUT81), .B(G97), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n209), .B(new_n540), .C1(new_n541), .C2(G33), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n506), .A2(G20), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n542), .A2(KEYINPUT20), .A3(new_n286), .A4(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT20), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n540), .A2(new_n209), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n202), .A2(KEYINPUT81), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT81), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n546), .B1(new_n550), .B2(new_n270), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n286), .A2(new_n543), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n545), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n300), .A2(G116), .A3(new_n532), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT88), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n300), .A2(KEYINPUT88), .A3(G116), .A4(new_n532), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n354), .A2(new_n506), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n554), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n278), .A2(G257), .A3(new_n470), .ZN(new_n561));
  XNOR2_X1  g0361(.A(KEYINPUT87), .B(G303), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n274), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G264), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n561), .B(new_n563), .C1(new_n280), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n282), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n282), .B1(new_n485), .B2(new_n483), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n500), .B1(G270), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n319), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n566), .A2(new_n568), .A3(G179), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n560), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n560), .A2(new_n569), .A3(KEYINPUT21), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n495), .A2(new_n348), .A3(new_n497), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n501), .B2(G200), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n578), .B(new_n521), .C1(new_n536), .C2(new_n537), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n566), .A2(new_n568), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n348), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n309), .B1(new_n566), .B2(new_n568), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n581), .A2(new_n560), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n539), .A2(new_n576), .A3(new_n579), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n304), .A2(new_n202), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n533), .B2(new_n202), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n291), .A2(new_n277), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n390), .B2(G107), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT82), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(G97), .A2(G107), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n204), .A2(KEYINPUT82), .A3(new_n591), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n550), .A2(KEYINPUT6), .A3(new_n203), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G20), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n589), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT83), .B1(new_n601), .B2(new_n286), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  AOI211_X1 g0403(.A(new_n603), .B(new_n358), .C1(new_n589), .C2(new_n600), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n587), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(new_n470), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT4), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n470), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n540), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n282), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n486), .A2(G257), .A3(new_n262), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n497), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n319), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n614), .B1(new_n282), .B2(new_n611), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n317), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n605), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n209), .B1(new_n597), .B2(new_n598), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n203), .B1(new_n373), .B2(new_n389), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(new_n624), .A3(new_n588), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n603), .B1(new_n625), .B2(new_n358), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n601), .A2(KEYINPUT83), .A3(new_n286), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n612), .A2(new_n615), .A3(new_n348), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(G200), .B2(new_n618), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n587), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G87), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n547), .A2(new_n549), .A3(new_n632), .A4(new_n203), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT19), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n209), .B1(new_n409), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n634), .B1(new_n541), .B2(new_n288), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n278), .A2(new_n209), .A3(G68), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n286), .B1(new_n354), .B2(new_n458), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n415), .A2(new_n470), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n465), .A2(G1698), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n271), .A2(new_n641), .A3(new_n273), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(G33), .A2(G116), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n282), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n484), .B2(G1), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n263), .A2(KEYINPUT84), .A3(G45), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G250), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n485), .A2(G274), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n262), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n646), .A2(new_n653), .A3(G190), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n533), .A2(G87), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n262), .B1(new_n643), .B2(new_n644), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n282), .B1(new_n650), .B2(new_n651), .ZN(new_n657));
  OAI21_X1  g0457(.A(G200), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n640), .A2(new_n654), .A3(new_n655), .A4(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(G169), .B1(new_n656), .B2(new_n657), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n646), .A2(new_n653), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n317), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT85), .ZN(new_n663));
  INV_X1    g0463(.A(new_n458), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n533), .A2(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n662), .A2(new_n663), .B1(new_n640), .B2(new_n665), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n660), .B(KEYINPUT85), .C1(new_n661), .C2(new_n317), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n659), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n622), .A2(new_n631), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT86), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT86), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n622), .A2(new_n671), .A3(new_n631), .A4(new_n668), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n585), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n482), .A2(new_n673), .ZN(G372));
  NOR2_X1   g0474(.A1(new_n399), .A2(new_n400), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT94), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n480), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT94), .A4(new_n464), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n679), .A2(new_n454), .B1(new_n449), .B2(new_n433), .ZN(new_n680));
  INV_X1    g0480(.A(new_n384), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n321), .B1(new_n682), .B2(new_n316), .ZN(new_n683));
  INV_X1    g0483(.A(new_n482), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n640), .A2(new_n655), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n654), .A2(new_n658), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n640), .A2(new_n665), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n662), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n605), .A2(new_n621), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n662), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n620), .B1(new_n628), .B2(new_n587), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n689), .B1(new_n693), .B2(new_n668), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n575), .A2(new_n574), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n518), .A2(new_n286), .A3(new_n520), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n530), .A2(new_n534), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT92), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(new_n699), .B2(new_n535), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n696), .B(new_n572), .C1(new_n700), .C2(new_n503), .ZN(new_n701));
  INV_X1    g0501(.A(new_n659), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n691), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n700), .B2(new_n578), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n701), .A2(new_n704), .A3(new_n622), .A4(new_n631), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n695), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n683), .B1(new_n684), .B2(new_n707), .ZN(G369));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n263), .A2(new_n209), .A3(G13), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n713));
  INV_X1    g0513(.A(G213), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G343), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT95), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n718), .A2(new_n560), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n710), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT96), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n710), .A2(new_n719), .A3(new_n583), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n709), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n504), .A2(new_n538), .A3(new_n717), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n579), .B1(new_n700), .B2(new_n717), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n539), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n539), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n576), .A2(new_n718), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n725), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(G399));
  INV_X1    g0532(.A(new_n213), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G41), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n633), .A2(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n206), .B2(new_n735), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n668), .A2(new_n605), .A3(new_n621), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n691), .B1(new_n740), .B2(KEYINPUT26), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n689), .B1(new_n693), .B2(new_n688), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n718), .B1(new_n743), .B2(new_n705), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n707), .A2(new_n718), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n670), .A2(new_n672), .ZN(new_n748));
  INV_X1    g0548(.A(new_n585), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(new_n717), .ZN(new_n750));
  INV_X1    g0550(.A(new_n661), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n573), .A2(new_n495), .A3(new_n618), .A4(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT30), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n580), .A2(new_n317), .A3(new_n661), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(KEYINPUT30), .A3(new_n618), .A4(new_n495), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n751), .A2(G179), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n498), .A2(new_n757), .A3(new_n616), .A4(new_n580), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n754), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n718), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n750), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G330), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n747), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n739), .B1(new_n769), .B2(G1), .ZN(G364));
  NAND2_X1  g0570(.A1(new_n721), .A2(new_n722), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n209), .A2(G13), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n263), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OR3_X1    g0575(.A1(new_n775), .A2(new_n734), .A3(KEYINPUT97), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT97), .B1(new_n775), .B2(new_n734), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n772), .A2(new_n723), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n208), .B1(G20), .B2(new_n319), .ZN(new_n782));
  NAND2_X1  g0582(.A1(G20), .A2(G179), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n348), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n209), .A2(G179), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n348), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G50), .A2(new_n786), .B1(new_n789), .B2(G107), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n348), .A2(G179), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n209), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G97), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n785), .A2(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n790), .B(new_n794), .C1(new_n240), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G190), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n799), .A2(KEYINPUT32), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G87), .ZN(new_n804));
  OAI21_X1  g0604(.A(KEYINPUT32), .B1(new_n799), .B2(new_n800), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n784), .A2(new_n798), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n783), .A2(new_n348), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n278), .B1(new_n807), .B2(new_n277), .C1(new_n809), .C2(new_n363), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n797), .A2(new_n801), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G317), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT33), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n812), .A2(KEYINPUT33), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n795), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n786), .A2(G326), .ZN(new_n816));
  INV_X1    g0616(.A(G303), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n802), .ZN(new_n818));
  INV_X1    g0618(.A(new_n799), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G329), .B1(G322), .B2(new_n808), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n274), .C1(new_n821), .C2(new_n807), .ZN(new_n822));
  INV_X1    g0622(.A(G294), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n792), .A2(new_n823), .B1(new_n788), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n818), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n782), .B1(new_n811), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n733), .A2(new_n274), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(G355), .B1(new_n506), .B2(new_n733), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n244), .A2(new_n484), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n733), .A2(new_n278), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n254), .A2(new_n256), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n206), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n829), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(G13), .A2(G33), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(G20), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n782), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n778), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n837), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n827), .B(new_n839), .C1(new_n771), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n781), .A2(new_n841), .ZN(G396));
  NAND3_X1  g0642(.A1(new_n477), .A2(new_n480), .A3(new_n717), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n579), .A2(new_n622), .A3(new_n631), .A4(new_n688), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n710), .B1(new_n538), .B2(new_n504), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n740), .A2(KEYINPUT26), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n691), .A3(new_n690), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n844), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT99), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT99), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n706), .A2(new_n852), .A3(new_n844), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n677), .A2(new_n464), .A3(new_n678), .A4(new_n718), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n477), .B(new_n480), .C1(new_n463), .C2(new_n717), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n854), .B1(new_n746), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n779), .B1(new_n858), .B2(new_n767), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n767), .B2(new_n858), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n782), .A2(new_n835), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n779), .B1(G77), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n786), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n824), .A2(new_n796), .B1(new_n863), .B2(new_n817), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G107), .B2(new_n803), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n809), .A2(new_n823), .B1(new_n799), .B2(new_n821), .ZN(new_n866));
  INV_X1    g0666(.A(new_n807), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n278), .B(new_n866), .C1(G116), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n788), .A2(new_n632), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n865), .A2(new_n794), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n867), .A2(G159), .B1(G143), .B2(new_n808), .ZN(new_n872));
  INV_X1    g0672(.A(G137), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n872), .B1(new_n863), .B2(new_n873), .C1(new_n289), .C2(new_n796), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT34), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n789), .A2(G68), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n274), .B1(new_n819), .B2(G132), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n793), .A2(G58), .B1(new_n803), .B2(G50), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n874), .A2(new_n875), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n871), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n862), .B1(new_n882), .B2(new_n782), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n857), .B2(new_n836), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n860), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(G384));
  OR2_X1    g0686(.A1(new_n599), .A2(KEYINPUT35), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n599), .A2(KEYINPUT35), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(G116), .A3(new_n210), .A4(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT36), .Z(new_n890));
  OAI211_X1 g0690(.A(new_n207), .B(G77), .C1(new_n363), .C2(new_n240), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n263), .B(G13), .C1(new_n891), .C2(new_n239), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n675), .A2(new_n715), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n452), .A2(new_n717), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n450), .A2(new_n454), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n450), .B2(new_n454), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n480), .A2(new_n718), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT100), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n854), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n380), .A2(new_n286), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT16), .B1(new_n377), .B2(new_n367), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n356), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n715), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n407), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n353), .A2(new_n381), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n388), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n397), .B1(new_n388), .B2(new_n715), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT37), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n911), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n910), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n407), .A2(new_n908), .B1(new_n918), .B2(new_n915), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(KEYINPUT38), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n894), .B1(new_n903), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n916), .A2(new_n911), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT101), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n917), .B1(new_n916), .B2(new_n911), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n397), .A2(new_n715), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n384), .B2(new_n675), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n910), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n920), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT102), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n915), .A2(new_n918), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n909), .B2(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n715), .A2(new_n906), .B1(new_n353), .B2(new_n381), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n917), .B1(new_n938), .B2(new_n913), .ZN(new_n939));
  INV_X1    g0739(.A(new_n918), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT38), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n407), .B2(new_n908), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT39), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT102), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n920), .A2(new_n932), .A3(new_n944), .A4(new_n933), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n935), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n450), .A2(new_n718), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n923), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n683), .B1(new_n747), .B2(new_n684), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n855), .A2(new_n856), .ZN(new_n952));
  INV_X1    g0752(.A(new_n898), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n450), .A2(new_n454), .A3(new_n896), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n922), .A2(new_n766), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n764), .B1(new_n673), .B2(new_n717), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n857), .B1(new_n897), .B2(new_n898), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n958), .A2(new_n959), .A3(new_n957), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n920), .A2(new_n932), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n956), .A2(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n684), .B2(new_n958), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(new_n482), .A3(new_n766), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(G330), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n951), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n263), .B2(new_n773), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n951), .A2(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n893), .B1(new_n968), .B2(new_n969), .ZN(G367));
  AOI22_X1  g0770(.A1(new_n819), .A2(G137), .B1(G150), .B2(new_n808), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n971), .B(new_n278), .C1(new_n238), .C2(new_n807), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n796), .A2(new_n800), .B1(new_n802), .B2(new_n363), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n789), .A2(G77), .ZN(new_n974));
  INV_X1    g0774(.A(G143), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n863), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n792), .A2(new_n240), .ZN(new_n977));
  NOR4_X1   g0777(.A1(new_n972), .A2(new_n973), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT110), .Z(new_n979));
  NAND3_X1  g0779(.A1(new_n803), .A2(KEYINPUT46), .A3(G116), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT108), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n793), .A2(G107), .B1(new_n795), .B2(G294), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G311), .A2(new_n786), .B1(new_n789), .B2(new_n550), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT46), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n802), .B2(new_n506), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT109), .B(G317), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n799), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n274), .B1(new_n807), .B2(new_n824), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n562), .C2(new_n808), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n982), .A2(new_n983), .A3(new_n985), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n979), .B1(new_n981), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT47), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n782), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n688), .B1(new_n685), .B2(new_n717), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n691), .A2(new_n717), .A3(new_n685), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n837), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n233), .A2(new_n831), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(new_n838), .C1(new_n213), .C2(new_n458), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT107), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n1000), .A2(new_n1001), .A3(new_n778), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n993), .A2(new_n996), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n631), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n717), .B1(new_n628), .B2(new_n587), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1004), .A2(new_n693), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n622), .A2(new_n717), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n731), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT45), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n731), .A2(new_n1008), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT44), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n1011), .A2(new_n728), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n728), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n727), .B(new_n730), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n723), .A2(KEYINPUT104), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n723), .A2(KEYINPUT104), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1022), .A2(new_n768), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n769), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT105), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n734), .B(KEYINPUT41), .Z(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n768), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT105), .B1(new_n1030), .B2(new_n1027), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n774), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1008), .A2(new_n727), .A3(new_n730), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT42), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1006), .A2(new_n538), .A3(new_n504), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n718), .B1(new_n1036), .B2(new_n622), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1034), .B2(KEYINPUT42), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n994), .A2(new_n995), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1035), .A2(new_n1038), .B1(KEYINPUT43), .B2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(KEYINPUT43), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n728), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n1008), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1042), .B1(KEYINPUT103), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1044), .A2(KEYINPUT103), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT106), .B1(new_n1033), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n775), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1049), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT106), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1003), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT111), .ZN(G387));
  INV_X1    g0856(.A(new_n1023), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1022), .A2(new_n768), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n734), .B(KEYINPUT115), .Z(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1020), .A2(new_n1021), .A3(new_n775), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n274), .B1(new_n819), .B2(G150), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n277), .B2(new_n802), .C1(new_n202), .C2(new_n788), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT112), .Z(new_n1064));
  NOR2_X1   g0864(.A1(new_n792), .A2(new_n458), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n238), .B2(new_n809), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT113), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n795), .A2(new_n456), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n786), .A2(G159), .B1(new_n867), .B2(G68), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1064), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT114), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n278), .B1(new_n819), .B2(G326), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n792), .A2(new_n824), .B1(new_n802), .B2(new_n823), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n986), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n867), .A2(new_n562), .B1(new_n1075), .B2(new_n808), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n786), .A2(G322), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n821), .C2(new_n796), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n1079), .B2(new_n1078), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT49), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1073), .B1(new_n506), .B2(new_n788), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n782), .B1(new_n1072), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n831), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n229), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n832), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n736), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n828), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n736), .B(new_n484), .C1(new_n240), .C2(new_n277), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT50), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n287), .B2(G50), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n456), .A2(KEYINPUT50), .A3(new_n238), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1090), .A2(new_n1095), .B1(G107), .B2(new_n213), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n778), .B1(new_n1096), .B2(new_n838), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1085), .B(new_n1097), .C1(new_n727), .C2(new_n840), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1061), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1060), .A2(new_n1099), .ZN(G393));
  OAI21_X1  g0900(.A(new_n1057), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n1024), .A3(new_n1059), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1008), .A2(new_n840), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n838), .B1(new_n213), .B2(new_n541), .C1(new_n237), .C2(new_n1086), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n779), .A2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n786), .A2(G150), .B1(G159), .B2(new_n808), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT51), .Z(new_n1107));
  OAI221_X1 g0907(.A(new_n278), .B1(new_n799), .B2(new_n975), .C1(new_n287), .C2(new_n807), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n796), .A2(new_n238), .B1(new_n802), .B2(new_n240), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n792), .A2(new_n277), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1110), .A2(new_n869), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1107), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n786), .A2(G317), .B1(G311), .B2(new_n808), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT52), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n793), .A2(G116), .B1(new_n803), .B2(G283), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n562), .A2(new_n795), .B1(new_n789), .B2(G107), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n867), .A2(G294), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n278), .B1(new_n819), .B2(G322), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1113), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1105), .B1(new_n1121), .B2(new_n782), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1016), .A2(new_n775), .B1(new_n1103), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1102), .A2(new_n1123), .ZN(G390));
  AOI21_X1  g0924(.A(new_n901), .B1(new_n744), .B2(new_n857), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n961), .B1(new_n450), .B2(new_n718), .C1(new_n1125), .C2(new_n899), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n852), .B1(new_n706), .B2(new_n844), .ZN(new_n1127));
  AOI211_X1 g0927(.A(KEYINPUT99), .B(new_n843), .C1(new_n695), .C2(new_n705), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n902), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n899), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n947), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1126), .B1(new_n1131), .B2(new_n946), .ZN(new_n1132));
  NOR4_X1   g0932(.A1(new_n958), .A2(new_n899), .A3(new_n709), .A4(new_n952), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n709), .B1(new_n750), .B2(new_n765), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(new_n1130), .A3(new_n857), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1136), .B(new_n1126), .C1(new_n1131), .C2(new_n946), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1134), .A2(new_n775), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n779), .B1(new_n456), .B2(new_n861), .ZN(new_n1140));
  INV_X1    g0940(.A(G132), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n809), .A2(new_n1141), .B1(new_n807), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n274), .B(new_n1143), .C1(G125), .C2(new_n819), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n802), .A2(new_n289), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G137), .A2(new_n795), .B1(new_n789), .B2(G50), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n792), .A2(new_n800), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G128), .B2(new_n786), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1111), .B1(G283), .B2(new_n786), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n203), .B2(new_n796), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n807), .A2(new_n541), .B1(new_n799), .B2(new_n823), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n278), .B(new_n1153), .C1(G116), .C2(new_n808), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n804), .A3(new_n877), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1150), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1140), .B1(new_n1156), .B2(new_n782), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n946), .B2(new_n836), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1138), .A2(new_n1139), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1139), .B1(new_n1138), .B2(new_n1158), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT116), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1135), .A2(new_n482), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n683), .B(new_n1164), .C1(new_n747), .C2(new_n684), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n899), .B1(new_n767), .B2(new_n952), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1136), .A3(new_n1125), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1130), .B1(new_n1135), .B2(new_n857), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1129), .B1(new_n1168), .B2(new_n1133), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1165), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1163), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1134), .A2(new_n1170), .A3(new_n1137), .ZN(new_n1173));
  AND4_X1   g0973(.A1(new_n1162), .A2(new_n1172), .A3(new_n1059), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1059), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1162), .B1(new_n1176), .B2(new_n1173), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1161), .B1(new_n1174), .B2(new_n1177), .ZN(G378));
  NAND2_X1  g0978(.A1(new_n305), .A2(new_n715), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n316), .A2(new_n322), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n316), .B2(new_n322), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  OR3_X1    g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n962), .B2(G330), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n955), .A2(new_n766), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n909), .A2(new_n936), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1189), .A2(new_n910), .B1(new_n909), .B2(new_n919), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n957), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n960), .A2(new_n961), .ZN(new_n1192));
  AND4_X1   g0992(.A1(G330), .A2(new_n1191), .A3(new_n1192), .A4(new_n1186), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n949), .B1(new_n1187), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(G330), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1186), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1191), .A2(new_n1192), .A3(new_n1186), .A4(G330), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1197), .A2(new_n948), .A3(new_n923), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1194), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n775), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n779), .B1(G50), .B2(new_n861), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT119), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n278), .A2(G41), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n824), .B2(new_n799), .C1(new_n458), .C2(new_n807), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n977), .B(new_n1205), .C1(G77), .C2(new_n803), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n789), .A2(G58), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n796), .B2(new_n202), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G116), .B2(new_n786), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n808), .A2(G107), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT118), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1206), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT58), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1204), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n238), .C1(G33), .C2(G41), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n786), .A2(G125), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n796), .B2(new_n1141), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n867), .A2(G137), .B1(G128), .B2(new_n808), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n802), .B2(new_n1142), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G150), .C2(new_n793), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n789), .A2(G159), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n819), .C2(G124), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1217), .B1(new_n1213), .B2(new_n1212), .C1(new_n1224), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1203), .B1(new_n1229), .B2(new_n782), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1186), .B2(new_n836), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1201), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1165), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1173), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1200), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1175), .B1(new_n1238), .B2(new_n1234), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1232), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G375));
  NAND2_X1  g1041(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n775), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n779), .B1(G68), .B2(new_n861), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n795), .A2(G116), .B1(new_n867), .B2(G107), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT121), .Z(new_n1246));
  OAI21_X1  g1046(.A(new_n274), .B1(new_n799), .B2(new_n817), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G283), .B2(new_n808), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G294), .A2(new_n786), .B1(new_n803), .B2(G97), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n974), .A4(new_n1066), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n786), .A2(G132), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n800), .B2(new_n802), .C1(new_n796), .C2(new_n1142), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n793), .A2(G50), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n867), .A2(G150), .B1(G137), .B2(new_n808), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n274), .B1(new_n819), .B2(G128), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1207), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1246), .A2(new_n1250), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1244), .B1(new_n1257), .B2(new_n782), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1130), .B2(new_n836), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1243), .A2(new_n1259), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(KEYINPUT122), .Z(new_n1261));
  NOR2_X1   g1061(.A1(new_n1242), .A2(new_n1233), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT120), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1171), .A2(new_n1028), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(G381));
  XOR2_X1   g1065(.A(new_n1240), .B(KEYINPUT123), .Z(new_n1266));
  NAND4_X1  g1066(.A1(new_n1099), .A2(new_n1060), .A3(new_n841), .A4(new_n781), .ZN(new_n1267));
  OR3_X1    g1067(.A1(G390), .A2(G384), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1176), .A2(new_n1173), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1138), .A2(new_n1158), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1268), .A2(G381), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1266), .A2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(G387), .A2(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT124), .ZN(G407));
  NOR2_X1   g1075(.A1(new_n714), .A2(G343), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1271), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n714), .B1(new_n1266), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G407), .A2(new_n1279), .ZN(G409));
  INV_X1    g1080(.A(new_n1271), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1201), .B(new_n1231), .C1(new_n1235), .C2(new_n1027), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1240), .A2(G378), .A3(KEYINPUT125), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT125), .B1(new_n1240), .B2(G378), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1175), .B1(new_n1262), .B2(KEYINPUT60), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1171), .A2(KEYINPUT60), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1263), .B2(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1289), .A2(new_n1261), .A3(G384), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1289), .B2(new_n1261), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1286), .A2(new_n1277), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G2897), .B(new_n1276), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1289), .A2(new_n1261), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n885), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1289), .A2(new_n1261), .A3(G384), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1276), .A2(G2897), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1240), .A2(G378), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT125), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1240), .A2(G378), .A3(KEYINPUT125), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1305), .A2(new_n1306), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1302), .B1(new_n1307), .B2(new_n1276), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1286), .A2(new_n1309), .A3(new_n1277), .A4(new_n1292), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1294), .A2(new_n1295), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(G393), .A2(G396), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1267), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G390), .B1(new_n1313), .B2(KEYINPUT111), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(G390), .B2(new_n1313), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1055), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1033), .A2(KEYINPUT106), .A3(new_n1049), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1053), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1313), .A2(KEYINPUT111), .ZN(new_n1320));
  MUX2_X1   g1120(.A(new_n1320), .B(new_n1313), .S(G390), .Z(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1321), .A3(new_n1003), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1316), .A2(KEYINPUT126), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT126), .B1(new_n1316), .B2(new_n1322), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1311), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1286), .A2(new_n1277), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT61), .B1(new_n1327), .B2(new_n1302), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1293), .A2(new_n1329), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1316), .A2(new_n1322), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1286), .A2(KEYINPUT63), .A3(new_n1277), .A4(new_n1292), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1328), .A2(new_n1330), .A3(new_n1331), .A4(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1326), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT127), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1326), .A2(KEYINPUT127), .A3(new_n1333), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(G405));
  OAI22_X1  g1138(.A1(new_n1284), .A2(new_n1285), .B1(new_n1240), .B2(new_n1271), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1339), .B(new_n1292), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1325), .B(new_n1340), .ZN(G402));
endmodule


