//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT79), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212));
  OAI22_X1  g011(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(KEYINPUT22), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(KEYINPUT22), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n208), .B(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT24), .ZN(new_n220));
  XOR2_X1   g019(.A(G183gat), .B(G190gat), .Z(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(KEYINPUT24), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  INV_X1    g022(.A(G169gat), .ZN(new_n224));
  INV_X1    g023(.A(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(new_n227), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT66), .Z(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n230), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n236), .B(KEYINPUT68), .C1(new_n233), .C2(new_n227), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n229), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n227), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n235), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT64), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n242), .A2(new_n246), .A3(new_n235), .A4(new_n243), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n247), .A3(new_n222), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(new_n223), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n248), .B2(new_n223), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n241), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n254));
  AOI21_X1  g053(.A(G190gat), .B1(new_n254), .B2(KEYINPUT69), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT27), .B(G183gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(KEYINPUT69), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(KEYINPUT28), .A3(new_n219), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n226), .A2(KEYINPUT26), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n235), .B(new_n262), .C1(new_n233), .C2(KEYINPUT26), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n218), .B2(new_n219), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n253), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(KEYINPUT78), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT78), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n240), .A2(new_n251), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n265), .B1(new_n272), .B2(new_n250), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n250), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n276), .A2(new_n240), .A3(new_n251), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT77), .B1(new_n277), .B2(new_n265), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT77), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n253), .A2(new_n279), .A3(new_n266), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT29), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n268), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n217), .B1(new_n275), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n268), .B1(new_n278), .B2(new_n280), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n273), .A2(KEYINPUT29), .A3(new_n269), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n217), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n205), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n205), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n274), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(new_n268), .B2(new_n282), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n287), .B(new_n290), .C1(new_n292), .C2(new_n217), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(new_n293), .A3(KEYINPUT30), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n284), .A2(new_n288), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n290), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299));
  XOR2_X1   g098(.A(G127gat), .B(G134gat), .Z(new_n300));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT70), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT1), .B1(new_n303), .B2(KEYINPUT70), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OR3_X1    g106(.A1(new_n303), .A2(KEYINPUT71), .A3(KEYINPUT1), .ZN(new_n308));
  INV_X1    g107(.A(new_n300), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G141gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G148gat), .ZN(new_n313));
  INV_X1    g112(.A(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G141gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n313), .A2(new_n315), .B1(KEYINPUT2), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(KEYINPUT80), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(G155gat), .A3(G162gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT81), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT81), .B1(new_n317), .B2(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n319), .A2(new_n316), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n317), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n311), .B1(new_n331), .B2(KEYINPUT3), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n326), .A2(new_n327), .B1(new_n317), .B2(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n299), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n305), .A2(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n333), .B2(new_n334), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n328), .A2(new_n334), .A3(new_n330), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT82), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n331), .A2(new_n337), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(KEYINPUT4), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(new_n331), .B2(new_n337), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n333), .B(new_n337), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(new_n342), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT85), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n331), .A2(new_n337), .A3(new_n346), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT4), .B1(new_n333), .B2(new_n311), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n346), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n333), .A2(new_n311), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(KEYINPUT85), .B(new_n365), .C1(new_n344), .C2(KEYINPUT4), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n363), .B(new_n366), .C1(new_n336), .C2(new_n340), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n342), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OR3_X1    g168(.A1(new_n354), .A2(new_n359), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n359), .B1(new_n354), .B2(new_n369), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(KEYINPUT6), .B(new_n359), .C1(new_n354), .C2(new_n369), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n298), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G22gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT31), .B(G50gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n216), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n381));
  INV_X1    g180(.A(G228gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT86), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n216), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n208), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT86), .A3(new_n215), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n281), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n386), .A2(KEYINPUT87), .A3(new_n281), .A4(new_n388), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n334), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n384), .B1(new_n393), .B2(new_n331), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n334), .B1(new_n216), .B2(KEYINPUT29), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n331), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n382), .B(new_n383), .C1(new_n396), .C2(new_n381), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n380), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n394), .A2(new_n397), .A3(new_n380), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n379), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n378), .A3(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G15gat), .B(G43gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n267), .A2(new_n311), .ZN(new_n408));
  AND2_X1   g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n273), .A2(new_n337), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n411), .B2(KEYINPUT32), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n407), .A2(KEYINPUT72), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(KEYINPUT72), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(KEYINPUT33), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(KEYINPUT32), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT74), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n409), .B1(new_n408), .B2(new_n410), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(KEYINPUT73), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(KEYINPUT73), .A3(new_n421), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT34), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n422), .B2(KEYINPUT73), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n424), .B2(new_n425), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n420), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n420), .ZN(new_n432));
  INV_X1    g231(.A(new_n427), .ZN(new_n433));
  INV_X1    g232(.A(new_n425), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n423), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n435), .A3(new_n428), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n404), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n376), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT35), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT35), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n376), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n376), .A2(new_n404), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n375), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n290), .B1(new_n295), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT38), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n216), .B1(new_n285), .B2(new_n286), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT37), .B(new_n449), .C1(new_n292), .C2(new_n216), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n445), .A2(new_n451), .A3(new_n293), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT37), .B1(new_n284), .B2(new_n288), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n448), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n367), .A2(new_n343), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT88), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT88), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n367), .A2(new_n460), .A3(new_n343), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT39), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n457), .B1(new_n462), .B2(new_n359), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n367), .A2(new_n460), .A3(new_n343), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n460), .B1(new_n367), .B2(new_n343), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(KEYINPUT89), .A3(new_n358), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n464), .B1(new_n352), .B2(new_n342), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n459), .A2(new_n461), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT40), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  INV_X1    g272(.A(new_n471), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n473), .B(new_n474), .C1(new_n463), .C2(new_n468), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n294), .A2(new_n372), .A3(new_n297), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT90), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n462), .A2(new_n457), .A3(new_n359), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT89), .B1(new_n467), .B2(new_n358), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n471), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n473), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n469), .A2(KEYINPUT40), .A3(new_n471), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n482), .A2(new_n477), .A3(KEYINPUT90), .A4(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n456), .B1(new_n478), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n404), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n444), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n489));
  INV_X1    g288(.A(new_n431), .ZN(new_n490));
  INV_X1    g289(.A(new_n436), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n431), .A2(KEYINPUT36), .A3(new_n436), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n442), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G43gat), .B(G50gat), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n496), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  NOR3_X1   g296(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n498), .B(KEYINPUT91), .Z(new_n499));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OAI221_X1 g300(.A(new_n497), .B1(KEYINPUT15), .B2(new_n496), .C1(new_n499), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G29gat), .ZN(new_n503));
  INV_X1    g302(.A(G36gat), .ZN(new_n504));
  OAI22_X1  g303(.A1(new_n501), .A2(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(KEYINPUT15), .A3(new_n496), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G1gat), .B2(new_n510), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(G8gat), .Z(new_n514));
  NAND3_X1  g313(.A1(new_n502), .A2(KEYINPUT17), .A3(new_n506), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n507), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT18), .A3(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n507), .B(new_n514), .Z(new_n522));
  XOR2_X1   g321(.A(new_n520), .B(KEYINPUT13), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n520), .A3(new_n518), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n521), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G197gat), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT11), .B(G169gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT12), .Z(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n521), .A2(new_n535), .A3(new_n524), .A4(new_n527), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n495), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  INV_X1    g341(.A(G92gat), .ZN(new_n543));
  AOI22_X1  g342(.A1(KEYINPUT8), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G99gat), .B(G106gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n509), .A2(new_n515), .A3(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n507), .A2(new_n547), .B1(KEYINPUT41), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(new_n549), .B2(new_n551), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT99), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n550), .A2(KEYINPUT41), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT97), .ZN(new_n558));
  XOR2_X1   g357(.A(G134gat), .B(G162gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT98), .Z(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n553), .B2(new_n554), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n556), .B1(new_n555), .B2(new_n561), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n568));
  INV_X1    g367(.A(G57gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(G64gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT92), .B(G57gat), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(G64gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n568), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(KEYINPUT92), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G57gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n580), .A3(G64gat), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n569), .A2(G64gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n574), .A2(new_n575), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(KEYINPUT93), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n577), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n573), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n575), .ZN(new_n588));
  XOR2_X1   g387(.A(G57gat), .B(G64gat), .Z(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(KEYINPUT9), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT94), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n593));
  AOI211_X1 g392(.A(new_n593), .B(new_n590), .C1(new_n577), .C2(new_n585), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n548), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI221_X4 g394(.A(new_n568), .B1(new_n574), .B2(new_n575), .C1(new_n581), .C2(new_n582), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT93), .B1(new_n583), .B2(new_n584), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n598), .A2(new_n547), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT10), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n593), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n586), .A2(KEYINPUT94), .A3(new_n591), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n547), .A2(KEYINPUT10), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n567), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n605), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n599), .B1(new_n604), .B2(new_n548), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT100), .B(new_n609), .C1(new_n610), .C2(KEYINPUT10), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n609), .B1(new_n610), .B2(KEYINPUT10), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n608), .B(KEYINPUT101), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n617), .B1(new_n623), .B2(new_n614), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n517), .B1(new_n604), .B2(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n604), .B2(KEYINPUT21), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n592), .A2(new_n594), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT21), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n627), .ZN(new_n632));
  INV_X1    g431(.A(G127gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n633), .B1(new_n629), .B2(new_n632), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n636), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n604), .A2(KEYINPUT21), .A3(new_n628), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n641));
  OAI21_X1  g440(.A(G127gat), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n642), .B2(new_n634), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n644));
  INV_X1    g443(.A(G155gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n638), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n636), .B1(new_n635), .B2(new_n637), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n642), .A2(new_n639), .A3(new_n634), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n626), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n647), .B1(new_n638), .B2(new_n643), .ZN(new_n654));
  INV_X1    g453(.A(new_n626), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n646), .A3(new_n650), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n652), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n653), .B1(new_n652), .B2(new_n657), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n566), .B(new_n625), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n538), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n445), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  INV_X1    g463(.A(new_n298), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n538), .A2(new_n665), .A3(new_n661), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n662), .A2(new_n669), .A3(new_n665), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NOR4_X1   g471(.A1(new_n666), .A2(new_n669), .A3(KEYINPUT42), .A4(new_n667), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT103), .B1(new_n666), .B2(G8gat), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n666), .A2(KEYINPUT103), .A3(G8gat), .ZN(new_n675));
  OAI22_X1  g474(.A1(new_n672), .A2(new_n673), .B1(new_n674), .B2(new_n675), .ZN(G1325gat));
  INV_X1    g475(.A(G15gat), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n490), .A2(new_n491), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n494), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n492), .A2(KEYINPUT104), .A3(new_n493), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n538), .A2(new_n661), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n680), .B1(new_n677), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n680), .B(KEYINPUT105), .C1(new_n677), .C2(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1326gat));
  AND2_X1   g489(.A1(new_n538), .A2(new_n404), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n661), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n652), .A2(new_n657), .ZN(new_n695));
  INV_X1    g494(.A(new_n653), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n652), .A2(new_n653), .A3(new_n657), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n625), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n699), .A2(new_n566), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n538), .A2(new_n503), .A3(new_n445), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n376), .A2(new_n437), .A3(new_n440), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n440), .B1(new_n376), .B2(new_n437), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT106), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n439), .A2(new_n708), .A3(new_n441), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n482), .A2(new_n477), .A3(new_n483), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT90), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n455), .B1(new_n713), .B2(new_n484), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n443), .B1(new_n714), .B2(new_n404), .ZN(new_n715));
  INV_X1    g514(.A(new_n684), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n710), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n704), .B1(new_n717), .B2(new_n566), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n566), .A2(new_n704), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n495), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n537), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n699), .A2(new_n722), .A3(new_n700), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n724), .A2(new_n445), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n703), .B1(new_n725), .B2(new_n503), .ZN(G1328gat));
  AND2_X1   g525(.A1(new_n538), .A2(new_n701), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n504), .A3(new_n665), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(KEYINPUT46), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n724), .A2(new_n665), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n729), .B(new_n730), .C1(new_n731), .C2(new_n504), .ZN(G1329gat));
  INV_X1    g531(.A(G43gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n727), .A2(new_n733), .A3(new_n679), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n718), .A2(new_n720), .A3(new_n684), .A4(new_n723), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G43gat), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n734), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1330gat));
  NOR2_X1   g539(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n741));
  NOR4_X1   g540(.A1(new_n699), .A2(G50gat), .A3(new_n566), .A4(new_n700), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n691), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n720), .A3(new_n404), .A4(new_n723), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n744), .B1(new_n743), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n699), .A2(new_n566), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n717), .A2(new_n537), .A3(new_n750), .A4(new_n625), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n445), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(new_n571), .Z(G1332gat));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n665), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT49), .B(G64gat), .Z(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n754), .B2(new_n756), .ZN(G1333gat));
  NAND2_X1  g556(.A1(new_n751), .A2(new_n684), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n678), .A2(G71gat), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n758), .A2(G71gat), .B1(new_n751), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n751), .A2(new_n404), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  INV_X1    g562(.A(new_n566), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n699), .A2(new_n537), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n486), .A2(new_n487), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n684), .B1(new_n766), .B2(new_n443), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n764), .B(new_n765), .C1(new_n767), .C2(new_n710), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n700), .ZN(new_n770));
  INV_X1    g569(.A(new_n717), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n771), .A2(new_n772), .A3(new_n764), .A4(new_n765), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OR4_X1    g573(.A1(G85gat), .A2(new_n770), .A3(new_n375), .A4(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n699), .A2(new_n537), .A3(new_n625), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n721), .A2(new_n445), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT108), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G85gat), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(KEYINPUT108), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  NAND4_X1  g580(.A1(new_n769), .A2(new_n773), .A3(new_n665), .A4(new_n700), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n543), .ZN(new_n783));
  NAND2_X1  g582(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n298), .A2(new_n543), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n718), .A2(new_n720), .A3(new_n776), .A4(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n783), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n784), .B1(new_n783), .B2(new_n788), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(G1337gat));
  OR4_X1    g590(.A1(G99gat), .A2(new_n770), .A3(new_n678), .A4(new_n774), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n721), .A2(new_n684), .A3(new_n776), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G99gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1338gat));
  NAND4_X1  g594(.A1(new_n718), .A2(new_n720), .A3(new_n404), .A4(new_n776), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT53), .B1(new_n797), .B2(KEYINPUT110), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n487), .A2(G106gat), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n769), .A2(new_n773), .A3(new_n700), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n800), .B(new_n797), .C1(KEYINPUT110), .C2(KEYINPUT53), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(G1339gat));
  INV_X1    g603(.A(new_n699), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n621), .B(new_n609), .C1(new_n610), .C2(KEYINPUT10), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT54), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n613), .B1(new_n620), .B2(new_n567), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n611), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n622), .C1(new_n601), .C2(new_n606), .ZN(new_n812));
  INV_X1    g611(.A(new_n617), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n806), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n612), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n819));
  INV_X1    g618(.A(new_n817), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(KEYINPUT111), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT112), .B1(new_n822), .B2(new_n618), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n824), .B(new_n619), .C1(new_n818), .C2(new_n821), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n537), .B(new_n815), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n519), .A2(new_n520), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n522), .A2(new_n523), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n532), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n536), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n700), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n764), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n566), .A2(new_n830), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n815), .B(new_n834), .C1(new_n823), .C2(new_n825), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n805), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n660), .A2(new_n537), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n375), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n437), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n665), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n722), .A2(G113gat), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT113), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n404), .B1(new_n837), .B2(new_n839), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n665), .A2(new_n375), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n679), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n722), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n845), .A2(new_n849), .ZN(G1340gat));
  INV_X1    g649(.A(G120gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n848), .A2(new_n851), .A3(new_n625), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n842), .A2(new_n700), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(G1341gat));
  NOR3_X1   g653(.A1(new_n848), .A2(new_n633), .A3(new_n805), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT114), .Z(new_n856));
  NAND2_X1  g655(.A1(new_n842), .A2(new_n699), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(G127gat), .B1(new_n858), .B2(KEYINPUT115), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n858), .A2(KEYINPUT115), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(G1342gat));
  NAND2_X1  g660(.A1(new_n298), .A2(new_n764), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT116), .Z(new_n863));
  OR3_X1    g662(.A1(new_n841), .A2(G134gat), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n848), .B2(new_n566), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n684), .A2(new_n487), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(new_n840), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n537), .A2(new_n312), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT119), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n870), .A2(new_n298), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n684), .A2(new_n375), .A3(new_n665), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n837), .A2(new_n839), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n404), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n404), .A2(KEYINPUT57), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n822), .A2(new_n618), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n537), .A2(new_n815), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n832), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n566), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n699), .B1(new_n882), .B2(new_n835), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n883), .B2(new_n838), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT117), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n886), .B(new_n878), .C1(new_n883), .C2(new_n838), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n875), .B1(new_n877), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G141gat), .B1(new_n889), .B2(new_n722), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(KEYINPUT118), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n895), .B(new_n875), .C1(new_n877), .C2(new_n888), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n537), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G141gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n874), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n893), .B1(new_n899), .B2(KEYINPUT58), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n873), .B1(new_n897), .B2(G141gat), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(KEYINPUT120), .A3(new_n891), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n892), .B1(new_n900), .B2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n870), .A2(new_n298), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n904), .B(G148gat), .C1(new_n905), .C2(new_n700), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n876), .A2(new_n878), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n883), .A2(new_n838), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT57), .B1(new_n908), .B2(new_n404), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n700), .A3(new_n875), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n314), .B1(new_n911), .B2(KEYINPUT59), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n894), .A2(new_n904), .A3(new_n700), .A4(new_n896), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(G1345gat));
  NAND3_X1  g713(.A1(new_n905), .A2(new_n645), .A3(new_n699), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n894), .A2(new_n699), .A3(new_n896), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n645), .ZN(G1346gat));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n764), .A3(new_n896), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G162gat), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n863), .A2(G162gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n870), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT121), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(G1347gat));
  AOI21_X1  g722(.A(new_n445), .B1(new_n837), .B2(new_n839), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n924), .A2(new_n665), .A3(new_n437), .ZN(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n537), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n665), .A2(new_n375), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n678), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n846), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n722), .A2(new_n224), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(G1348gat));
  INV_X1    g730(.A(new_n929), .ZN(new_n932));
  OAI21_X1  g731(.A(G176gat), .B1(new_n932), .B2(new_n625), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n925), .A2(new_n225), .A3(new_n700), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1349gat));
  AOI21_X1  g734(.A(new_n218), .B1(new_n929), .B2(new_n699), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n699), .A2(new_n256), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n925), .B2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT60), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n938), .B(new_n940), .ZN(G1350gat));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n219), .B1(new_n929), .B2(new_n764), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n219), .A3(new_n764), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n944), .A2(new_n945), .A3(new_n942), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n950), .ZN(G1351gat));
  AND3_X1   g750(.A1(new_n869), .A2(new_n665), .A3(new_n924), .ZN(new_n952));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952), .B2(new_n537), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n684), .A2(new_n927), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n910), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n537), .A2(G197gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  INV_X1    g756(.A(G204gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n952), .A2(new_n958), .A3(new_n700), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT62), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n955), .B2(new_n700), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n960), .A2(new_n961), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n910), .A2(new_n699), .A3(new_n954), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G211gat), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n964), .A2(KEYINPUT126), .A3(new_n965), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n964), .B2(new_n965), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n963), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n952), .A2(new_n210), .A3(new_n699), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1354gat));
  AOI21_X1  g774(.A(G218gat), .B1(new_n952), .B2(new_n764), .ZN(new_n976));
  XOR2_X1   g775(.A(new_n976), .B(KEYINPUT127), .Z(new_n977));
  NOR2_X1   g776(.A1(new_n566), .A2(new_n211), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n955), .B2(new_n978), .ZN(G1355gat));
endmodule


