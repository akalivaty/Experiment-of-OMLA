//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202));
  NOR4_X1   g001(.A1(KEYINPUT91), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT91), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT92), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT88), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n208), .A2(new_n209), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n208), .B2(new_n214), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n218));
  OAI21_X1  g017(.A(G36gat), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT90), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(G43gat), .A2(G50gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G43gat), .A2(G50gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT15), .ZN(new_n225));
  OAI211_X1 g024(.A(KEYINPUT90), .B(G36gat), .C1(new_n217), .C2(new_n218), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n227), .A3(new_n223), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n221), .A2(new_n225), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n215), .A2(new_n216), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n221), .A2(new_n226), .ZN(new_n231));
  NOR3_X1   g030(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(new_n212), .B2(new_n213), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(new_n225), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n202), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G15gat), .B(G22gat), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(KEYINPUT93), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT93), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT16), .B1(new_n241), .B2(G1gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n238), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n237), .B1(new_n243), .B2(KEYINPUT94), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(G1gat), .B2(new_n238), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n245), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n208), .A2(new_n214), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT92), .ZN(new_n251));
  INV_X1    g050(.A(new_n231), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n208), .A2(new_n209), .A3(new_n214), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n225), .A2(new_n228), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT15), .B(new_n224), .C1(new_n231), .C2(new_n233), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(KEYINPUT17), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n236), .A2(new_n249), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G229gat), .A2(G233gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT95), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n255), .A2(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n248), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n258), .A2(KEYINPUT18), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT18), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n260), .B(KEYINPUT13), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n255), .A2(new_n246), .A3(new_n247), .A4(new_n256), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G113gat), .B(G141gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G169gat), .B(G197gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT12), .ZN(new_n276));
  AND4_X1   g075(.A1(new_n263), .A2(new_n266), .A3(new_n270), .A4(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n269), .B1(new_n264), .B2(new_n265), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n278), .B2(new_n263), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT32), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT23), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n284), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n285), .B2(new_n282), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT24), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n287), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n294), .A2(KEYINPUT64), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(KEYINPUT64), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n292), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n287), .A2(new_n300), .A3(KEYINPUT25), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n287), .A2(new_n300), .A3(KEYINPUT65), .A4(KEYINPUT25), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G113gat), .B(G120gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(KEYINPUT1), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT68), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n306), .B2(KEYINPUT1), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G134gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OR4_X1    g111(.A1(new_n309), .A2(new_n306), .A3(new_n311), .A4(KEYINPUT1), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT67), .B1(new_n318), .B2(KEYINPUT26), .ZN(new_n321));
  OAI221_X1 g120(.A(new_n315), .B1(KEYINPUT26), .B2(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G183gat), .ZN(new_n323));
  OR3_X1    g122(.A1(new_n323), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT27), .B1(new_n323), .B2(KEYINPUT66), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n288), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT27), .B(G183gat), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n331), .B2(KEYINPUT28), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n322), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n305), .A2(new_n314), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT69), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n305), .A2(new_n333), .ZN(new_n336));
  INV_X1    g135(.A(new_n314), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n305), .A2(new_n339), .A3(new_n314), .A4(new_n333), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n281), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n343), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT33), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n345), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(KEYINPUT33), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n344), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n344), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n338), .A2(new_n340), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n359), .A2(new_n342), .A3(new_n335), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n360), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n341), .B2(new_n343), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n364), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n353), .B(new_n366), .C1(new_n356), .C2(new_n357), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT73), .B(KEYINPUT22), .Z(new_n369));
  NAND2_X1  g168(.A1(G211gat), .A2(G218gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G211gat), .ZN(new_n372));
  INV_X1    g171(.A(G218gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n370), .ZN(new_n375));
  XOR2_X1   g174(.A(G197gat), .B(G204gat), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n370), .B(new_n374), .C1(new_n369), .C2(new_n376), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n305), .A2(new_n333), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n305), .B2(new_n333), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n381), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n305), .A2(new_n333), .A3(new_n382), .ZN(new_n387));
  INV_X1    g186(.A(new_n333), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n296), .A2(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n304), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n387), .B(new_n380), .C1(new_n390), .C2(new_n384), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT74), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n383), .A2(new_n385), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT74), .A3(new_n380), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT75), .ZN(new_n397));
  XOR2_X1   g196(.A(G8gat), .B(G36gat), .Z(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT76), .ZN(new_n399));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT75), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n393), .A2(new_n403), .A3(new_n395), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n397), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(G141gat), .B(G148gat), .Z(new_n406));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n407));
  OAI211_X1 g206(.A(G155gat), .B(G162gat), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409));
  NAND2_X1  g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(G155gat), .B2(G162gat), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n406), .A2(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G141gat), .B(G148gat), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n413), .A2(KEYINPUT78), .ZN(new_n414));
  INV_X1    g213(.A(G155gat), .ZN(new_n415));
  INV_X1    g214(.A(G162gat), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n413), .A2(KEYINPUT78), .B1(new_n417), .B2(new_n410), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n408), .A2(new_n412), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n314), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT79), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n314), .A2(new_n423), .A3(new_n419), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n412), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n414), .A2(new_n418), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n314), .B1(KEYINPUT3), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n419), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n314), .A2(KEYINPUT4), .A3(new_n419), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n425), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n421), .B(new_n424), .C1(new_n419), .C2(new_n314), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n427), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT5), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n314), .A2(new_n423), .A3(new_n419), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n423), .B1(new_n314), .B2(new_n419), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT4), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT5), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n420), .A2(new_n422), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n442), .A2(new_n434), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT0), .ZN(new_n448));
  XNOR2_X1  g247(.A(G57gat), .B(G85gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n446), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n438), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT4), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n430), .A2(KEYINPUT3), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n337), .A2(new_n455), .A3(new_n433), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n426), .A3(new_n435), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT5), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n450), .B(new_n445), .C1(new_n453), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n450), .B1(new_n439), .B2(new_n445), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n452), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT30), .B1(new_n396), .B2(new_n401), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465));
  AOI211_X1 g264(.A(new_n465), .B(new_n402), .C1(new_n393), .C2(new_n395), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G78gat), .B(G106gat), .ZN(new_n468));
  INV_X1    g267(.A(G50gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n433), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n433), .A2(KEYINPUT83), .A3(new_n474), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n381), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(G228gat), .A2(G233gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n432), .B1(new_n381), .B2(KEYINPUT29), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n430), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n378), .A2(KEYINPUT82), .A3(new_n379), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n474), .B1(new_n378), .B2(KEYINPUT82), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n432), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n486), .A2(new_n430), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n380), .B1(new_n433), .B2(new_n474), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n480), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G22gat), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n483), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n483), .B2(new_n489), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n473), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n483), .A2(new_n489), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G22gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n483), .A2(new_n489), .A3(new_n490), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n496), .A3(new_n472), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT35), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  AND4_X1   g297(.A1(new_n405), .A2(new_n463), .A3(new_n467), .A4(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n368), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n365), .A2(new_n367), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n463), .A2(new_n498), .A3(new_n467), .A4(new_n405), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT86), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n464), .ZN(new_n506));
  INV_X1    g305(.A(new_n466), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n405), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT80), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n460), .B(new_n459), .C1(new_n462), .C2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n462), .A2(new_n509), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n452), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n361), .A2(new_n363), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n361), .B2(new_n363), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n358), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n493), .A2(new_n497), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n367), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT35), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n519), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n442), .A2(new_n456), .A3(new_n444), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n427), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n524), .A2(new_n427), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT39), .B1(new_n437), .B2(new_n427), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n526), .B(new_n450), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n462), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n427), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(KEYINPUT39), .C1(new_n427), .C2(new_n437), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(KEYINPUT40), .A3(new_n450), .A4(new_n526), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n467), .A2(new_n405), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n523), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n397), .A2(KEYINPUT37), .A3(new_n404), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT37), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n396), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(KEYINPUT38), .A3(new_n402), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n386), .B2(new_n391), .ZN(new_n542));
  AOI211_X1 g341(.A(new_n401), .B(new_n542), .C1(new_n396), .C2(new_n539), .ZN(new_n543));
  OAI22_X1  g342(.A1(new_n538), .A2(new_n541), .B1(new_n543), .B2(KEYINPUT38), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n396), .A2(new_n401), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n452), .B(new_n545), .C1(new_n461), .C2(new_n462), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT84), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n519), .B(new_n549), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n537), .A2(new_n548), .B1(new_n513), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n518), .A2(new_n367), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT36), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n365), .A2(new_n554), .A3(new_n367), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n280), .B1(new_n522), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT96), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G57gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G64gat), .ZN(new_n563));
  INV_X1    g362(.A(G64gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(G57gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n563), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n567), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n567), .ZN(new_n572));
  NOR2_X1   g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT97), .B1(new_n569), .B2(new_n567), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n568), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n571), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(KEYINPUT98), .B(new_n568), .C1(new_n575), .C2(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G127gat), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n249), .B1(new_n582), .B2(new_n581), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G127gat), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n589), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n590), .A2(new_n591), .A3(new_n587), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(new_n415), .ZN(new_n595));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n586), .A2(new_n587), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(new_n592), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT7), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(G85gat), .A3(G92gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G99gat), .B(G106gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n608), .B1(new_n607), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n236), .A2(new_n257), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n261), .A2(new_n615), .B1(KEYINPUT41), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT99), .Z(new_n622));
  AND2_X1   g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n622), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n628), .B1(new_n623), .B2(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n602), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n579), .A2(new_n580), .A3(new_n615), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n615), .B1(new_n579), .B2(new_n580), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n635), .A2(new_n636), .A3(KEYINPUT10), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n580), .A4(new_n615), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n634), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n634), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(new_n635), .B2(new_n636), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G120gat), .B(G148gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT100), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT101), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n640), .A2(new_n642), .A3(new_n648), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT102), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n643), .A2(new_n653), .A3(new_n649), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n633), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n561), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n512), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n239), .ZN(G1324gat));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  INV_X1    g460(.A(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n536), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n662), .A2(KEYINPUT42), .A3(new_n536), .A4(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(G8gat), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(G1325gat));
  OR3_X1    g468(.A1(new_n658), .A2(G15gat), .A3(new_n502), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n365), .A2(new_n554), .A3(new_n367), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n554), .B1(new_n518), .B2(new_n367), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT103), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n553), .A2(new_n674), .A3(new_n555), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n658), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n677), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n550), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NOR3_X1   g480(.A1(new_n602), .A2(new_n632), .A3(new_n656), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n559), .B2(new_n560), .ZN(new_n684));
  INV_X1    g483(.A(new_n512), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n217), .A2(new_n218), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT45), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(KEYINPUT45), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n500), .B1(new_n368), .B2(new_n499), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT86), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n690), .B(new_n521), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n551), .A2(new_n675), .A3(new_n673), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n690), .B1(new_n505), .B2(new_n521), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n631), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n631), .A2(KEYINPUT44), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n522), .B2(new_n556), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n655), .B(KEYINPUT104), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n280), .A3(new_n602), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n699), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n512), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n688), .B(new_n689), .C1(new_n686), .C2(new_n707), .ZN(G1328gat));
  INV_X1    g507(.A(new_n684), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n536), .A2(new_n206), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n709), .A2(KEYINPUT46), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n706), .B2(new_n508), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT46), .B1(new_n709), .B2(new_n710), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(G1329gat));
  OAI21_X1  g513(.A(G43gat), .B1(new_n706), .B2(new_n676), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n502), .A2(G43gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n709), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n706), .B2(new_n519), .ZN(new_n720));
  INV_X1    g519(.A(new_n550), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(G50gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n684), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(KEYINPUT48), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n699), .A2(new_n550), .A3(new_n702), .A4(new_n705), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n725), .A2(KEYINPUT106), .A3(G50gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n723), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT106), .B1(new_n725), .B2(G50gat), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n724), .B1(new_n729), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n522), .A2(KEYINPUT105), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n694), .A3(new_n693), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n266), .A2(new_n263), .A3(new_n270), .ZN(new_n733));
  INV_X1    g532(.A(new_n276), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n278), .A2(new_n263), .A3(new_n276), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n633), .A2(new_n703), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n732), .A2(KEYINPUT107), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n512), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(new_n562), .ZN(G1332gat));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n508), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  AND2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n746), .B2(new_n747), .ZN(G1333gat));
  AND2_X1   g549(.A1(new_n741), .A2(new_n742), .ZN(new_n751));
  INV_X1    g550(.A(G71gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n752), .A3(new_n368), .ZN(new_n753));
  OAI21_X1  g552(.A(G71gat), .B1(new_n743), .B2(new_n676), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n753), .B2(new_n754), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(G1334gat));
  NAND2_X1  g557(.A1(new_n751), .A2(new_n550), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n602), .A2(new_n737), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n656), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n699), .A2(new_n702), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n699), .A2(new_n766), .A3(new_n702), .A4(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n512), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n631), .B(new_n761), .C1(new_n695), .C2(new_n696), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT51), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n732), .A2(new_n772), .A3(new_n631), .A4(new_n761), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n774), .A2(new_n610), .A3(new_n685), .A4(new_n656), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n769), .A2(new_n775), .ZN(G1336gat));
  NOR3_X1   g575(.A1(new_n703), .A2(new_n508), .A3(G92gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G92gat), .B1(new_n764), .B2(new_n508), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n768), .B2(new_n508), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n770), .B(new_n783), .Z(new_n784));
  XOR2_X1   g583(.A(new_n777), .B(KEYINPUT110), .Z(new_n785));
  AOI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n780), .B1(new_n781), .B2(new_n786), .ZN(G1337gat));
  XNOR2_X1  g586(.A(KEYINPUT112), .B(G99gat), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n774), .A2(new_n368), .A3(new_n656), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n768), .A2(new_n676), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(new_n788), .ZN(G1338gat));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AOI211_X1 g592(.A(new_n701), .B(new_n762), .C1(new_n697), .C2(new_n698), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n523), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n703), .A2(G106gat), .A3(new_n519), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n771), .A2(new_n773), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n792), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G106gat), .B1(new_n764), .B2(new_n519), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n801), .A2(KEYINPUT113), .A3(new_n798), .A4(new_n797), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n765), .A2(new_n550), .A3(new_n767), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n804), .A2(G106gat), .B1(new_n784), .B2(new_n796), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n805), .B2(new_n798), .ZN(G1339gat));
  AOI21_X1  g605(.A(new_n260), .B1(new_n258), .B2(new_n262), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n262), .A2(new_n268), .A3(new_n267), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n275), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n652), .A2(new_n736), .A3(new_n654), .A4(new_n809), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n640), .A2(new_n642), .A3(new_n648), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n634), .C1(new_n637), .C2(new_n639), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n638), .A2(new_n641), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n637), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n581), .A2(new_n616), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT10), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n579), .A2(new_n580), .A3(new_n615), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n641), .B1(new_n820), .B2(new_n638), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n814), .B(new_n649), .C1(new_n816), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n811), .B1(new_n812), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n815), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n813), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n812), .B1(new_n640), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n648), .B1(new_n821), .B2(new_n813), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n826), .A2(KEYINPUT114), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT114), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n810), .B1(new_n830), .B2(new_n280), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT115), .B(new_n810), .C1(new_n830), .C2(new_n280), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n632), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n830), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n836), .A2(new_n736), .A3(new_n631), .A4(new_n809), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n602), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AND4_X1   g637(.A1(new_n280), .A2(new_n602), .A3(new_n632), .A4(new_n655), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT116), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n834), .A2(new_n632), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n827), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n826), .A2(KEYINPUT114), .A3(new_n827), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n737), .A3(new_n823), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT115), .B1(new_n847), .B2(new_n810), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n837), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n602), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852));
  INV_X1    g651(.A(new_n839), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n840), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n721), .A2(new_n368), .ZN(new_n856));
  NOR4_X1   g655(.A1(new_n855), .A2(new_n512), .A3(new_n536), .A4(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n280), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT117), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT116), .B(new_n839), .C1(new_n849), .C2(new_n850), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n520), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n863), .A2(KEYINPUT118), .A3(new_n685), .A4(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n840), .A2(new_n854), .A3(new_n685), .A4(new_n864), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n536), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n280), .A2(G113gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n860), .B1(new_n870), .B2(new_n871), .ZN(G1340gat));
  AOI21_X1  g671(.A(G120gat), .B1(new_n869), .B2(new_n656), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n857), .A2(G120gat), .A3(new_n704), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1341gat));
  NAND3_X1  g676(.A1(new_n869), .A2(new_n589), .A3(new_n602), .ZN(new_n878));
  OAI21_X1  g677(.A(G127gat), .B1(new_n858), .B2(new_n850), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  INV_X1    g679(.A(KEYINPUT56), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n536), .A2(new_n632), .A3(G134gat), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n865), .B2(new_n868), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n857), .A2(new_n631), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n881), .A2(new_n884), .B1(new_n885), .B2(G134gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n866), .A2(new_n867), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n866), .A2(new_n867), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n882), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n887), .B1(new_n890), .B2(KEYINPUT56), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n884), .A2(KEYINPUT120), .A3(new_n881), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n895), .B(new_n886), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1343gat));
  NOR2_X1   g696(.A1(new_n855), .A2(new_n519), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n676), .A2(new_n685), .A3(new_n508), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n831), .A2(new_n632), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n602), .B1(new_n902), .B2(new_n837), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n550), .B1(new_n903), .B2(new_n839), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(KEYINPUT57), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G141gat), .B1(new_n906), .B2(new_n280), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n676), .A2(new_n523), .ZN(new_n908));
  AND4_X1   g707(.A1(new_n685), .A2(new_n863), .A3(new_n508), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n280), .A2(G141gat), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n909), .A2(new_n910), .B1(KEYINPUT122), .B2(KEYINPUT58), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g711(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n912), .B(new_n913), .ZN(G1344gat));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(G148gat), .C1(new_n906), .C2(new_n655), .ZN(new_n916));
  INV_X1    g715(.A(G148gat), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n898), .A2(KEYINPUT57), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n904), .A2(new_n899), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n901), .A2(new_n655), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n916), .B1(new_n922), .B2(new_n915), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n909), .A2(new_n917), .A3(new_n656), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1345gat));
  AOI21_X1  g724(.A(G155gat), .B1(new_n909), .B2(new_n602), .ZN(new_n926));
  INV_X1    g725(.A(new_n906), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n602), .A2(G155gat), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT123), .Z(new_n929));
  AOI21_X1  g728(.A(new_n926), .B1(new_n927), .B2(new_n929), .ZN(G1346gat));
  AOI21_X1  g729(.A(G162gat), .B1(new_n909), .B2(new_n631), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n632), .A2(new_n416), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n927), .B2(new_n932), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n685), .A2(new_n508), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT124), .Z(new_n935));
  NAND4_X1  g734(.A1(new_n863), .A2(new_n721), .A3(new_n368), .A4(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(new_n316), .A3(new_n280), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n855), .A2(new_n685), .A3(new_n508), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n864), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n737), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n941), .B2(new_n316), .ZN(G1348gat));
  OAI21_X1  g741(.A(G176gat), .B1(new_n936), .B2(new_n703), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n656), .A2(new_n317), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n939), .B2(new_n944), .ZN(G1349gat));
  OAI21_X1  g744(.A(G183gat), .B1(new_n936), .B2(new_n850), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n602), .A2(new_n329), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n936), .B2(new_n632), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n951));
  OR2_X1    g750(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n953));
  NAND2_X1  g752(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n330), .A3(new_n631), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n951), .A2(new_n953), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n955), .B(new_n956), .C1(new_n957), .C2(new_n952), .ZN(G1351gat));
  NAND3_X1  g757(.A1(new_n920), .A2(new_n676), .A3(new_n935), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(new_n280), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n938), .A2(new_n737), .A3(new_n908), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n938), .A2(new_n908), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(G204gat), .A3(new_n655), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  OAI21_X1  g765(.A(G204gat), .B1(new_n959), .B2(new_n703), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1353gat));
  OAI21_X1  g767(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n959), .B2(new_n850), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n972));
  NAND2_X1  g771(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n970), .B(new_n973), .C1(new_n959), .C2(new_n850), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n938), .A2(new_n372), .A3(new_n602), .A4(new_n908), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n959), .B2(new_n632), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n631), .A2(new_n373), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n964), .B2(new_n978), .ZN(G1355gat));
endmodule


