//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G110), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n192), .B(G119), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G128), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n191), .B(new_n193), .C1(new_n196), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT23), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n195), .A3(new_n194), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n205), .A2(KEYINPUT74), .A3(new_n191), .A4(new_n193), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n194), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n191), .A2(KEYINPUT24), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G110), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT72), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(new_n208), .B2(new_n210), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n202), .A2(new_n206), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G125), .B(G140), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT16), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n218));
  INV_X1    g032(.A(G140), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G125), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n217), .A2(G146), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(G125), .ZN(new_n223));
  INV_X1    g037(.A(G125), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G140), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT75), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(new_n222), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G953), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(G221), .A3(G234), .ZN(new_n234));
  XOR2_X1   g048(.A(new_n234), .B(KEYINPUT22), .Z(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G137), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n234), .B(KEYINPUT22), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n205), .A2(new_n193), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G110), .ZN(new_n243));
  OR3_X1    g057(.A1(new_n212), .A2(new_n213), .A3(new_n207), .ZN(new_n244));
  AOI21_X1  g058(.A(G146), .B1(new_n217), .B2(new_n220), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n243), .B(new_n244), .C1(new_n245), .C2(new_n221), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n232), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT77), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT76), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n240), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n236), .A2(new_n239), .A3(KEYINPUT76), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n232), .A2(new_n246), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT77), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n232), .A2(new_n241), .A3(new_n255), .A4(new_n246), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n248), .A2(new_n254), .A3(new_n188), .A4(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT78), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT25), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(KEYINPUT77), .A2(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n261));
  INV_X1    g075(.A(new_n259), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n261), .A2(new_n188), .A3(new_n262), .A4(new_n256), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n190), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n256), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n265), .A2(G902), .A3(new_n189), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n230), .A2(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n230), .A2(G143), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G146), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .A4(G128), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n269), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(G137), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(G137), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n283), .A2(new_n284), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n282), .A2(G137), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n238), .A2(G134), .ZN(new_n289));
  OAI21_X1  g103(.A(G131), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n274), .A2(new_n276), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n192), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(new_n278), .A3(KEYINPUT67), .A4(new_n271), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n280), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT0), .B(G128), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n272), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n192), .A2(KEYINPUT0), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT0), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G128), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n293), .A2(new_n303), .A3(KEYINPUT64), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n283), .A2(new_n286), .A3(new_n284), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G131), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n287), .ZN(new_n308));
  AND4_X1   g122(.A1(KEYINPUT0), .A2(new_n274), .A3(new_n276), .A4(G128), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n296), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n198), .ZN(new_n314));
  NAND2_X1  g128(.A1(G116), .A2(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT2), .A2(G113), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT2), .A2(G113), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n314), .B(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n320));
  INV_X1    g134(.A(G113), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(G116), .A2(G119), .ZN(new_n323));
  NOR2_X1   g137(.A1(G116), .A2(G119), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n322), .B(new_n316), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n319), .A2(new_n325), .A3(KEYINPUT66), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT66), .B1(new_n319), .B2(new_n325), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n312), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n296), .A2(new_n311), .A3(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT28), .ZN(new_n333));
  INV_X1    g147(.A(G237), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n233), .A3(G210), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT27), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT26), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n335), .A2(KEYINPUT27), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(KEYINPUT27), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n341), .A3(G101), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G101), .B1(new_n337), .B2(new_n341), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n331), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n333), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n188), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n293), .A2(new_n192), .B1(KEYINPUT1), .B2(new_n270), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n291), .B1(new_n278), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT65), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n311), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n309), .B1(new_n299), .B2(new_n304), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT65), .A3(new_n308), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n328), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n331), .B1(new_n359), .B2(KEYINPUT69), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT69), .ZN(new_n361));
  AOI211_X1 g175(.A(new_n361), .B(new_n328), .C1(new_n356), .C2(new_n358), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT28), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT68), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n343), .B2(new_n344), .ZN(new_n365));
  INV_X1    g179(.A(new_n344), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT68), .A3(new_n342), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n350), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n296), .A2(new_n311), .A3(KEYINPUT30), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n357), .A2(KEYINPUT65), .A3(new_n308), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT65), .B1(new_n357), .B2(new_n308), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n373), .A2(new_n374), .A3(new_n354), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n329), .B(new_n372), .C1(new_n375), .C2(KEYINPUT30), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n331), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n377), .B2(new_n346), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n352), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G472), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT71), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n369), .B1(KEYINPUT28), .B2(new_n332), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n382), .B2(new_n348), .ZN(new_n383));
  INV_X1    g197(.A(new_n368), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n350), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n361), .B1(new_n375), .B2(new_n328), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n311), .A2(new_n355), .ZN(new_n387));
  INV_X1    g201(.A(new_n354), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n358), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT69), .A3(new_n329), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n331), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n385), .B1(new_n391), .B2(KEYINPUT28), .ZN(new_n392));
  INV_X1    g206(.A(new_n331), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n296), .A2(new_n311), .A3(KEYINPUT30), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n393), .B1(new_n396), .B2(new_n329), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n347), .B1(new_n397), .B2(new_n345), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n383), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G472), .ZN(new_n401));
  NOR2_X1   g215(.A1(G472), .A2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT31), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n397), .B2(new_n345), .ZN(new_n405));
  AND4_X1   g219(.A1(new_n404), .A2(new_n376), .A3(new_n331), .A4(new_n345), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n389), .A2(new_n329), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n393), .B1(new_n408), .B2(new_n361), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n349), .B1(new_n409), .B2(new_n390), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n368), .B1(new_n410), .B2(new_n369), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n403), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n381), .A2(new_n401), .B1(new_n412), .B2(KEYINPUT32), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n376), .A2(new_n331), .A3(new_n345), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT31), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n397), .A2(new_n404), .A3(new_n345), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n384), .B1(new_n363), .B2(new_n350), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n402), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT70), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n422));
  OAI211_X1 g236(.A(KEYINPUT70), .B(new_n402), .C1(new_n417), .C2(new_n418), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n268), .B1(new_n413), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G214), .B1(G237), .B2(G902), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G122), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G104), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT3), .B1(new_n430), .B2(G107), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n432));
  INV_X1    g246(.A(G107), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(G104), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(G107), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(G101), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n326), .B2(new_n327), .ZN(new_n439));
  INV_X1    g253(.A(G101), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n431), .A2(new_n434), .A3(new_n440), .A4(new_n435), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n441), .A2(KEYINPUT4), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n436), .A2(G101), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(KEYINPUT4), .A3(new_n441), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n439), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT5), .B1(new_n323), .B2(new_n324), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n313), .A2(KEYINPUT5), .A3(G119), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(G113), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n325), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n430), .A2(G107), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n433), .A2(G104), .ZN(new_n454));
  OAI21_X1  g268(.A(G101), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n441), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n429), .B1(new_n448), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n438), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n319), .A2(new_n325), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n319), .A2(new_n325), .A3(KEYINPUT66), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n443), .B1(new_n442), .B2(new_n444), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n457), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n428), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n357), .A2(new_n224), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n273), .A2(new_n279), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n224), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n353), .A2(new_n278), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT84), .B1(new_n475), .B2(G125), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(G224), .A3(new_n233), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n233), .A2(G224), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n471), .A2(new_n479), .A3(new_n474), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n482), .B(new_n429), .C1(new_n448), .C2(new_n457), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n470), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n470), .A2(new_n481), .A3(KEYINPUT85), .A4(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n479), .A2(KEYINPUT7), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n477), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n471), .A2(new_n474), .A3(new_n476), .A4(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n428), .B(KEYINPUT8), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n452), .A2(new_n456), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n457), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n469), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n188), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n427), .B1(new_n488), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n427), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n503), .B(new_n500), .C1(new_n486), .C2(new_n487), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n426), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n506));
  INV_X1    g320(.A(new_n456), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n475), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n472), .A2(new_n456), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n506), .B1(new_n510), .B2(new_n308), .ZN(new_n511));
  INV_X1    g325(.A(new_n308), .ZN(new_n512));
  AOI211_X1 g326(.A(KEYINPUT12), .B(new_n512), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n357), .B(new_n438), .C1(new_n465), .C2(new_n466), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT10), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n280), .A2(KEYINPUT10), .A3(new_n507), .A4(new_n295), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n515), .A2(new_n512), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(G110), .B(G140), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n233), .A2(G227), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT83), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT83), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n514), .A2(new_n519), .A3(new_n526), .A4(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n357), .A2(new_n438), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n445), .B2(new_n447), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n517), .A2(new_n518), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n308), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n519), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n525), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G469), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n188), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n519), .A2(new_n531), .A3(new_n523), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n523), .B1(new_n514), .B2(new_n519), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(KEYINPUT82), .B(G469), .C1(new_n539), .C2(G902), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n519), .A2(new_n531), .A3(new_n523), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n514), .A2(new_n519), .ZN(new_n542));
  OAI211_X1 g356(.A(G469), .B(new_n541), .C1(new_n542), .C2(new_n523), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT82), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n535), .A2(new_n188), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n536), .A2(new_n540), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT9), .B(G234), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT79), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G221), .B1(new_n551), .B2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n334), .A2(new_n233), .A3(G214), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(new_n275), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G131), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n554), .B(G143), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n285), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n221), .A2(new_n245), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n560), .B(new_n561), .C1(new_n559), .C2(new_n556), .ZN(new_n562));
  XNOR2_X1  g376(.A(G113), .B(G122), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(new_n430), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n231), .B1(new_n230), .B2(new_n216), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT18), .A2(G131), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n555), .A2(KEYINPUT87), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT87), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n557), .A2(new_n568), .B1(KEYINPUT18), .B2(G131), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n562), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n564), .B1(new_n562), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n188), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G475), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n556), .A2(new_n558), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n226), .A2(KEYINPUT19), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n227), .A2(new_n229), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n230), .B(new_n577), .C1(new_n578), .C2(KEYINPUT19), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n579), .A3(new_n222), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n580), .A2(new_n570), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n571), .B1(new_n581), .B2(new_n564), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT20), .ZN(new_n583));
  NOR2_X1   g397(.A1(G475), .A2(G902), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n583), .B1(new_n582), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n575), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(G234), .A2(G237), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(G952), .A3(new_n233), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(G902), .A3(G953), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT21), .B(G898), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(G128), .B(G143), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT13), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n192), .A2(KEYINPUT13), .A3(G143), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n282), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n596), .A2(new_n598), .B1(new_n282), .B2(new_n595), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT88), .ZN(new_n600));
  INV_X1    g414(.A(G122), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(KEYINPUT88), .A2(G122), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G116), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n313), .A2(G122), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n605), .A2(new_n433), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n433), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n599), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OR3_X1    g423(.A1(new_n601), .A2(KEYINPUT14), .A3(G116), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(KEYINPUT14), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n313), .B1(new_n602), .B2(new_n603), .ZN(new_n613));
  OAI21_X1  g427(.A(G107), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n595), .B(new_n282), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n433), .A3(new_n606), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n551), .A2(new_n187), .A3(G953), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n609), .A2(new_n619), .A3(new_n617), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G478), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(KEYINPUT15), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n623), .B(new_n625), .Z(new_n626));
  NOR3_X1   g440(.A1(new_n587), .A2(new_n594), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n505), .A2(new_n553), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n425), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G101), .ZN(G3));
  NOR3_X1   g445(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT89), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n488), .A2(new_n427), .A3(new_n501), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT89), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n426), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT90), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT90), .ZN(new_n637));
  INV_X1    g451(.A(new_n426), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n504), .B2(KEYINPUT89), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n488), .A2(new_n501), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n503), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n633), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n637), .B(new_n639), .C1(new_n642), .C2(KEYINPUT89), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n623), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(KEYINPUT93), .A3(new_n624), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT93), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n623), .B2(G478), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n622), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n619), .B1(new_n609), .B2(new_n617), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT91), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(KEYINPUT92), .A3(KEYINPUT33), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT92), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n621), .A2(new_n622), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(KEYINPUT91), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n656), .B2(new_n655), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n654), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n188), .A2(G478), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n650), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n587), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n594), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n188), .B1(new_n417), .B2(new_n418), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n421), .A2(new_n666), .A3(new_n423), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n553), .A2(new_n268), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n645), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT34), .B(G104), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT94), .B(KEYINPUT95), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(new_n587), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n626), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n594), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n645), .A2(new_n669), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT35), .B(G107), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  INV_X1    g494(.A(new_n423), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n369), .B1(new_n391), .B2(KEYINPUT28), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n415), .B(new_n416), .C1(new_n682), .C2(new_n384), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT70), .B1(new_n683), .B2(new_n402), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n260), .A2(new_n263), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n189), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n252), .A2(KEYINPUT36), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n253), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n189), .A2(G902), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n685), .A2(KEYINPUT96), .A3(new_n666), .A4(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n421), .A2(new_n666), .A3(new_n423), .A4(new_n692), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT96), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n693), .A2(new_n696), .A3(new_n629), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT37), .B(G110), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  INV_X1    g513(.A(new_n692), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n413), .B2(new_n424), .ZN(new_n701));
  INV_X1    g515(.A(new_n553), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n701), .A2(new_n702), .A3(new_n643), .A4(new_n636), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT97), .B(G900), .Z(new_n704));
  AOI21_X1  g518(.A(new_n590), .B1(new_n704), .B2(new_n592), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n676), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT98), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n192), .ZN(G30));
  XNOR2_X1  g524(.A(new_n642), .B(KEYINPUT99), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT38), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n705), .B(KEYINPUT39), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n702), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT40), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n683), .A2(KEYINPUT32), .A3(new_n402), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n397), .A2(new_n345), .B1(new_n368), .B2(new_n332), .ZN(new_n717));
  OAI21_X1  g531(.A(G472), .B1(new_n717), .B2(G902), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n424), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n587), .A2(new_n626), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n426), .A3(new_n700), .A4(new_n720), .ZN(new_n721));
  OR3_X1    g535(.A1(new_n712), .A2(new_n715), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G143), .ZN(G45));
  NOR2_X1   g537(.A1(new_n663), .A2(new_n705), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n703), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n230), .ZN(G48));
  NAND2_X1  g541(.A1(new_n534), .A2(new_n188), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n552), .A3(new_n536), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n425), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n636), .A2(new_n643), .A3(new_n664), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT41), .B(G113), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND3_X1  g550(.A1(new_n636), .A2(new_n643), .A3(new_n677), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n313), .ZN(G18));
  NAND2_X1  g553(.A1(new_n701), .A2(new_n627), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n636), .A2(new_n643), .A3(new_n731), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n198), .ZN(G21));
  INV_X1    g557(.A(new_n266), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT100), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n687), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT100), .B1(new_n264), .B2(new_n266), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n382), .A2(new_n384), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n402), .B1(new_n417), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n666), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n751), .A2(new_n594), .A3(new_n730), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n643), .A3(new_n636), .A4(new_n720), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT101), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  AND4_X1   g569(.A1(new_n666), .A2(new_n724), .A3(new_n692), .A4(new_n750), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n636), .A2(new_n643), .A3(new_n756), .A4(new_n731), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  OAI21_X1  g572(.A(KEYINPUT102), .B1(new_n537), .B2(new_n538), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT102), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n541), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(G469), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n536), .A2(new_n546), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT103), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n536), .A2(new_n762), .A3(KEYINPUT103), .A4(new_n546), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n502), .A2(new_n504), .A3(new_n638), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(new_n768), .A3(new_n552), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n425), .A3(new_n724), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n771));
  INV_X1    g585(.A(new_n748), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n419), .A2(new_n422), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n716), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n774), .A2(KEYINPUT105), .B1(new_n401), .B2(new_n381), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT105), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n776), .A3(new_n716), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n772), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n552), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n765), .B2(new_n766), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n780), .A2(new_n768), .A3(new_n781), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n770), .A2(new_n771), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n285), .ZN(G33));
  NAND3_X1  g598(.A1(new_n769), .A2(new_n425), .A3(new_n706), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  OAI21_X1  g600(.A(G469), .B1(new_n539), .B2(KEYINPUT45), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n759), .A2(new_n761), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(KEYINPUT45), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n545), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT46), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n536), .B1(new_n790), .B2(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n552), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n713), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n667), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n675), .A2(new_n662), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT43), .Z(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n799), .A3(new_n692), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT44), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n796), .A2(new_n768), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT106), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(new_n238), .ZN(G39));
  XNOR2_X1  g618(.A(new_n793), .B(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n413), .A2(new_n424), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n768), .A2(new_n268), .A3(new_n724), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  NOR3_X1   g623(.A1(new_n798), .A2(new_n638), .A3(new_n779), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n729), .A2(new_n536), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n810), .B(new_n748), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT107), .Z(new_n815));
  AOI21_X1  g629(.A(new_n719), .B1(new_n813), .B2(new_n812), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n712), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n799), .A2(new_n590), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n731), .A2(new_n768), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n778), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT48), .Z(new_n823));
  AOI21_X1  g637(.A(KEYINPUT115), .B1(new_n233), .B2(G952), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n719), .A2(new_n819), .A3(new_n268), .A4(new_n589), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n825), .A2(new_n587), .A3(new_n662), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n824), .B(new_n826), .C1(KEYINPUT115), .C2(new_n233), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n818), .A2(new_n730), .A3(new_n751), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n645), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT116), .Z(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n712), .A2(new_n638), .A3(new_n828), .ZN(new_n832));
  NOR2_X1   g646(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n662), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n825), .A2(new_n675), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n666), .A2(new_n692), .A3(new_n750), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n820), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n805), .B1(new_n552), .B2(new_n811), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n818), .A2(new_n638), .A3(new_n642), .A4(new_n751), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n834), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n831), .B1(new_n847), .B2(KEYINPUT51), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n846), .B2(new_n850), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n806), .A2(new_n702), .A3(new_n692), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n644), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n636), .A2(new_n643), .A3(new_n720), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n692), .A2(new_n705), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n719), .A2(new_n780), .A3(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n857), .A2(new_n724), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n643), .A2(new_n636), .A3(new_n731), .A4(new_n756), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n857), .B2(new_n706), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n719), .A2(new_n780), .A3(new_n860), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n703), .A2(new_n725), .B1(new_n866), .B2(new_n858), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n757), .B1(new_n703), .B2(new_n707), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n587), .A2(new_n626), .A3(new_n705), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n641), .A2(new_n426), .A3(new_n872), .A4(new_n633), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT109), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n768), .A2(KEYINPUT109), .A3(new_n872), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n701), .A2(new_n875), .A3(new_n702), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n769), .A2(new_n756), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n785), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n783), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n505), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n594), .B1(new_n676), .B2(new_n663), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n667), .A2(new_n668), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n697), .A2(new_n630), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT108), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n697), .A2(new_n630), .A3(new_n883), .A4(KEYINPUT108), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n753), .B1(new_n741), .B2(new_n740), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n732), .B1(new_n733), .B2(new_n737), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n880), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n855), .B1(new_n871), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n880), .A2(new_n888), .A3(new_n891), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT52), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n869), .B1(new_n867), .B2(new_n868), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(KEYINPUT53), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n902), .B2(KEYINPUT110), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT110), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n901), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n854), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(G952), .A2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n817), .B1(new_n907), .B2(new_n908), .ZN(G75));
  NOR2_X1   g723(.A1(new_n233), .A2(G952), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(G210), .A2(G902), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n899), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n481), .B(KEYINPUT55), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT118), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n470), .A2(new_n483), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT117), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n915), .B(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n918), .A2(KEYINPUT56), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n911), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n899), .A2(KEYINPUT119), .A3(new_n912), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT119), .B1(new_n899), .B2(new_n912), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT120), .B(new_n918), .C1(new_n923), .C2(new_n924), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n920), .B1(new_n927), .B2(new_n928), .ZN(G51));
  NOR2_X1   g743(.A1(new_n902), .A2(new_n900), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n545), .B(KEYINPUT57), .Z(new_n931));
  OAI21_X1  g745(.A(new_n534), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n899), .A2(G902), .A3(new_n789), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n910), .B1(new_n932), .B2(new_n933), .ZN(G54));
  NAND4_X1  g748(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n935));
  INV_X1    g749(.A(new_n582), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(KEYINPUT121), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(KEYINPUT121), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n911), .B1(new_n935), .B2(new_n936), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G60));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT59), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n654), .B(new_n943), .C1(new_n657), .C2(new_n659), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n911), .B1(new_n930), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n903), .A2(new_n906), .A3(new_n943), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(new_n660), .ZN(G63));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n187), .A2(new_n188), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n899), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n951), .ZN(new_n953));
  AOI211_X1 g767(.A(KEYINPUT123), .B(new_n953), .C1(new_n893), .C2(new_n898), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n689), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n871), .A2(new_n855), .A3(new_n892), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT53), .B1(new_n894), .B2(new_n897), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT123), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n899), .A2(new_n948), .A3(new_n951), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n265), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n955), .A2(new_n961), .A3(new_n911), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n955), .A2(new_n961), .A3(KEYINPUT61), .A4(new_n911), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(G66));
  AND2_X1   g780(.A1(new_n888), .A2(new_n891), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n233), .ZN(new_n968));
  INV_X1    g782(.A(new_n593), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(G224), .A3(G953), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n917), .B1(G898), .B2(new_n233), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G69));
  AOI21_X1  g789(.A(new_n233), .B1(G227), .B2(G900), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n808), .A2(new_n785), .A3(new_n802), .ZN(new_n977));
  INV_X1    g791(.A(new_n783), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n868), .A2(new_n726), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n795), .A2(new_n858), .A3(new_n821), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n396), .B(KEYINPUT125), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n577), .B1(new_n578), .B2(KEYINPUT19), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n983), .B(new_n984), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n233), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n976), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n714), .B1(new_n663), .B2(new_n676), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n989), .A2(new_n425), .A3(new_n768), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n808), .A2(new_n802), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n722), .A2(new_n979), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(KEYINPUT62), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n994));
  AOI21_X1  g808(.A(G953), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n988), .B1(new_n995), .B2(new_n985), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n988), .B(KEYINPUT126), .C1(new_n995), .C2(new_n985), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g814(.A(KEYINPUT127), .B(G900), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n985), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n976), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1000), .A2(new_n1003), .ZN(G72));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n982), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n967), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n397), .A2(new_n346), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n911), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n993), .A2(new_n967), .A3(new_n994), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n346), .B(new_n397), .C1(new_n1012), .C2(new_n1006), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n377), .A2(new_n346), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1007), .B1(new_n1014), .B2(new_n414), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n899), .A2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1011), .A2(new_n1013), .A3(new_n1016), .ZN(G57));
endmodule


