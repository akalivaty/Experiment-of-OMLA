//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n187));
  OAI21_X1  g001(.A(G214), .B1(G237), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT87), .Z(new_n189));
  XNOR2_X1  g003(.A(G143), .B(G146), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  OAI211_X1 g006(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n192), .C2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT67), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n191), .B1(new_n194), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n190), .A2(new_n199), .A3(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT0), .B(G128), .Z(new_n203));
  NAND3_X1  g017(.A1(new_n191), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT0), .B(G128), .C1(new_n190), .C2(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT75), .B(G125), .ZN(new_n208));
  MUX2_X1   g022(.A(new_n201), .B(new_n207), .S(new_n208), .Z(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G224), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n209), .B(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT81), .B(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  AOI21_X1  g028(.A(G101), .B1(new_n213), .B2(G107), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT82), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n214), .A2(new_n215), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(KEYINPUT81), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G104), .ZN(new_n226));
  AOI21_X1  g040(.A(G107), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT84), .B1(new_n228), .B2(G104), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT84), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n216), .A3(G107), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n223), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n236));
  INV_X1    g050(.A(G113), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(G119), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT5), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n236), .A2(new_n241), .B1(new_n243), .B2(new_n235), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n234), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT89), .ZN(new_n246));
  XNOR2_X1  g060(.A(G110), .B(G122), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n248));
  INV_X1    g062(.A(G101), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n228), .A2(G104), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n220), .A2(KEYINPUT82), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n225), .A2(G104), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n216), .A2(KEYINPUT81), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n228), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n253), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n224), .A2(new_n226), .A3(G107), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n260));
  OAI22_X1  g074(.A1(new_n227), .A2(new_n220), .B1(new_n260), .B2(new_n250), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n249), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT83), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n222), .B(new_n258), .C1(new_n227), .C2(new_n220), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G101), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT4), .A4(new_n223), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n270), .A3(G101), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n243), .B1(new_n272), .B2(new_n235), .ZN(new_n273));
  INV_X1    g087(.A(G119), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G116), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n242), .B(KEYINPUT68), .C1(new_n239), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n248), .B1(new_n269), .B2(new_n279), .ZN(new_n280));
  AOI211_X1 g094(.A(KEYINPUT88), .B(new_n278), .C1(new_n264), .C2(new_n268), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n246), .B(new_n247), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n246), .B1(new_n280), .B2(new_n281), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n247), .B(KEYINPUT90), .Z(new_n284));
  AOI22_X1  g098(.A1(new_n282), .A2(KEYINPUT6), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n283), .A2(KEYINPUT6), .A3(new_n284), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n212), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n209), .B(new_n288), .Z(new_n289));
  XNOR2_X1  g103(.A(new_n234), .B(new_n244), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n247), .B(KEYINPUT8), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n292), .B2(new_n282), .ZN(new_n293));
  OAI21_X1  g107(.A(G210), .B1(G237), .B2(G902), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n287), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n287), .B2(new_n293), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n189), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT15), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G478), .ZN(new_n299));
  AND2_X1   g113(.A1(KEYINPUT65), .A2(G134), .ZN(new_n300));
  NOR2_X1   g114(.A1(KEYINPUT65), .A2(G134), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n192), .A2(G128), .ZN(new_n303));
  INV_X1    g117(.A(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G143), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT96), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n303), .B2(new_n305), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n192), .A2(KEYINPUT13), .A3(G128), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT95), .A3(new_n305), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT13), .B1(new_n192), .B2(G128), .ZN(new_n313));
  OAI221_X1 g127(.A(G134), .B1(KEYINPUT95), .B2(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G122), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT94), .B1(new_n315), .B2(G116), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n238), .A3(G122), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n238), .A2(G122), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n320), .A2(G107), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n321), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n228), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n310), .B(new_n314), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT9), .B(G234), .ZN(new_n326));
  INV_X1    g140(.A(G217), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n326), .A2(new_n327), .A3(G953), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT14), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n316), .B2(new_n318), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT97), .B1(new_n330), .B2(new_n321), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n320), .A2(new_n329), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n330), .A2(KEYINPUT97), .A3(new_n321), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n228), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n309), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT65), .B(G134), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n307), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n310), .ZN(new_n339));
  INV_X1    g153(.A(new_n322), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n325), .B(new_n328), .C1(new_n335), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT98), .ZN(new_n343));
  INV_X1    g157(.A(new_n341), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n334), .A2(new_n332), .A3(new_n331), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G107), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT98), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n325), .A4(new_n328), .ZN(new_n349));
  INV_X1    g163(.A(new_n328), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n341), .B1(G107), .B2(new_n345), .ZN(new_n351));
  INV_X1    g165(.A(new_n325), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n343), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G902), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n299), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n355), .A3(new_n299), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(KEYINPUT99), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT99), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n354), .A2(new_n355), .A3(new_n299), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(new_n356), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n210), .A2(G952), .ZN(new_n363));
  NAND2_X1  g177(.A1(G234), .A2(G237), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT21), .B(G898), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(G902), .A3(G953), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G237), .A2(G953), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(G143), .A3(G214), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(G143), .B1(new_n370), .B2(G214), .ZN(new_n373));
  OAI21_X1  g187(.A(G131), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  INV_X1    g189(.A(G131), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n371), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT17), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT16), .ZN(new_n380));
  AND2_X1   g194(.A1(KEYINPUT75), .A2(G125), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT75), .A2(G125), .ZN(new_n382));
  OAI21_X1  g196(.A(G140), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G125), .A2(G140), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n380), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G140), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n208), .A2(new_n380), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n195), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n208), .A2(new_n380), .A3(new_n387), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n384), .B1(new_n208), .B2(G140), .ZN(new_n391));
  OAI211_X1 g205(.A(G146), .B(new_n390), .C1(new_n391), .C2(new_n380), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n375), .A2(new_n371), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT17), .A3(G131), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n379), .A2(new_n389), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(G146), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT76), .ZN(new_n398));
  NAND2_X1  g212(.A1(G125), .A2(G140), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n385), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT76), .B1(new_n401), .B2(new_n384), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n397), .B1(new_n403), .B2(new_n195), .ZN(new_n404));
  AOI211_X1 g218(.A(KEYINPUT77), .B(G146), .C1(new_n400), .C2(new_n402), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n396), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n372), .A2(new_n373), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT18), .A2(G131), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT91), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT91), .ZN(new_n411));
  INV_X1    g225(.A(new_n409), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n393), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n409), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n395), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT93), .B(G104), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n420), .B(new_n395), .C1(new_n407), .C2(new_n416), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G475), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n391), .A2(KEYINPUT92), .A3(KEYINPUT19), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n383), .A2(KEYINPUT19), .A3(new_n385), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT19), .B1(new_n400), .B2(new_n402), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n195), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n374), .A2(new_n377), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(new_n392), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n410), .A2(new_n413), .B1(new_n408), .B2(new_n409), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n433), .A2(new_n435), .B1(new_n436), .B2(new_n406), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n423), .B1(new_n437), .B2(new_n420), .ZN(new_n438));
  NOR2_X1   g252(.A1(G475), .A2(G902), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT20), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n442), .A3(new_n439), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n426), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AND4_X1   g258(.A1(new_n359), .A2(new_n362), .A3(new_n369), .A4(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G221), .B1(new_n326), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n271), .A2(new_n207), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n269), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT11), .ZN(new_n451));
  OR2_X1    g265(.A1(KEYINPUT65), .A2(G134), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT65), .A2(G134), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(G137), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G137), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G134), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n451), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT11), .B1(new_n337), .B2(new_n455), .ZN(new_n458));
  OAI21_X1  g272(.A(G131), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n451), .B1(new_n302), .B2(G137), .ZN(new_n460));
  INV_X1    g274(.A(new_n456), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n302), .B2(G137), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n376), .B(new_n460), .C1(new_n462), .C2(new_n451), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n304), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n200), .B1(new_n466), .B2(new_n190), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n223), .A2(new_n233), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n201), .A2(KEYINPUT10), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n223), .A2(new_n233), .ZN(new_n470));
  OAI22_X1  g284(.A1(new_n468), .A2(KEYINPUT10), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n450), .A2(new_n465), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n210), .A2(G227), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT80), .ZN(new_n475));
  XNOR2_X1  g289(.A(G110), .B(G140), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n448), .B1(new_n264), .B2(new_n268), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n464), .B1(new_n478), .B2(new_n471), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n201), .B1(new_n223), .B2(new_n233), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n464), .B1(new_n482), .B2(new_n468), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n223), .A2(new_n233), .A3(new_n467), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n234), .B2(new_n201), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT12), .A3(new_n464), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n477), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n355), .B1(new_n481), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G469), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n483), .A2(new_n484), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT12), .B1(new_n487), .B2(new_n464), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(KEYINPUT86), .A3(new_n488), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n473), .A4(new_n477), .ZN(new_n498));
  INV_X1    g312(.A(new_n477), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n465), .B1(new_n450), .B2(new_n472), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n478), .A2(new_n464), .A3(new_n471), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT85), .B(G469), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n355), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n447), .B1(new_n492), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n445), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n187), .B1(new_n297), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n304), .B2(G119), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n274), .A2(KEYINPUT72), .A3(G128), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n304), .A2(G119), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT24), .B(G110), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n274), .A2(G128), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n304), .A2(KEYINPUT23), .A3(G119), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n274), .A2(G128), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n517), .B(new_n518), .C1(new_n519), .C2(KEYINPUT23), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n516), .B1(G110), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n392), .B(new_n521), .C1(new_n404), .C2(new_n405), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n389), .A2(new_n392), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n514), .A2(new_n515), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT73), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n514), .A2(new_n526), .A3(new_n515), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT74), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n520), .A2(new_n528), .A3(G110), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n520), .B2(G110), .ZN(new_n530));
  OAI22_X1  g344(.A1(new_n525), .A2(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n522), .B1(new_n523), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT22), .B(G137), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n522), .B(new_n535), .C1(new_n523), .C2(new_n531), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n327), .B1(G234), .B2(new_n355), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G902), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT79), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n355), .A3(new_n538), .ZN(new_n545));
  NOR2_X1   g359(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n546), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n537), .A2(new_n355), .A3(new_n538), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n544), .B1(new_n551), .B2(new_n540), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT66), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n337), .A2(new_n554), .A3(new_n455), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n302), .A2(G137), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT66), .B1(new_n455), .B2(G134), .ZN(new_n557));
  OAI211_X1 g371(.A(G131), .B(new_n555), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n463), .A2(new_n201), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n206), .B1(new_n459), .B2(new_n463), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT30), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n300), .A2(new_n301), .A3(new_n455), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT11), .B1(new_n563), .B2(new_n461), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n376), .B1(new_n564), .B2(new_n460), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n457), .A2(new_n458), .A3(G131), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n207), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n463), .A2(new_n201), .A3(new_n558), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n277), .B1(new_n561), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT69), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n277), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n273), .A2(new_n276), .A3(KEYINPUT69), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n567), .A2(new_n574), .A3(new_n568), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n370), .A2(G210), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT27), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT26), .B(G101), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT31), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n570), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n277), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT30), .B1(new_n559), .B2(new_n560), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n567), .A2(new_n562), .A3(new_n568), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT31), .B1(new_n587), .B2(new_n580), .ZN(new_n588));
  INV_X1    g402(.A(new_n579), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT28), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n277), .B1(new_n559), .B2(new_n560), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(new_n575), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n559), .A2(new_n560), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT28), .B1(new_n593), .B2(new_n574), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n589), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n583), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(G472), .A2(G902), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT32), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT70), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT70), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n601), .B(KEYINPUT32), .C1(new_n596), .C2(new_n597), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT29), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n589), .B1(new_n575), .B2(new_n590), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n606), .B2(new_n592), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n579), .B1(new_n570), .B2(new_n575), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT71), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n573), .B(new_n572), .C1(new_n559), .C2(new_n560), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n590), .B1(new_n610), .B2(new_n575), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n606), .A2(new_n611), .A3(new_n604), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(G902), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n591), .A2(new_n575), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n605), .B1(new_n614), .B2(new_n590), .ZN(new_n615));
  INV_X1    g429(.A(new_n575), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n589), .B1(new_n587), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT71), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n615), .A2(new_n617), .A3(new_n618), .A4(new_n604), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n609), .A2(new_n613), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n596), .A2(new_n597), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n620), .A2(G472), .B1(new_n621), .B2(KEYINPUT32), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n553), .B1(new_n603), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n359), .A2(new_n362), .A3(new_n369), .A4(new_n444), .ZN(new_n624));
  AOI211_X1 g438(.A(G902), .B(new_n504), .C1(new_n498), .C2(new_n502), .ZN(new_n625));
  INV_X1    g439(.A(G469), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n478), .A2(new_n471), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n627), .A2(new_n465), .B1(new_n488), .B2(new_n485), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n480), .B1(new_n628), .B2(new_n477), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n626), .B1(new_n629), .B2(new_n355), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n446), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n294), .ZN(new_n633));
  INV_X1    g447(.A(new_n212), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n282), .A2(KEYINPUT6), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n283), .A2(new_n284), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n283), .A2(KEYINPUT6), .A3(new_n284), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n292), .A2(new_n282), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n355), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n633), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n287), .A2(new_n293), .A3(new_n294), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n632), .A2(new_n644), .A3(KEYINPUT100), .A4(new_n189), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n509), .A2(new_n623), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G101), .ZN(G3));
  INV_X1    g461(.A(new_n188), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n642), .B2(new_n643), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n596), .A2(new_n355), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G472), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n598), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n631), .A2(new_n652), .A3(new_n553), .ZN(new_n653));
  INV_X1    g467(.A(new_n369), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n655));
  AOI21_X1  g469(.A(G478), .B1(new_n354), .B2(new_n355), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n342), .A2(KEYINPUT33), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n328), .B(KEYINPUT101), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n347), .B2(new_n325), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n657), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n659), .B1(new_n351), .B2(new_n352), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n663), .A2(KEYINPUT102), .A3(KEYINPUT33), .A4(new_n342), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT33), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n662), .A2(new_n664), .B1(new_n354), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(G478), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(G902), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n656), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n655), .B1(new_n669), .B2(new_n444), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n662), .A2(new_n664), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n354), .A2(new_n665), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n672), .A3(new_n668), .ZN(new_n673));
  INV_X1    g487(.A(new_n656), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n441), .A2(new_n443), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n425), .B2(new_n424), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT103), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n654), .B1(new_n670), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n649), .A2(new_n653), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G104), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G6));
  XOR2_X1   g497(.A(new_n369), .B(KEYINPUT105), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n444), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n359), .B2(new_n362), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n649), .A2(new_n653), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  NAND2_X1  g503(.A1(new_n551), .A2(new_n540), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n536), .A2(KEYINPUT36), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n532), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n532), .A2(new_n691), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n543), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n652), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n509), .A2(new_n645), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  OAI211_X1 g515(.A(new_n696), .B(new_n446), .C1(new_n625), .C2(new_n630), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n603), .B2(new_n622), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n365), .B(KEYINPUT107), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n707));
  OR3_X1    g521(.A1(new_n368), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n444), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n359), .B2(new_n362), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n703), .A2(new_n649), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  XNOR2_X1  g527(.A(new_n709), .B(KEYINPUT39), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n507), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n715), .B(KEYINPUT40), .Z(new_n716));
  INV_X1    g530(.A(new_n600), .ZN(new_n717));
  INV_X1    g531(.A(new_n602), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n596), .A2(KEYINPUT32), .A3(new_n597), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n587), .A2(new_n616), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n589), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n610), .A2(new_n575), .A3(new_n589), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n355), .ZN(new_n723));
  OAI21_X1  g537(.A(G472), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n717), .A2(new_n718), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n444), .B1(new_n359), .B2(new_n362), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n696), .A2(new_n648), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n716), .A2(new_n726), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n644), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n192), .ZN(G45));
  NAND3_X1  g547(.A1(new_n675), .A2(new_n677), .A3(new_n709), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n703), .A2(new_n649), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G146), .ZN(G48));
  AOI21_X1  g551(.A(G902), .B1(new_n498), .B2(new_n502), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n506), .B(new_n446), .C1(new_n626), .C2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n623), .A2(new_n649), .A3(new_n679), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND4_X1  g557(.A1(new_n623), .A2(new_n649), .A3(new_n686), .A4(new_n740), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  NAND2_X1  g559(.A1(new_n603), .A2(new_n622), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n624), .A2(new_n697), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n649), .A2(new_n746), .A3(new_n740), .A4(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT109), .B(G119), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G21));
  AND2_X1   g564(.A1(new_n498), .A2(new_n502), .ZN(new_n751));
  OAI21_X1  g565(.A(G469), .B1(new_n751), .B2(G902), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n446), .A3(new_n506), .A4(new_n684), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n589), .B1(new_n611), .B2(new_n594), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n588), .A3(KEYINPUT110), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n583), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT110), .B1(new_n754), .B2(new_n588), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n597), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n552), .A3(new_n651), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n649), .A3(new_n727), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n651), .A3(new_n696), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n734), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n649), .A2(new_n764), .A3(new_n740), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n734), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n620), .A2(G472), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n598), .A2(new_n599), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n719), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n552), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n642), .A2(new_n507), .A3(new_n643), .A4(new_n188), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT111), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n642), .A2(new_n507), .A3(new_n643), .A4(new_n188), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n553), .B1(new_n622), .B2(new_n770), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n768), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n623), .A3(new_n735), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n774), .A2(new_n778), .B1(new_n779), .B2(new_n767), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n376), .ZN(G33));
  NAND3_X1  g595(.A1(new_n775), .A2(new_n623), .A3(new_n711), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  INV_X1    g597(.A(new_n629), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n784), .A2(KEYINPUT45), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(KEYINPUT45), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(G469), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(G469), .A2(G902), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n788), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n506), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n446), .A3(new_n714), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n793), .A2(new_n446), .A3(new_n714), .A4(new_n795), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n675), .A2(new_n444), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT43), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n697), .B1(new_n651), .B2(new_n598), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT44), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n295), .A2(new_n296), .A3(new_n648), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n802), .A2(KEYINPUT44), .A3(new_n803), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(KEYINPUT115), .B(new_n807), .C1(new_n810), .C2(new_n811), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n799), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(new_n455), .ZN(G39));
  NAND2_X1  g631(.A1(new_n793), .A2(new_n446), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT47), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n793), .A2(KEYINPUT47), .A3(new_n446), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n806), .A2(new_n746), .A3(new_n552), .A4(new_n734), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(new_n387), .ZN(G42));
  NAND2_X1  g639(.A1(new_n752), .A2(new_n506), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT49), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n603), .A2(new_n552), .A3(new_n725), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n189), .A2(new_n446), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n827), .A2(new_n800), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n731), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n731), .A2(new_n648), .A3(new_n740), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n834));
  INV_X1    g648(.A(new_n704), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n802), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n759), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n833), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT50), .Z(new_n840));
  NOR2_X1   g654(.A1(new_n806), .A2(new_n739), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n828), .A2(new_n365), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n843), .A2(new_n677), .A3(new_n675), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n841), .A2(new_n836), .ZN(new_n845));
  INV_X1    g659(.A(new_n763), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n820), .B(new_n821), .C1(new_n446), .C2(new_n826), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n838), .A2(new_n805), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n844), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n840), .A2(KEYINPUT51), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  INV_X1    g666(.A(new_n709), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n694), .B(new_n853), .C1(new_n551), .C2(new_n540), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n726), .A2(new_n507), .A3(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n188), .B(new_n727), .C1(new_n295), .C2(new_n296), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT116), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n854), .B(new_n446), .C1(new_n630), .C2(new_n625), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n603), .B2(new_n725), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n649), .A4(new_n727), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n712), .A2(new_n736), .A3(new_n765), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT52), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n863), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n857), .A2(new_n861), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n357), .A2(new_n358), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n444), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n444), .B2(new_n669), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(new_n684), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n644), .A3(new_n189), .A4(new_n653), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n646), .A2(new_n699), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n774), .A2(new_n778), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n779), .A2(new_n767), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n741), .A2(new_n744), .A3(new_n748), .A4(new_n761), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n710), .A2(new_n870), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n805), .A2(new_n703), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n775), .A2(new_n764), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n782), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n852), .B1(new_n869), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n780), .A2(new_n883), .A3(new_n879), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n868), .A3(new_n864), .A4(new_n875), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n866), .B1(new_n712), .B2(new_n765), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(KEYINPUT53), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n886), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n782), .A2(new_n881), .A3(new_n882), .A4(KEYINPUT53), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n780), .A2(new_n893), .A3(new_n889), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n748), .A2(new_n761), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(KEYINPUT117), .A3(new_n741), .A4(new_n744), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n879), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n894), .A2(new_n899), .A3(new_n875), .ZN(new_n900));
  INV_X1    g714(.A(new_n869), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n900), .A2(new_n901), .B1(new_n888), .B2(new_n852), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n892), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT51), .B1(new_n840), .B2(new_n850), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n845), .A2(new_n777), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT48), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n670), .A2(new_n678), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n843), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n838), .A2(new_n649), .A3(new_n740), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n908), .A2(new_n363), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  NOR4_X1   g726(.A1(new_n851), .A2(new_n905), .A3(new_n906), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n831), .B1(new_n913), .B2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n902), .A2(new_n355), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n916), .B2(G210), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n285), .A2(new_n286), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n212), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n917), .B(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n210), .A2(G952), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT119), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n921), .A2(new_n924), .ZN(G51));
  NOR3_X1   g739(.A1(new_n902), .A2(new_n355), .A3(new_n787), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n646), .A2(new_n699), .A3(new_n874), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n896), .B2(new_n898), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(new_n868), .A3(new_n864), .A4(new_n894), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n886), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT54), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n904), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n788), .B(KEYINPUT57), .Z(new_n933));
  AOI21_X1  g747(.A(new_n751), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n926), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n930), .B(new_n903), .ZN(new_n937));
  INV_X1    g751(.A(new_n933), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n503), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT120), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n922), .B1(new_n936), .B2(new_n940), .ZN(G54));
  NAND3_X1  g755(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  INV_X1    g756(.A(new_n438), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n922), .ZN(G60));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n666), .B1(new_n905), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n666), .A2(new_n949), .ZN(new_n951));
  AOI211_X1 g765(.A(new_n924), .B(new_n950), .C1(new_n932), .C2(new_n951), .ZN(G63));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n930), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g771(.A(KEYINPUT121), .B(new_n955), .C1(new_n886), .C2(new_n929), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n924), .B1(new_n959), .B2(new_n539), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n692), .A2(new_n693), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT122), .Z(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n957), .B2(new_n958), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n960), .B(new_n963), .C1(new_n964), .C2(KEYINPUT61), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT121), .B1(new_n902), .B2(new_n955), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n930), .A2(new_n953), .A3(new_n956), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n539), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n963), .A2(new_n968), .A3(new_n923), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n964), .A3(new_n923), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n965), .A2(new_n972), .ZN(G66));
  AOI21_X1  g787(.A(new_n210), .B1(new_n367), .B2(G224), .ZN(new_n974));
  INV_X1    g788(.A(new_n879), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n875), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n976), .B2(new_n210), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n918), .B1(G898), .B2(new_n210), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n977), .B(new_n978), .Z(G69));
  NOR2_X1   g793(.A1(new_n561), .A2(new_n569), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n432), .B(KEYINPUT124), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n732), .B2(new_n863), .ZN(new_n984));
  OAI211_X1 g798(.A(KEYINPUT62), .B(new_n865), .C1(new_n729), .C2(new_n731), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n824), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n987));
  INV_X1    g801(.A(new_n816), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n872), .A2(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n872), .A2(KEYINPUT125), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n989), .A2(new_n507), .A3(new_n714), .A4(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n623), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n992), .A3(new_n806), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n987), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n816), .A2(KEYINPUT126), .A3(new_n993), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n986), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n982), .B1(new_n997), .B2(new_n210), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n210), .B1(G227), .B2(G900), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n982), .B1(new_n705), .B2(new_n210), .ZN(new_n1000));
  INV_X1    g814(.A(new_n799), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n649), .A2(new_n777), .A3(new_n727), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n780), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n782), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n822), .B2(new_n823), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1003), .A2(new_n865), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(new_n816), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1000), .B1(new_n1007), .B2(new_n210), .ZN(new_n1008));
  OR3_X1    g822(.A1(new_n998), .A2(new_n999), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n999), .B1(new_n998), .B2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(G72));
  INV_X1    g825(.A(new_n976), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1012), .B(new_n986), .C1(new_n995), .C2(new_n996), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n721), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n720), .A2(new_n589), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1006), .A2(new_n816), .A3(new_n976), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1015), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1020), .A2(new_n721), .A3(new_n1022), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n922), .B1(new_n891), .B2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1017), .A2(new_n1018), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1027));
  INV_X1    g841(.A(new_n721), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1029));
  OAI21_X1  g843(.A(KEYINPUT127), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1026), .A2(new_n1030), .ZN(G57));
endmodule


