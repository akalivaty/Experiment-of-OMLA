//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(KEYINPUT2), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT74), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n210), .B1(new_n204), .B2(KEYINPUT2), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n204), .A2(new_n210), .A3(KEYINPUT2), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n202), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT73), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n204), .A2(KEYINPUT72), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT73), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT72), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(G155gat), .A3(G162gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n215), .A2(new_n216), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n209), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223));
  INV_X1    g022(.A(G113gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G120gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(G120gat), .ZN(new_n226));
  INV_X1    g025(.A(G120gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT68), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n231));
  INV_X1    g030(.A(G134gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G127gat), .ZN(new_n233));
  INV_X1    g032(.A(G127gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G134gat), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n225), .A2(new_n228), .A3(new_n237), .A4(new_n226), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n230), .A2(new_n231), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n235), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(KEYINPUT1), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n222), .A2(KEYINPUT3), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n213), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n203), .B1(new_n244), .B2(new_n211), .ZN(new_n245));
  INV_X1    g044(.A(new_n221), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n245), .A2(new_n246), .B1(new_n203), .B2(new_n208), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT76), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n229), .A2(KEYINPUT68), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n238), .A2(new_n231), .A3(new_n236), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n242), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n251), .B1(new_n254), .B2(new_n222), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n247), .A2(KEYINPUT76), .A3(new_n239), .A4(new_n242), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(KEYINPUT4), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT78), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n254), .A2(new_n222), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n257), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n258), .B1(new_n257), .B2(new_n261), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n250), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G225gat), .A2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT39), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n254), .A2(new_n222), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n255), .A2(new_n256), .A3(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n270), .A2(new_n266), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n267), .B(new_n273), .C1(new_n272), .C2(new_n271), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n264), .A2(new_n268), .A3(new_n266), .ZN(new_n275));
  XNOR2_X1  g074(.A(G1gat), .B(G29gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT0), .ZN(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G85gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  AND3_X1   g078(.A1(new_n275), .A2(KEYINPUT81), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT81), .B1(new_n275), .B2(new_n279), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n274), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT40), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n274), .B(KEYINPUT40), .C1(new_n280), .C2(new_n281), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G226gat), .ZN(new_n290));
  INV_X1    g089(.A(G233gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT24), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G183gat), .ZN(new_n298));
  INV_X1    g097(.A(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT24), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT23), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n297), .A2(new_n302), .A3(new_n304), .A4(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n293), .B1(new_n308), .B2(KEYINPUT64), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n307), .A2(new_n304), .A3(new_n295), .A4(new_n296), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n300), .A2(KEYINPUT24), .A3(new_n301), .ZN(new_n311));
  OAI211_X1 g110(.A(KEYINPUT64), .B(new_n293), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT27), .B(G183gat), .Z(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(G190gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT27), .B(G183gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n299), .C1(KEYINPUT65), .C2(KEYINPUT28), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT66), .A4(KEYINPUT26), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT66), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT26), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n296), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n301), .B(new_n320), .C1(new_n321), .C2(new_n323), .ZN(new_n324));
  OAI22_X1  g123(.A1(new_n309), .A2(new_n313), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n292), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(KEYINPUT22), .B2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G211gat), .B(G218gat), .Z(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n324), .B1(new_n316), .B2(new_n318), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT64), .B1(new_n310), .B2(new_n311), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT25), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n338), .B2(new_n312), .ZN(new_n339));
  INV_X1    g138(.A(new_n292), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n327), .A2(new_n335), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n292), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n334), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n289), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n335), .B1(new_n327), .B2(new_n341), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n334), .A3(new_n344), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(KEYINPUT30), .A3(new_n348), .A4(new_n288), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n348), .A3(new_n288), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n351), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n266), .B1(new_n243), .B2(new_n249), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n262), .B2(new_n263), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT4), .B1(new_n255), .B2(new_n256), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n259), .A2(new_n260), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n358), .B1(new_n270), .B2(new_n266), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g165(.A(KEYINPUT77), .B(new_n358), .C1(new_n270), .C2(new_n266), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n360), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n279), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n356), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n284), .A2(new_n285), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n334), .A2(new_n326), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n247), .B1(new_n374), .B2(new_n248), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n334), .B1(new_n249), .B2(new_n326), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(G228gat), .A3(G233gat), .ZN(new_n378));
  INV_X1    g177(.A(G228gat), .ZN(new_n379));
  OAI22_X1  g178(.A1(new_n375), .A2(new_n376), .B1(new_n379), .B2(new_n291), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n373), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n373), .A3(new_n380), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G78gat), .B(G106gat), .Z(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT31), .B(G50gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n381), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n382), .A2(new_n388), .A3(new_n383), .A4(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n360), .B(new_n279), .C1(new_n366), .C2(new_n367), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n370), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n368), .A2(KEYINPUT6), .A3(new_n369), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT37), .B1(new_n348), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n347), .A2(new_n348), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n401), .B2(new_n398), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n289), .B(new_n403), .C1(new_n400), .C2(KEYINPUT37), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n351), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT37), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n346), .B1(new_n406), .B2(new_n288), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n400), .A2(KEYINPUT37), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n392), .B1(new_n397), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n254), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n325), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G227gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n291), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n339), .A2(new_n254), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT69), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT69), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n413), .A2(new_n416), .A3(new_n419), .A4(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT32), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G15gat), .B(G43gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n428), .A2(KEYINPUT70), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(KEYINPUT70), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(KEYINPUT33), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(KEYINPUT32), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n416), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n414), .B2(new_n291), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n436), .B(KEYINPUT34), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n429), .A2(new_n437), .A3(new_n433), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT36), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT36), .ZN(new_n442));
  INV_X1    g241(.A(new_n440), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n437), .B1(new_n429), .B2(new_n433), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n372), .A2(new_n411), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n395), .A2(new_n396), .ZN(new_n447));
  INV_X1    g246(.A(new_n356), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT79), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT79), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n450), .B(new_n356), .C1(new_n395), .C2(new_n396), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n392), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n390), .A2(new_n391), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n439), .A3(new_n440), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n447), .A2(new_n448), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT35), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n450), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n440), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(new_n392), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n447), .A2(KEYINPUT79), .A3(new_n448), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n457), .B1(new_n462), .B2(KEYINPUT35), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n465));
  OR2_X1    g264(.A1(G43gat), .A2(G50gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(G43gat), .A2(G50gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  NAND2_X1  g268(.A1(G29gat), .A2(G36gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(new_n471), .A3(new_n467), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT14), .ZN(new_n476));
  INV_X1    g275(.A(G29gat), .ZN(new_n477));
  INV_X1    g276(.A(G36gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n480));
  NOR3_X1   g279(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n475), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n473), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(KEYINPUT86), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n474), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n469), .B1(new_n489), .B2(new_n470), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n465), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n474), .B1(new_n481), .B2(KEYINPUT86), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n479), .A2(new_n486), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n470), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(KEYINPUT15), .A3(new_n468), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n496));
  NOR2_X1   g295(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n482), .B1(new_n497), .B2(new_n478), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n474), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n468), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n472), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n501), .A3(KEYINPUT17), .ZN(new_n502));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503));
  INV_X1    g302(.A(G1gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT16), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(G1gat), .B2(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G8gat), .ZN(new_n508));
  INV_X1    g307(.A(G8gat), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n506), .B(new_n509), .C1(G1gat), .C2(new_n503), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n502), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n501), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n510), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n512), .A2(KEYINPUT18), .A3(new_n513), .A4(new_n516), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n513), .B(KEYINPUT13), .Z(new_n521));
  INV_X1    g320(.A(new_n516), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n514), .A2(new_n515), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G169gat), .B(G197gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT12), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n525), .B(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n464), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT8), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n544));
  OR2_X1    g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n541), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G99gat), .B(G106gat), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G99gat), .B(G106gat), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n551), .B(new_n541), .C1(new_n546), .C2(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n491), .A2(new_n502), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT90), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT41), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n485), .A2(new_n490), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(new_n553), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n535), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n556), .A2(KEYINPUT41), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n491), .A2(new_n502), .A3(new_n553), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT8), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(G99gat), .B2(G106gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT91), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n543), .A2(new_n545), .A3(new_n544), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n551), .B1(new_n570), .B2(new_n541), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n549), .B(new_n540), .C1(new_n568), .C2(new_n569), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n514), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n564), .A2(new_n574), .A3(new_n557), .A4(new_n534), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n563), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n575), .ZN(new_n579));
  INV_X1    g378(.A(new_n563), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT93), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  AOI211_X1 g381(.A(new_n582), .B(new_n563), .C1(new_n560), .C2(new_n575), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G71gat), .ZN(new_n588));
  INV_X1    g387(.A(G78gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n591), .B(new_n590), .C1(new_n586), .C2(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n511), .B1(new_n598), .B2(new_n597), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT88), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G183gat), .B(G211gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT89), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n607), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n603), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G230gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n291), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n552), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n597), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n617), .B(new_n618), .C1(new_n571), .C2(new_n572), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n550), .B(new_n552), .C1(new_n616), .C2(new_n597), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT10), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n597), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n573), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n615), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n619), .A2(new_n620), .A3(new_n614), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G120gat), .B(G148gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT95), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n626), .A2(new_n627), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(KEYINPUT96), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n612), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n533), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n447), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n504), .ZN(G1324gat));
  NAND3_X1  g443(.A1(new_n533), .A2(new_n356), .A3(new_n641), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT16), .B(G8gat), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OR3_X1    g447(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(G8gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n646), .B1(new_n645), .B2(new_n648), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(G1325gat));
  NAND2_X1  g451(.A1(new_n445), .A2(new_n441), .ZN(new_n653));
  OAI21_X1  g452(.A(G15gat), .B1(new_n642), .B2(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n459), .A2(G15gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n654), .B1(new_n642), .B2(new_n655), .ZN(G1326gat));
  NOR2_X1   g455(.A1(new_n642), .A2(new_n454), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(G1327gat));
  INV_X1    g458(.A(KEYINPUT45), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n585), .A2(new_n640), .A3(new_n611), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n533), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n447), .A2(G29gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n576), .B(KEYINPUT92), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n581), .B2(new_n583), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT44), .B(new_n667), .C1(new_n453), .C2(new_n463), .ZN(new_n668));
  INV_X1    g467(.A(new_n640), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n531), .ZN(new_n671));
  INV_X1    g470(.A(new_n611), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT97), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n452), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(KEYINPUT98), .B(new_n392), .C1(new_n449), .C2(new_n451), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n446), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n679));
  INV_X1    g478(.A(new_n457), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n585), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n668), .B(new_n674), .C1(new_n682), .C2(KEYINPUT44), .ZN(new_n683));
  OAI21_X1  g482(.A(G29gat), .B1(new_n683), .B2(new_n447), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n533), .A2(KEYINPUT45), .A3(new_n661), .A4(new_n663), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n665), .A2(new_n684), .A3(new_n685), .ZN(G1328gat));
  NOR2_X1   g485(.A1(new_n448), .A2(G36gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n662), .A2(KEYINPUT46), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G36gat), .B1(new_n683), .B2(new_n448), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT46), .B1(new_n662), .B2(new_n688), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(G1329gat));
  INV_X1    g491(.A(G43gat), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(KEYINPUT99), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n683), .B2(new_n653), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n459), .A2(KEYINPUT99), .A3(G43gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n533), .A2(new_n661), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n696), .B1(new_n695), .B2(new_n698), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(G1330gat));
  OAI21_X1  g500(.A(G50gat), .B1(new_n683), .B2(new_n454), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n454), .A2(G50gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n533), .A2(new_n661), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n702), .A2(KEYINPUT48), .A3(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1331gat));
  NAND2_X1  g508(.A1(new_n678), .A2(new_n681), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n612), .A2(new_n669), .A3(new_n671), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n397), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g514(.A1(new_n712), .A2(new_n448), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(G1333gat));
  OR3_X1    g519(.A1(new_n712), .A2(G71gat), .A3(new_n459), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n712), .A2(new_n653), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n588), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT100), .B(KEYINPUT50), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1334gat));
  NOR2_X1   g524(.A1(new_n712), .A2(new_n454), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(new_n589), .ZN(G1335gat));
  NOR2_X1   g526(.A1(new_n671), .A2(new_n611), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n640), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n668), .B(new_n729), .C1(new_n682), .C2(KEYINPUT44), .ZN(new_n730));
  OAI21_X1  g529(.A(G85gat), .B1(new_n730), .B2(new_n447), .ZN(new_n731));
  AND4_X1   g530(.A1(KEYINPUT51), .A2(new_n710), .A3(new_n667), .A4(new_n728), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT51), .B1(new_n682), .B2(new_n728), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT101), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n682), .A2(new_n728), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n447), .A2(new_n669), .A3(G85gat), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT102), .Z(new_n742));
  OAI21_X1  g541(.A(new_n731), .B1(new_n740), .B2(new_n742), .ZN(G1336gat));
  OR2_X1    g542(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n744), .A2(new_n356), .A3(new_n668), .A4(new_n729), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n682), .A2(KEYINPUT51), .A3(new_n728), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n737), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n669), .A2(new_n448), .A3(G92gat), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n745), .A2(G92gat), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  INV_X1    g549(.A(new_n748), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n734), .B2(new_n739), .ZN(new_n752));
  OAI21_X1  g551(.A(G92gat), .B1(new_n730), .B2(new_n448), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n750), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n749), .A2(new_n750), .B1(new_n752), .B2(new_n754), .ZN(G1337gat));
  OAI21_X1  g554(.A(G99gat), .B1(new_n730), .B2(new_n653), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n459), .A2(G99gat), .A3(new_n669), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n740), .B2(new_n757), .ZN(G1338gat));
  NAND4_X1  g557(.A1(new_n744), .A2(new_n392), .A3(new_n668), .A4(new_n729), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n454), .A2(new_n669), .A3(G106gat), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n759), .A2(G106gat), .B1(new_n747), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  INV_X1    g561(.A(new_n760), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n734), .B2(new_n739), .ZN(new_n764));
  OAI21_X1  g563(.A(G106gat), .B1(new_n730), .B2(new_n454), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n762), .ZN(new_n766));
  OAI22_X1  g565(.A1(new_n761), .A2(new_n762), .B1(new_n764), .B2(new_n766), .ZN(G1339gat));
  NOR3_X1   g566(.A1(new_n612), .A2(new_n671), .A3(new_n640), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n770), .B(new_n615), .C1(new_n621), .C2(new_n625), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n632), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n619), .A2(new_n620), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n622), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n614), .B1(new_n775), .B2(new_n624), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n624), .A2(new_n614), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT54), .B1(new_n621), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n776), .A2(new_n778), .A3(KEYINPUT103), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT103), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n615), .B1(new_n573), .B2(new_n623), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n770), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n782), .B2(new_n626), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n773), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n532), .B1(new_n769), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n635), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT103), .B1(new_n776), .B2(new_n778), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(new_n780), .A3(new_n626), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n769), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n523), .ZN(new_n792));
  INV_X1    g591(.A(new_n521), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n516), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n513), .B1(new_n512), .B2(new_n516), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT104), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI211_X1 g596(.A(KEYINPUT104), .B(new_n513), .C1(new_n512), .C2(new_n516), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n530), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT105), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n670), .A2(new_n531), .ZN(new_n802));
  OAI211_X1 g601(.A(KEYINPUT105), .B(new_n530), .C1(new_n797), .C2(new_n798), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n785), .A2(new_n791), .B1(new_n804), .B2(new_n640), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n799), .A2(new_n800), .B1(new_n670), .B2(new_n531), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n784), .A2(new_n769), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n667), .A2(new_n791), .A3(new_n808), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n805), .A2(new_n667), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n768), .B1(new_n810), .B2(new_n672), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n392), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n397), .A2(new_n448), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n459), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n532), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT106), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n808), .A2(new_n671), .A3(new_n791), .ZN(new_n818));
  INV_X1    g617(.A(new_n639), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT96), .B1(new_n633), .B2(new_n635), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n806), .B(new_n803), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n667), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n772), .B1(new_n787), .B2(new_n788), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n578), .A2(new_n584), .B1(new_n823), .B2(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n789), .A2(new_n790), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n635), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n824), .A2(new_n826), .A3(new_n807), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n672), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n768), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n447), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n460), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(KEYINPUT107), .A3(new_n448), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT107), .B1(new_n831), .B2(new_n448), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n224), .B(new_n671), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n834), .ZN(G1340gat));
  OAI211_X1 g634(.A(new_n227), .B(new_n640), .C1(new_n832), .C2(new_n833), .ZN(new_n836));
  OAI21_X1  g635(.A(G120gat), .B1(new_n815), .B2(new_n669), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT108), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n838), .B(new_n839), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n815), .B2(new_n672), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n831), .A2(new_n234), .A3(new_n448), .A4(new_n611), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT109), .Z(G1342gat));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n585), .A2(new_n356), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n232), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT110), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(KEYINPUT110), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n845), .B1(new_n850), .B2(KEYINPUT56), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n848), .A2(KEYINPUT111), .A3(new_n852), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n815), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n232), .B1(new_n855), .B2(new_n667), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n850), .B2(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(G1343gat));
  INV_X1    g657(.A(new_n653), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n813), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n811), .B2(new_n454), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n454), .A2(new_n861), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n768), .B1(new_n828), .B2(KEYINPUT112), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n810), .A2(new_n866), .A3(new_n672), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n864), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n862), .B1(new_n868), .B2(KEYINPUT113), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n870), .B(new_n864), .C1(new_n865), .C2(new_n867), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n671), .B(new_n860), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n653), .A2(new_n392), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT114), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n653), .A2(new_n876), .A3(new_n392), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n830), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  OR4_X1    g677(.A1(G141gat), .A2(new_n878), .A3(new_n356), .A4(new_n532), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT58), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(KEYINPUT115), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n532), .A2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT115), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n830), .A2(new_n884), .A3(new_n875), .A4(new_n877), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n882), .A2(new_n448), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n888), .A3(KEYINPUT116), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n881), .A2(new_n891), .A3(new_n892), .ZN(G1344gat));
  AND2_X1   g692(.A1(new_n882), .A2(new_n885), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n669), .A2(G148gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n448), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G148gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n869), .A2(new_n871), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n859), .A3(new_n813), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n902), .B2(new_n640), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n768), .B(KEYINPUT118), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n807), .B1(new_n809), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n667), .A2(KEYINPUT119), .A3(new_n808), .A4(new_n791), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n822), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT120), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n672), .B1(new_n908), .B2(KEYINPUT120), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT57), .B1(new_n912), .B2(new_n392), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n828), .A2(new_n829), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n863), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n640), .B(new_n860), .C1(new_n913), .C2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n899), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n898), .B1(new_n903), .B2(new_n918), .ZN(G1345gat));
  AOI21_X1  g718(.A(new_n205), .B1(new_n902), .B2(new_n611), .ZN(new_n920));
  AND4_X1   g719(.A1(new_n205), .A2(new_n894), .A3(new_n448), .A4(new_n611), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n920), .A2(new_n921), .ZN(G1346gat));
  OAI211_X1 g721(.A(new_n667), .B(new_n860), .C1(new_n869), .C2(new_n871), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n206), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n924), .B2(new_n923), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n894), .A2(new_n206), .A3(new_n846), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n447), .A2(new_n356), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n459), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n812), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n305), .A3(new_n532), .ZN(new_n932));
  NOR4_X1   g731(.A1(new_n811), .A2(new_n397), .A3(new_n448), .A4(new_n455), .ZN(new_n933));
  AOI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n671), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n932), .A2(new_n934), .ZN(G1348gat));
  OAI21_X1  g734(.A(G176gat), .B1(new_n931), .B2(new_n669), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n306), .A3(new_n640), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT122), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n931), .B2(new_n672), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n672), .A2(new_n315), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n933), .A2(KEYINPUT123), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT123), .B1(new_n933), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n931), .B2(new_n585), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n299), .A3(new_n667), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n950), .B(new_n951), .C1(KEYINPUT61), .C2(new_n949), .ZN(G1351gat));
  NOR4_X1   g751(.A1(new_n811), .A2(new_n397), .A3(new_n448), .A4(new_n874), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT125), .ZN(new_n954));
  INV_X1    g753(.A(G197gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n671), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n859), .A2(new_n929), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n671), .B(new_n957), .C1(new_n913), .C2(new_n916), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G197gat), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n958), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(G1352gat));
  INV_X1    g762(.A(G204gat), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n953), .A2(new_n964), .A3(new_n640), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  INV_X1    g765(.A(new_n957), .ZN(new_n967));
  INV_X1    g766(.A(new_n904), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n906), .A2(new_n907), .ZN(new_n969));
  INV_X1    g768(.A(new_n822), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n611), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(new_n973), .B2(new_n909), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n861), .B1(new_n974), .B2(new_n454), .ZN(new_n975));
  AOI211_X1 g774(.A(new_n669), .B(new_n967), .C1(new_n975), .C2(new_n915), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n966), .B1(new_n976), .B2(new_n964), .ZN(G1353gat));
  OAI211_X1 g776(.A(new_n611), .B(new_n957), .C1(new_n913), .C2(new_n916), .ZN(new_n978));
  NOR2_X1   g777(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n978), .A2(G211gat), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n954), .A2(new_n329), .A3(new_n611), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n967), .B1(new_n975), .B2(new_n915), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n329), .B1(new_n982), .B2(new_n611), .ZN(new_n983));
  XNOR2_X1  g782(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n980), .B(new_n981), .C1(new_n983), .C2(new_n984), .ZN(G1354gat));
  NAND3_X1  g784(.A1(new_n954), .A2(new_n330), .A3(new_n667), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n982), .A2(new_n667), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(new_n330), .ZN(G1355gat));
endmodule


