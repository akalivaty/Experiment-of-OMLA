

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XNOR2_X1 U323 ( .A(n345), .B(n344), .ZN(n555) );
  XOR2_X2 U324 ( .A(KEYINPUT124), .B(n474), .Z(n561) );
  XOR2_X1 U325 ( .A(G99GAT), .B(G85GAT), .Z(n330) );
  NOR2_X1 U326 ( .A1(n529), .A2(n424), .ZN(n426) );
  XNOR2_X1 U327 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U328 ( .A(KEYINPUT36), .B(n555), .Z(n579) );
  AND2_X1 U329 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  AND2_X1 U330 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U331 ( .A(KEYINPUT37), .B(n445), .Z(n293) );
  OR2_X1 U332 ( .A1(n517), .A2(n421), .ZN(n294) );
  XOR2_X1 U333 ( .A(KEYINPUT47), .B(n464), .Z(n295) );
  XNOR2_X1 U334 ( .A(n329), .B(n328), .ZN(n456) );
  INV_X1 U335 ( .A(KEYINPUT114), .ZN(n458) );
  XNOR2_X1 U336 ( .A(n458), .B(KEYINPUT46), .ZN(n459) );
  XNOR2_X1 U337 ( .A(n460), .B(n459), .ZN(n461) );
  OR2_X1 U338 ( .A1(n527), .A2(n531), .ZN(n424) );
  INV_X1 U339 ( .A(KEYINPUT96), .ZN(n425) );
  XNOR2_X1 U340 ( .A(n330), .B(n291), .ZN(n316) );
  XNOR2_X1 U341 ( .A(n316), .B(n432), .ZN(n320) );
  AND2_X1 U342 ( .A1(n294), .A2(n427), .ZN(n428) );
  XNOR2_X1 U343 ( .A(n403), .B(n402), .ZN(n404) );
  OR2_X1 U344 ( .A1(n528), .A2(n467), .ZN(n468) );
  XNOR2_X1 U345 ( .A(n335), .B(n292), .ZN(n336) );
  XNOR2_X1 U346 ( .A(n468), .B(KEYINPUT54), .ZN(n469) );
  XNOR2_X1 U347 ( .A(n337), .B(n336), .ZN(n341) );
  XNOR2_X1 U348 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U349 ( .A(n446), .B(KEYINPUT38), .ZN(n447) );
  XOR2_X1 U350 ( .A(KEYINPUT28), .B(n470), .Z(n531) );
  XNOR2_X1 U351 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n475) );
  XNOR2_X1 U352 ( .A(n449), .B(G50GAT), .ZN(n450) );
  XNOR2_X1 U353 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U354 ( .A(n476), .B(n475), .ZN(G1351GAT) );
  XNOR2_X1 U355 ( .A(n451), .B(n450), .ZN(G1331GAT) );
  XOR2_X1 U356 ( .A(G141GAT), .B(G197GAT), .Z(n297) );
  XNOR2_X1 U357 ( .A(G36GAT), .B(G50GAT), .ZN(n296) );
  XNOR2_X1 U358 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U359 ( .A(n298), .B(G15GAT), .Z(n300) );
  XOR2_X1 U360 ( .A(G113GAT), .B(G1GAT), .Z(n360) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(n360), .ZN(n299) );
  XNOR2_X1 U362 ( .A(n300), .B(n299), .ZN(n306) );
  XOR2_X1 U363 ( .A(G29GAT), .B(G43GAT), .Z(n302) );
  XNOR2_X1 U364 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n301) );
  XNOR2_X1 U365 ( .A(n302), .B(n301), .ZN(n343) );
  XOR2_X1 U366 ( .A(n343), .B(KEYINPUT68), .Z(n304) );
  NAND2_X1 U367 ( .A1(G229GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U369 ( .A(n306), .B(n305), .Z(n314) );
  XOR2_X1 U370 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n308) );
  XNOR2_X1 U371 ( .A(G22GAT), .B(G8GAT), .ZN(n307) );
  XNOR2_X1 U372 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U373 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n310) );
  XNOR2_X1 U374 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n309) );
  XNOR2_X1 U375 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U377 ( .A(n314), .B(n313), .ZN(n568) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(G57GAT), .ZN(n315) );
  XNOR2_X1 U379 ( .A(n315), .B(KEYINPUT13), .ZN(n432) );
  XOR2_X1 U380 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n318) );
  XNOR2_X1 U381 ( .A(KEYINPUT70), .B(KEYINPUT33), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U383 ( .A(n320), .B(n319), .Z(n329) );
  XNOR2_X1 U384 ( .A(G106GAT), .B(G78GAT), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n321), .B(G148GAT), .ZN(n377) );
  XOR2_X1 U386 ( .A(G64GAT), .B(G92GAT), .Z(n323) );
  XNOR2_X1 U387 ( .A(G176GAT), .B(G204GAT), .ZN(n322) );
  XNOR2_X1 U388 ( .A(n323), .B(n322), .ZN(n409) );
  XNOR2_X1 U389 ( .A(n377), .B(n409), .ZN(n327) );
  XOR2_X1 U390 ( .A(KEYINPUT73), .B(KEYINPUT71), .Z(n325) );
  XNOR2_X1 U391 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n324) );
  XOR2_X1 U392 ( .A(n325), .B(n324), .Z(n326) );
  NAND2_X1 U393 ( .A1(n568), .A2(n456), .ZN(n490) );
  XOR2_X1 U394 ( .A(KEYINPUT77), .B(n330), .Z(n332) );
  XOR2_X1 U395 ( .A(G36GAT), .B(G190GAT), .Z(n407) );
  XNOR2_X1 U396 ( .A(G218GAT), .B(n407), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U398 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n334) );
  XNOR2_X1 U399 ( .A(G92GAT), .B(KEYINPUT76), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U401 ( .A(KEYINPUT75), .B(KEYINPUT9), .Z(n339) );
  XNOR2_X1 U402 ( .A(G134GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U404 ( .A(n341), .B(n340), .Z(n345) );
  XNOR2_X1 U405 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n342), .B(G162GAT), .ZN(n378) );
  XNOR2_X1 U407 ( .A(n343), .B(n378), .ZN(n344) );
  XOR2_X1 U408 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n347) );
  NAND2_X1 U409 ( .A1(G225GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U411 ( .A(G57GAT), .B(n348), .ZN(n367) );
  XOR2_X1 U412 ( .A(G155GAT), .B(G148GAT), .Z(n350) );
  XNOR2_X1 U413 ( .A(G127GAT), .B(G162GAT), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U415 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n352) );
  XNOR2_X1 U416 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U418 ( .A(n354), .B(n353), .Z(n365) );
  XNOR2_X1 U419 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n355), .B(KEYINPUT83), .ZN(n356) );
  XOR2_X1 U421 ( .A(n356), .B(KEYINPUT0), .Z(n358) );
  XNOR2_X1 U422 ( .A(G120GAT), .B(G134GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n401) );
  XNOR2_X1 U424 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n359), .B(KEYINPUT2), .ZN(n368) );
  XOR2_X1 U426 ( .A(G85GAT), .B(n368), .Z(n362) );
  XNOR2_X1 U427 ( .A(G29GAT), .B(n360), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n401), .B(n363), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n517) );
  XOR2_X1 U432 ( .A(G22GAT), .B(G155GAT), .Z(n440) );
  XOR2_X1 U433 ( .A(n368), .B(n440), .Z(n370) );
  NAND2_X1 U434 ( .A1(G228GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n382) );
  XOR2_X1 U436 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n372) );
  XNOR2_X1 U437 ( .A(G204GAT), .B(KEYINPUT85), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U439 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n374) );
  XNOR2_X1 U440 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n373) );
  XNOR2_X1 U441 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U442 ( .A(n376), .B(n375), .Z(n380) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U446 ( .A(KEYINPUT21), .B(G218GAT), .Z(n384) );
  XNOR2_X1 U447 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U449 ( .A(G197GAT), .B(n385), .Z(n405) );
  XOR2_X1 U450 ( .A(n386), .B(n405), .Z(n470) );
  XOR2_X1 U451 ( .A(G15GAT), .B(G127GAT), .Z(n441) );
  XOR2_X1 U452 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n388) );
  XNOR2_X1 U453 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n403) );
  XOR2_X1 U455 ( .A(n441), .B(n403), .Z(n390) );
  XNOR2_X1 U456 ( .A(G190GAT), .B(G99GAT), .ZN(n389) );
  XNOR2_X1 U457 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U458 ( .A(G71GAT), .B(G176GAT), .Z(n392) );
  NAND2_X1 U459 ( .A1(G227GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U461 ( .A(n394), .B(n393), .Z(n399) );
  XOR2_X1 U462 ( .A(G183GAT), .B(KEYINPUT20), .Z(n396) );
  XNOR2_X1 U463 ( .A(G43GAT), .B(KEYINPUT84), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U465 ( .A(G113GAT), .B(n397), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n529) );
  XOR2_X1 U468 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n402) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U470 ( .A(n407), .B(n406), .Z(n413) );
  XNOR2_X1 U471 ( .A(G8GAT), .B(G183GAT), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n408), .B(G211GAT), .ZN(n433) );
  XNOR2_X1 U473 ( .A(n409), .B(n433), .ZN(n411) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n467) );
  INV_X1 U476 ( .A(n467), .ZN(n520) );
  NAND2_X1 U477 ( .A1(n529), .A2(n520), .ZN(n414) );
  NAND2_X1 U478 ( .A1(n470), .A2(n414), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n415), .B(KEYINPUT25), .ZN(n420) );
  NOR2_X1 U480 ( .A1(n529), .A2(n470), .ZN(n417) );
  XNOR2_X1 U481 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n416) );
  XOR2_X1 U482 ( .A(n417), .B(n416), .Z(n567) );
  XOR2_X1 U483 ( .A(n467), .B(KEYINPUT94), .Z(n418) );
  XNOR2_X1 U484 ( .A(n418), .B(KEYINPUT27), .ZN(n422) );
  AND2_X1 U485 ( .A1(n567), .A2(n422), .ZN(n419) );
  NOR2_X1 U486 ( .A1(n420), .A2(n419), .ZN(n421) );
  NAND2_X1 U487 ( .A1(n422), .A2(n517), .ZN(n423) );
  XOR2_X1 U488 ( .A(n423), .B(KEYINPUT95), .Z(n527) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U490 ( .A(KEYINPUT98), .B(n428), .ZN(n488) );
  NOR2_X1 U491 ( .A1(n579), .A2(n488), .ZN(n444) );
  XOR2_X1 U492 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n430) );
  NAND2_X1 U493 ( .A1(G231GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U495 ( .A(n431), .B(KEYINPUT14), .Z(n435) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U498 ( .A(KEYINPUT15), .B(G64GAT), .Z(n437) );
  XNOR2_X1 U499 ( .A(G1GAT), .B(G78GAT), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U501 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n576) );
  NAND2_X1 U504 ( .A1(n444), .A2(n576), .ZN(n445) );
  NOR2_X1 U505 ( .A1(n490), .A2(n293), .ZN(n448) );
  INV_X1 U506 ( .A(KEYINPUT105), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n503) );
  NAND2_X1 U508 ( .A1(n503), .A2(n531), .ZN(n451) );
  XOR2_X1 U509 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n449) );
  INV_X1 U510 ( .A(n456), .ZN(n571) );
  NOR2_X1 U511 ( .A1(n579), .A2(n576), .ZN(n452) );
  XOR2_X1 U512 ( .A(KEYINPUT45), .B(n452), .Z(n453) );
  NOR2_X1 U513 ( .A1(n571), .A2(n453), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT116), .B(n454), .Z(n455) );
  NOR2_X1 U515 ( .A1(n568), .A2(n455), .ZN(n465) );
  XNOR2_X1 U516 ( .A(n576), .B(KEYINPUT113), .ZN(n560) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT64), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(KEYINPUT41), .ZN(n546) );
  NAND2_X1 U519 ( .A1(n568), .A2(n546), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n560), .A2(n461), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT115), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n463), .A2(n555), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n465), .A2(n295), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT48), .ZN(n528) );
  NOR2_X1 U525 ( .A1(n517), .A2(n469), .ZN(n566) );
  NAND2_X1 U526 ( .A1(n566), .A2(n470), .ZN(n472) );
  XOR2_X1 U527 ( .A(KEYINPUT123), .B(KEYINPUT55), .Z(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n473), .A2(n529), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n561), .A2(n555), .ZN(n476) );
  NAND2_X1 U531 ( .A1(n517), .A2(n503), .ZN(n480) );
  XOR2_X1 U532 ( .A(G29GAT), .B(KEYINPUT104), .Z(n478) );
  XNOR2_X1 U533 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n480), .B(n479), .ZN(G1328GAT) );
  NAND2_X1 U535 ( .A1(n546), .A2(n561), .ZN(n483) );
  XOR2_X1 U536 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(G176GAT), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  XNOR2_X1 U539 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n485) );
  NOR2_X1 U540 ( .A1(n555), .A2(n576), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U542 ( .A(n486), .B(KEYINPUT79), .ZN(n487) );
  NOR2_X1 U543 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U544 ( .A(KEYINPUT99), .B(n489), .ZN(n506) );
  NOR2_X1 U545 ( .A1(n490), .A2(n506), .ZN(n491) );
  XNOR2_X1 U546 ( .A(n491), .B(KEYINPUT100), .ZN(n499) );
  NAND2_X1 U547 ( .A1(n517), .A2(n499), .ZN(n492) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(n492), .ZN(n493) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  XOR2_X1 U550 ( .A(G8GAT), .B(KEYINPUT101), .Z(n495) );
  NAND2_X1 U551 ( .A1(n499), .A2(n520), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n495), .B(n494), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n497) );
  NAND2_X1 U554 ( .A1(n499), .A2(n529), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n498), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT103), .Z(n501) );
  NAND2_X1 U558 ( .A1(n499), .A2(n531), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(G1327GAT) );
  NAND2_X1 U560 ( .A1(n503), .A2(n520), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n503), .A2(n529), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(KEYINPUT40), .ZN(n505) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  INV_X1 U566 ( .A(n568), .ZN(n542) );
  NAND2_X1 U567 ( .A1(n546), .A2(n542), .ZN(n515) );
  NOR2_X1 U568 ( .A1(n506), .A2(n515), .ZN(n512) );
  NAND2_X1 U569 ( .A1(n517), .A2(n512), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  XOR2_X1 U571 ( .A(G64GAT), .B(KEYINPUT109), .Z(n510) );
  NAND2_X1 U572 ( .A1(n512), .A2(n520), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n529), .A2(n512), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U577 ( .A1(n512), .A2(n531), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  XOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT111), .Z(n519) );
  NOR2_X1 U580 ( .A1(n515), .A2(n293), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT110), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n517), .A2(n524), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n524), .A2(n520), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(KEYINPUT112), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n524), .A2(n529), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n531), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT117), .Z(n533) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n541), .A2(n529), .ZN(n530) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n538), .A2(n568), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U599 ( .A1(n538), .A2(n546), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n560), .A2(n538), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n555), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n541), .A2(n567), .ZN(n556) );
  NOR2_X1 U608 ( .A1(n542), .A2(n556), .ZN(n543) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n551) );
  INV_X1 U613 ( .A(n546), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n547), .A2(n556), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n576), .A2(n556), .ZN(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  INV_X1 U622 ( .A(n555), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n568), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT125), .Z(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT126), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(n565), .Z(n570) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n578) );
  INV_X1 U634 ( .A(n578), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n572), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  OR2_X1 U641 ( .A1(n578), .A2(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

