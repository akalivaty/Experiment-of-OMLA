//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n212), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n210), .B(new_n224), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT9), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n225), .B1(new_n206), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n253), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n265), .B(new_n225), .C1(new_n251), .C2(new_n206), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n202), .B1(new_n264), .B2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n265), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n267), .A2(new_n268), .B1(new_n202), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n250), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n262), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n257), .B2(new_n259), .ZN(new_n274));
  OAI211_X1 g0074(.A(KEYINPUT9), .B(new_n270), .C1(new_n274), .C2(new_n253), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT10), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n272), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n276), .A2(KEYINPUT10), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n284), .A3(G274), .ZN(new_n285));
  INV_X1    g0085(.A(G226), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n281), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G222), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G223), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n291), .B1(new_n218), .B2(new_n289), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(G190), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n278), .A2(new_n280), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n297), .B2(new_n296), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n272), .A2(new_n275), .A3(new_n277), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n279), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n270), .B1(new_n274), .B2(new_n253), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n305), .B(new_n306), .C1(G169), .C2(new_n296), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n300), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n285), .B1(new_n219), .B2(new_n287), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n289), .A2(G232), .A3(new_n290), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G107), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n310), .B(new_n315), .C1(new_n292), .C2(new_n213), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n309), .B1(new_n316), .B2(new_n295), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n304), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n264), .A2(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G77), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n266), .A2(new_n320), .B1(G77), .B2(new_n265), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G20), .A2(G77), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n254), .A2(new_n251), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(new_n258), .B2(new_n323), .C1(new_n255), .C2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n325), .B2(new_n252), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n318), .B(new_n327), .C1(G169), .C2(new_n317), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n316), .A2(new_n295), .ZN(new_n329));
  INV_X1    g0129(.A(new_n309), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(G190), .A3(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n331), .B(new_n326), .C1(new_n297), .C2(new_n317), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n289), .A2(G232), .A3(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n289), .A2(G226), .A3(new_n290), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n295), .ZN(new_n338));
  INV_X1    g0138(.A(G274), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n295), .A2(new_n339), .A3(new_n281), .ZN(new_n340));
  INV_X1    g0140(.A(new_n287), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(G238), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT13), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n338), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT69), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n212), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n255), .B(KEYINPUT67), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n218), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n212), .B1(new_n264), .B2(G20), .ZN(new_n354));
  OR3_X1    g0154(.A1(new_n265), .A2(KEYINPUT12), .A3(G68), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT12), .B1(new_n265), .B2(G68), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n267), .A2(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT11), .B1(new_n352), .B2(new_n252), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n349), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n359), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n361), .A2(KEYINPUT69), .A3(new_n353), .A4(new_n357), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n348), .A2(G190), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n347), .A2(G200), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n333), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n308), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(new_n362), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  INV_X1    g0168(.A(new_n346), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n345), .B1(new_n338), .B2(new_n342), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(G169), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT70), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n344), .B2(new_n346), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT70), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n368), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n374), .A2(new_n368), .B1(new_n347), .B2(new_n304), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n367), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n366), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n289), .A2(G226), .A3(G1698), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n311), .A2(new_n313), .A3(G223), .A4(new_n290), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G87), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n295), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n339), .B1(new_n226), .B2(new_n283), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n341), .A2(G232), .B1(new_n388), .B2(new_n282), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n387), .A2(G190), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n297), .B1(new_n387), .B2(new_n389), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n289), .A2(new_n393), .A3(G20), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n314), .B2(new_n254), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n398), .B2(new_n201), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n261), .A2(G159), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n254), .B1(new_n230), .B2(new_n397), .ZN(new_n403));
  INV_X1    g0203(.A(G159), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n323), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT71), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n402), .A4(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n393), .B1(new_n289), .B2(G20), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n314), .A2(KEYINPUT7), .A3(new_n254), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n212), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n399), .A2(new_n401), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n413), .A3(new_n252), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n259), .A2(new_n319), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n415), .A2(new_n266), .B1(new_n265), .B2(new_n259), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n392), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n406), .A2(new_n402), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n411), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n253), .B1(new_n422), .B2(KEYINPUT16), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n416), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(KEYINPUT17), .A3(new_n392), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT72), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n420), .A2(new_n425), .A3(KEYINPUT72), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n414), .A2(new_n417), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n387), .A2(new_n389), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G169), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n304), .B2(new_n432), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n434), .A3(KEYINPUT18), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n381), .A2(new_n382), .A3(new_n430), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n377), .A2(new_n379), .ZN(new_n441));
  INV_X1    g0241(.A(new_n367), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n308), .A3(new_n365), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n428), .A2(new_n429), .A3(new_n439), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT73), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT77), .B1(new_n448), .B2(G41), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  INV_X1    g0250(.A(G41), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(KEYINPUT76), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n450), .B(new_n451), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n264), .B(G45), .C1(new_n451), .C2(KEYINPUT5), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n449), .A2(new_n388), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n457), .B1(new_n462), .B2(KEYINPUT77), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(KEYINPUT78), .A3(new_n388), .A4(new_n456), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n454), .A2(KEYINPUT76), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n467));
  AOI21_X1  g0267(.A(G41), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n458), .B1(new_n468), .B2(new_n450), .ZN(new_n469));
  INV_X1    g0269(.A(new_n456), .ZN(new_n470));
  OAI211_X1 g0270(.A(G270), .B(new_n284), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n289), .A2(G257), .A3(new_n290), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n314), .A2(G303), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(new_n292), .C2(new_n221), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n295), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(G200), .B1(new_n465), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n265), .A2(G116), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n264), .A2(KEYINPUT74), .A3(G33), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT74), .B1(new_n264), .B2(G33), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n266), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n481), .B2(G116), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n254), .C1(G33), .C2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G20), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n252), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n471), .A2(new_n475), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n461), .A2(new_n464), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(G190), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n477), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n373), .B1(new_n482), .B2(new_n490), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n465), .B2(new_n476), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT79), .A2(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n499), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n497), .C1(new_n465), .C2(new_n476), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n493), .A2(new_n491), .A3(G179), .A4(new_n494), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n496), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n311), .A2(new_n313), .A3(G244), .A4(new_n290), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(KEYINPUT75), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(KEYINPUT75), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n289), .A2(G244), .A3(new_n290), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n508), .A2(new_n483), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n295), .ZN(new_n513));
  OAI211_X1 g0313(.A(G257), .B(new_n284), .C1(new_n469), .C2(new_n470), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n494), .A2(new_n304), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n484), .A2(new_n220), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G97), .A2(G107), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n220), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n522));
  OAI21_X1  g0322(.A(G107), .B1(new_n394), .B2(new_n395), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n253), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n269), .A2(new_n484), .ZN(new_n525));
  INV_X1    g0325(.A(new_n481), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(new_n484), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n513), .A2(new_n514), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n465), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n515), .B(new_n528), .C1(new_n530), .C2(G169), .ZN(new_n531));
  OAI21_X1  g0331(.A(G200), .B1(new_n465), .B2(new_n529), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n524), .A2(new_n527), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n494), .A2(G190), .A3(new_n513), .A4(new_n514), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT25), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n265), .B2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n220), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n481), .A2(G107), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n311), .A2(new_n313), .A3(new_n254), .A4(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT22), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n289), .A2(new_n544), .A3(new_n254), .A4(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G20), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT23), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n254), .B2(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n220), .A2(KEYINPUT23), .A3(G20), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT24), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n546), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n541), .B1(new_n557), .B2(new_n252), .ZN(new_n558));
  OAI211_X1 g0358(.A(G264), .B(new_n284), .C1(new_n469), .C2(new_n470), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n289), .A2(G257), .A3(G1698), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n289), .A2(G250), .A3(new_n290), .ZN(new_n561));
  INV_X1    g0361(.A(G294), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(new_n561), .C1(new_n251), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n295), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(G200), .B1(new_n465), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n494), .A2(G190), .A3(new_n559), .A4(new_n564), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n558), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n556), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n555), .B1(new_n546), .B2(new_n552), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n252), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n540), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n373), .B1(new_n465), .B2(new_n565), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n494), .A2(new_n304), .A3(new_n559), .A4(new_n564), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G45), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n215), .B1(new_n576), .B2(G1), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n264), .A2(new_n339), .A3(G45), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n284), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n311), .A2(new_n313), .A3(G238), .A4(new_n290), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n311), .A2(new_n313), .A3(G244), .A4(G1698), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n547), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n580), .B1(new_n583), .B2(new_n295), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n297), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(G190), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n254), .B1(new_n336), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n518), .A2(new_n214), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n311), .A2(new_n313), .A3(new_n254), .A4(G68), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n588), .B1(new_n255), .B2(new_n484), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n252), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n479), .A2(new_n480), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n267), .A2(G87), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n324), .A2(new_n269), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n586), .A2(new_n587), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n324), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n267), .A2(new_n602), .A3(new_n596), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n595), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n584), .A2(G169), .ZN(new_n605));
  AOI211_X1 g0405(.A(G179), .B(new_n580), .C1(new_n583), .C2(new_n295), .ZN(new_n606));
  OR3_X1    g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n568), .A2(new_n575), .A3(new_n601), .A4(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n447), .A2(new_n505), .A3(new_n536), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT80), .ZN(G372));
  INV_X1    g0410(.A(KEYINPUT26), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT81), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n585), .B2(new_n599), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n587), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n594), .A2(new_n252), .B1(new_n269), .B2(new_n324), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n597), .C1(new_n584), .C2(new_n297), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n612), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n607), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n611), .B1(new_n618), .B2(new_n531), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT83), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n621), .B(new_n611), .C1(new_n618), .C2(new_n531), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n607), .A2(new_n601), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n531), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(KEYINPUT82), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n616), .A2(new_n612), .B1(G190), .B2(new_n584), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n586), .A2(KEYINPUT81), .A3(new_n600), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n531), .A2(new_n631), .A3(new_n568), .A4(new_n535), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n575), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n447), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT84), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n431), .A2(KEYINPUT18), .A3(new_n434), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT18), .B1(new_n431), .B2(new_n434), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n437), .A2(KEYINPUT84), .A3(new_n438), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n363), .A2(new_n364), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n443), .B1(new_n643), .B2(new_n328), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n642), .B1(new_n644), .B2(new_n430), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n300), .A2(new_n303), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n307), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n636), .A2(new_n647), .ZN(G369));
  NAND3_X1  g0448(.A1(new_n264), .A2(new_n254), .A3(G13), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n649), .A2(KEYINPUT85), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(KEYINPUT85), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n655), .A3(G213), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n492), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n502), .A2(new_n503), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n493), .A2(new_n494), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n501), .B1(new_n662), .B2(new_n497), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n660), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n504), .B2(new_n660), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n659), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n572), .A2(new_n658), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n568), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n669), .B2(new_n575), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n659), .B1(new_n661), .B2(new_n663), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT86), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT86), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n676), .B(new_n659), .C1(new_n661), .C2(new_n663), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n667), .B1(new_n678), .B2(new_n670), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(G399));
  NOR2_X1   g0480(.A1(new_n590), .A2(G116), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n207), .A2(new_n451), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n231), .B2(new_n682), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n465), .B1(new_n529), .B2(new_n565), .ZN(new_n686));
  INV_X1    g0486(.A(new_n584), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n304), .B(new_n687), .C1(new_n465), .C2(new_n476), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n494), .A2(G179), .A3(new_n475), .A4(new_n471), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT87), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n493), .A2(KEYINPUT87), .A3(G179), .A4(new_n494), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n565), .A2(new_n687), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n692), .A2(new_n530), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n689), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n494), .A2(new_n513), .A3(new_n514), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n698), .A2(new_n565), .A3(new_n687), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n692), .A3(KEYINPUT30), .A4(new_n693), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n659), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n608), .A2(new_n505), .A3(new_n536), .A4(new_n659), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(KEYINPUT31), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n701), .A2(KEYINPUT31), .ZN(new_n704));
  OAI21_X1  g0504(.A(G330), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n632), .A2(new_n633), .ZN(new_n706));
  INV_X1    g0506(.A(new_n628), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n624), .A2(new_n611), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT26), .B1(new_n618), .B2(new_n531), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n659), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n635), .A2(new_n714), .A3(new_n659), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n705), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n685), .B1(new_n716), .B2(G1), .ZN(G364));
  INV_X1    g0517(.A(G13), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n264), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n682), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n289), .A2(new_n207), .ZN(new_n724));
  INV_X1    g0524(.A(G355), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n724), .A2(new_n725), .B1(G116), .B2(new_n207), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n248), .A2(new_n576), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n314), .A2(new_n207), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n576), .B2(new_n232), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n225), .B1(G20), .B2(new_n373), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n723), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G190), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n254), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n304), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n254), .A2(G190), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G322), .A2(new_n742), .B1(new_n746), .B2(G329), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n254), .B1(new_n744), .B2(G190), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n562), .B2(new_n748), .ZN(new_n749));
  OR3_X1    g0549(.A1(new_n297), .A2(KEYINPUT90), .A3(G179), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT90), .B1(new_n297), .B2(G179), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(new_n743), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n749), .B1(G283), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n254), .A2(new_n304), .A3(new_n297), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT89), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT89), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(G190), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n738), .A3(new_n757), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G326), .A2(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT88), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n740), .A2(new_n743), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(new_n740), .B2(new_n743), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n754), .B(new_n763), .C1(new_n764), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n750), .A2(new_n739), .A3(new_n751), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n314), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT91), .Z(new_n775));
  NOR2_X1   g0575(.A1(new_n745), .A2(new_n404), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n777), .B1(new_n220), .B2(new_n752), .C1(new_n770), .C2(new_n218), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n772), .A2(new_n214), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n748), .A2(new_n484), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n289), .B1(new_n741), .B2(new_n229), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n782), .B1(new_n202), .B2(new_n758), .C1(new_n212), .C2(new_n760), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n771), .A2(new_n775), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n737), .B1(new_n784), .B2(new_n734), .ZN(new_n785));
  INV_X1    g0585(.A(new_n733), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n665), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT92), .Z(new_n788));
  INV_X1    g0588(.A(new_n666), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n723), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G330), .B2(new_n665), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(new_n791), .ZN(G396));
  INV_X1    g0592(.A(KEYINPUT96), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n658), .A2(new_n327), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n332), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n328), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n329), .A2(new_n330), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n326), .B1(new_n797), .B2(new_n373), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(new_n318), .A3(new_n659), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n793), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n332), .A2(new_n794), .B1(new_n798), .B2(new_n318), .ZN(new_n801));
  AND3_X1   g0601(.A1(new_n798), .A2(new_n318), .A3(new_n659), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n801), .A2(new_n802), .A3(KEYINPUT96), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n659), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(KEYINPUT97), .B1(new_n635), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT97), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n807), .B(new_n804), .C1(new_n626), .C2(new_n634), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n800), .A2(new_n803), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n635), .B2(new_n659), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n705), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n705), .B1(new_n809), .B2(new_n812), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n722), .C2(new_n721), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n734), .A2(new_n731), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n723), .B1(G77), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n769), .A2(G159), .B1(G143), .B2(new_n742), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n758), .C1(new_n822), .C2(new_n760), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT95), .Z(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n752), .A2(new_n212), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n289), .B1(new_n748), .B2(new_n229), .C1(new_n827), .C2(new_n745), .ZN(new_n828));
  INV_X1    g0628(.A(new_n772), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n826), .B(new_n828), .C1(G50), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n759), .A2(G303), .B1(G116), .B2(new_n769), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT93), .B(G283), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n760), .B2(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT94), .Z(new_n836));
  OAI221_X1 g0636(.A(new_n314), .B1(new_n745), .B2(new_n764), .C1(new_n741), .C2(new_n562), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n780), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n753), .A2(G87), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n838), .B(new_n839), .C1(new_n220), .C2(new_n772), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n831), .A2(new_n832), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n819), .B1(new_n841), .B2(new_n734), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n732), .B2(new_n811), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n817), .A2(new_n843), .ZN(G384));
  NAND2_X1  g0644(.A1(new_n397), .A2(G77), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n231), .A2(new_n845), .B1(G50), .B2(new_n212), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(G1), .A3(new_n718), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT98), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(G116), .A3(new_n228), .A4(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT36), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n423), .B1(KEYINPUT16), .B2(new_n422), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n417), .ZN(new_n856));
  INV_X1    g0656(.A(new_n656), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n445), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n434), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(new_n858), .A3(new_n418), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n656), .B1(new_n414), .B2(new_n417), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n424), .B2(new_n392), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT37), .B1(new_n431), .B2(new_n434), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n865), .A2(KEYINPUT100), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT100), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n860), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT38), .B1(new_n860), .B2(new_n869), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n799), .B1(new_n806), .B2(new_n808), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT99), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n380), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n378), .B1(new_n376), .B2(new_n372), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT99), .B1(new_n876), .B2(new_n367), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n367), .A2(new_n659), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n643), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n441), .A2(new_n878), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n872), .A2(new_n873), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n642), .A2(new_n656), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n870), .A2(new_n871), .A3(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n640), .A2(new_n641), .A3(new_n420), .A4(new_n425), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n864), .ZN(new_n890));
  INV_X1    g0690(.A(new_n864), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n418), .C1(new_n435), .C2(new_n637), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT84), .B1(new_n431), .B2(new_n434), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n867), .B2(new_n868), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n860), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT39), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n888), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n875), .A2(new_n877), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n658), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT101), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n883), .A2(new_n905), .A3(new_n884), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n886), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT103), .ZN(new_n908));
  INV_X1    g0708(.A(new_n711), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n658), .B1(new_n909), .B2(new_n634), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n714), .ZN(new_n911));
  AOI211_X1 g0711(.A(KEYINPUT29), .B(new_n658), .C1(new_n626), .C2(new_n634), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n447), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT102), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT102), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n447), .B(new_n915), .C1(new_n911), .C2(new_n912), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n647), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n908), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT40), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n870), .A2(new_n871), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n882), .B(new_n811), .C1(new_n703), .C2(new_n704), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n898), .A2(new_n899), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n703), .A2(new_n704), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n810), .B1(new_n880), .B2(new_n881), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT40), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n440), .A2(new_n446), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n929), .B2(new_n924), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n922), .A2(new_n447), .A3(new_n925), .A4(new_n927), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(G330), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n918), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n264), .B2(new_n719), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n918), .A2(new_n932), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n854), .B1(new_n934), .B2(new_n935), .ZN(G367));
  OAI221_X1 g0736(.A(new_n735), .B1(new_n207), .B2(new_n324), .C1(new_n240), .C2(new_n728), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n723), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n752), .A2(new_n484), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n289), .B(new_n939), .C1(G317), .C2(new_n746), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT112), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n741), .A2(new_n773), .B1(new_n748), .B2(new_n220), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n770), .A2(new_n834), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(G311), .C2(new_n759), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT46), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n829), .A2(G116), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n946), .A2(new_n947), .B1(new_n760), .B2(new_n562), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n941), .A2(KEYINPUT112), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n942), .A2(new_n945), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n770), .A2(new_n202), .B1(new_n404), .B2(new_n760), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT113), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n759), .A2(G143), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n748), .A2(new_n212), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n289), .B1(new_n741), .B2(new_n822), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G137), .B2(new_n746), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G58), .A2(new_n829), .B1(new_n753), .B2(G77), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n954), .A2(new_n955), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n951), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT47), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n938), .B1(new_n961), .B2(new_n734), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n659), .A2(new_n600), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n628), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n618), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n962), .B1(new_n786), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT111), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n678), .A2(new_n670), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n677), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n676), .B1(new_n971), .B2(new_n659), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n670), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n973), .A2(KEYINPUT110), .A3(new_n666), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n666), .B1(new_n973), .B2(KEYINPUT110), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(KEYINPUT110), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n789), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n973), .A2(KEYINPUT110), .A3(new_n666), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n968), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n705), .A2(new_n713), .A3(new_n715), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n967), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT109), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n528), .A2(new_n658), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n531), .A2(new_n535), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n533), .B1(new_n698), .B2(new_n373), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(new_n515), .A3(new_n658), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n985), .B1(new_n679), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n667), .ZN(new_n992));
  AND4_X1   g0792(.A1(new_n985), .A2(new_n973), .A3(new_n992), .A4(new_n990), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n984), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n973), .A2(new_n992), .ZN(new_n995));
  INV_X1    g0795(.A(new_n990), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT109), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n679), .A2(new_n985), .A3(new_n990), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT45), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(KEYINPUT44), .A3(new_n996), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n679), .B2(new_n990), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n994), .A2(new_n999), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n672), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n994), .A2(new_n999), .A3(new_n673), .A4(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n976), .A2(new_n980), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n716), .A2(KEYINPUT111), .A3(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n983), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n716), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n682), .B(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n721), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n987), .A2(KEYINPUT104), .A3(new_n989), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT104), .B1(new_n987), .B2(new_n989), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n673), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT105), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n531), .C1(new_n1018), .C2(new_n575), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT104), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n990), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n575), .B1(new_n1023), .B2(new_n1015), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n531), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT105), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1021), .A2(new_n1026), .A3(new_n659), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n1028));
  OR2_X1    g0828(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n973), .A2(new_n996), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n678), .A2(new_n670), .A3(new_n990), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1030), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1027), .A2(new_n1028), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT107), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n965), .B(KEYINPUT43), .Z(new_n1037));
  AOI22_X1  g0837(.A1(new_n1034), .A2(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1027), .A2(new_n1033), .A3(KEYINPUT107), .A4(new_n1028), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1019), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1042));
  AND4_X1   g0842(.A1(new_n1019), .A2(new_n1041), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n966), .B1(new_n1014), .B2(new_n1044), .ZN(G387));
  OAI22_X1  g0845(.A1(new_n724), .A2(new_n681), .B1(G107), .B2(new_n207), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n237), .A2(new_n576), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n681), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n1048), .C1(G68), .C2(G77), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n258), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n728), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1046), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n723), .B1(new_n1053), .B2(new_n736), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT114), .Z(new_n1055));
  NOR2_X1   g0855(.A1(new_n748), .A2(new_n324), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n289), .B1(new_n745), .B2(new_n822), .C1(new_n741), .C2(new_n202), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n759), .C2(G159), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n772), .A2(new_n218), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n939), .B(new_n1059), .C1(G68), .C2(new_n769), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n258), .C2(new_n760), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT115), .Z(new_n1062));
  AOI21_X1  g0862(.A(new_n289), .B1(new_n746), .B2(G326), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n772), .A2(new_n562), .B1(new_n748), .B2(new_n834), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n759), .A2(G322), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n769), .A2(G303), .B1(G317), .B2(new_n742), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n764), .C2(new_n760), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1063), .B1(new_n486), .B2(new_n752), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1062), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1055), .B1(new_n734), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n670), .B2(new_n786), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n722), .B1(new_n981), .B2(new_n982), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n716), .A2(new_n1007), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1076), .B1(new_n720), .B2(new_n981), .C1(new_n1077), .C2(new_n1078), .ZN(G393));
  AND2_X1   g0879(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n981), .A2(new_n982), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1009), .B(new_n722), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1018), .A2(new_n733), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n735), .B1(new_n484), .B2(new_n207), .C1(new_n244), .C2(new_n728), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n723), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n759), .A2(G317), .B1(G311), .B2(new_n742), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT117), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT52), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n289), .B1(new_n746), .B2(G322), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n486), .B2(new_n748), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n770), .A2(new_n562), .B1(new_n772), .B2(new_n834), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(G107), .C2(new_n753), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1088), .B(new_n1092), .C1(new_n773), .C2(new_n760), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1087), .A2(KEYINPUT52), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n758), .A2(new_n822), .B1(new_n741), .B2(new_n404), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n769), .A2(new_n259), .B1(G68), .B2(new_n829), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n748), .A2(new_n218), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n314), .B(new_n1099), .C1(G143), .C2(new_n746), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1098), .A2(new_n839), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n202), .C2(new_n760), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1093), .A2(new_n1094), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1085), .B1(new_n1104), .B2(new_n734), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1080), .A2(new_n721), .B1(new_n1083), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1082), .A2(new_n1106), .ZN(G390));
  INV_X1    g0907(.A(new_n882), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n802), .B1(new_n910), .B2(new_n811), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n923), .B1(new_n658), .B2(new_n902), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n903), .B1(new_n873), .B2(new_n882), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n901), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n705), .A2(new_n1108), .A3(new_n810), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n814), .A2(new_n811), .A3(new_n882), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1115), .B(new_n1110), .C1(new_n1111), .C2(new_n901), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n929), .A2(new_n705), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n647), .B(new_n1118), .C1(new_n914), .C2(new_n916), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1108), .B1(new_n705), .B2(new_n810), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n873), .B1(new_n1121), .B2(new_n1113), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1115), .A2(new_n1109), .A3(new_n1120), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1114), .A2(new_n1116), .A3(new_n1119), .A4(new_n1124), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n722), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1114), .A2(new_n721), .A3(new_n1116), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n723), .B1(new_n259), .B2(new_n818), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n314), .B1(new_n745), .B2(new_n562), .C1(new_n741), .C2(new_n486), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1099), .B(new_n1131), .C1(new_n759), .C2(G283), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n826), .B(new_n779), .C1(G97), .C2(new_n769), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n220), .C2(new_n760), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n752), .A2(new_n202), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n314), .B1(new_n746), .B2(G125), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n404), .B2(new_n748), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT54), .B(G143), .Z(new_n1138));
  AOI211_X1 g0938(.A(new_n1135), .B(new_n1137), .C1(new_n769), .C2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n772), .A2(new_n822), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT53), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n821), .C2(new_n760), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n758), .A2(new_n1143), .B1(new_n741), .B2(new_n827), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT118), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1134), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1130), .B1(new_n1146), .B2(new_n734), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n901), .B2(new_n732), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1128), .A2(new_n1129), .A3(new_n1148), .ZN(G378));
  NAND3_X1  g0949(.A1(new_n922), .A2(G330), .A3(new_n927), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n306), .A2(new_n857), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT120), .Z(new_n1152));
  XOR2_X1   g0952(.A(new_n308), .B(new_n1152), .Z(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n922), .A2(G330), .A3(new_n927), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n907), .A2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n885), .A2(KEYINPUT101), .B1(new_n903), .B2(new_n901), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1161), .A2(new_n906), .A3(new_n1158), .A4(new_n1156), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1162), .A3(new_n721), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n723), .B1(G50), .B2(new_n818), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G125), .A2(new_n759), .B1(new_n761), .B2(G132), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n741), .A2(new_n1143), .B1(new_n748), .B2(new_n822), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n829), .B2(new_n1138), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(new_n821), .C2(new_n770), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n753), .A2(G159), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n746), .C2(G124), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n955), .B1(new_n758), .B2(new_n486), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT119), .Z(new_n1175));
  OAI22_X1  g0975(.A1(new_n770), .A2(new_n324), .B1(new_n229), .B2(new_n752), .ZN(new_n1176));
  INV_X1    g0976(.A(G283), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n745), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n289), .A2(G41), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n220), .B2(new_n741), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1176), .A2(new_n1059), .A3(new_n1178), .A4(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1175), .B(new_n1181), .C1(new_n484), .C2(new_n760), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT58), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1173), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1185), .B1(new_n1183), .B2(new_n1182), .C1(new_n1179), .C2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1164), .B1(new_n1187), .B2(new_n734), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1155), .B2(new_n732), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT121), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1163), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1127), .A2(new_n1119), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1193), .A2(KEYINPUT57), .A3(new_n1162), .A4(new_n1160), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n722), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n907), .A2(new_n1159), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1161), .A2(new_n906), .B1(new_n1158), .B2(new_n1156), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1193), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1192), .B1(new_n1195), .B2(new_n1199), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n1108), .A2(new_n731), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n723), .B1(G68), .B2(new_n818), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT122), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n761), .A2(G116), .B1(G107), .B2(new_n769), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT123), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n218), .A2(new_n752), .B1(new_n772), .B2(new_n484), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n314), .B1(new_n745), .B2(new_n773), .C1(new_n741), .C2(new_n1177), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n1056), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1204), .A2(KEYINPUT123), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n759), .A2(G294), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n772), .A2(new_n404), .B1(new_n1143), .B2(new_n745), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT124), .Z(new_n1213));
  NOR2_X1   g1013(.A1(new_n752), .A2(new_n229), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n289), .B1(new_n748), .B2(new_n202), .C1(new_n741), .C2(new_n821), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(G150), .C2(new_n769), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G132), .A2(new_n759), .B1(new_n761), .B2(new_n1138), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1213), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1211), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1203), .B1(new_n1219), .B2(new_n734), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1124), .A2(new_n721), .B1(new_n1201), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1125), .A2(new_n1013), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(G381));
  OR2_X1    g1024(.A1(G375), .A2(G378), .ZN(new_n1225));
  OR2_X1    g1025(.A1(G393), .A2(G396), .ZN(new_n1226));
  OR4_X1    g1026(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1226), .ZN(new_n1227));
  OR3_X1    g1027(.A1(new_n1225), .A2(G387), .A3(new_n1227), .ZN(G407));
  OAI211_X1 g1028(.A(G407), .B(G213), .C1(G343), .C2(new_n1225), .ZN(G409));
  INV_X1    g1029(.A(KEYINPUT61), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n917), .B1(new_n929), .B2(new_n705), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1231), .A2(KEYINPUT60), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1232), .A2(new_n722), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1221), .ZN(new_n1237));
  INV_X1    g1037(.A(G384), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(G384), .A3(new_n1221), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n657), .A2(G213), .A3(G2897), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1241), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G384), .B1(new_n1236), .B2(new_n1221), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1221), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1245), .B(new_n1238), .C1(new_n1233), .C2(new_n1235), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1243), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1242), .A2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G378), .B(new_n1192), .C1(new_n1195), .C2(new_n1199), .ZN(new_n1249));
  INV_X1    g1049(.A(G378), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1198), .A2(new_n1013), .A3(new_n1193), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n1191), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1249), .A2(new_n1252), .B1(G213), .B2(new_n657), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1230), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n657), .A2(G213), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1256), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G390), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G387), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT125), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1012), .B1(new_n1009), .B2(new_n716), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n721), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(new_n966), .A3(G390), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1264), .A2(new_n1265), .A3(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(G393), .B(G396), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G390), .B1(new_n1268), .B2(new_n966), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(KEYINPUT125), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1264), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1255), .A2(new_n1262), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1259), .A2(KEYINPUT62), .A3(new_n1261), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1253), .B2(new_n1260), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1282), .A2(new_n1254), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1281), .B1(new_n1285), .B2(new_n1279), .ZN(G405));
  NAND2_X1  g1086(.A1(G375), .A2(new_n1250), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT127), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1249), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1279), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1249), .A2(new_n1288), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1291), .A2(new_n1278), .A3(new_n1274), .A4(new_n1277), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1290), .A2(new_n1261), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1261), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1287), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1279), .A2(new_n1289), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1270), .A2(new_n1273), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1291), .B1(new_n1297), .B2(new_n1278), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1260), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1287), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1290), .A2(new_n1292), .A3(new_n1261), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1302), .ZN(G402));
endmodule


