

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U321 ( .A(KEYINPUT41), .B(n572), .ZN(n558) );
  XNOR2_X1 U322 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n428) );
  XNOR2_X1 U323 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U324 ( .A(n429), .B(n428), .ZN(n449) );
  XNOR2_X1 U325 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U326 ( .A(n380), .B(n379), .ZN(n572) );
  NOR2_X1 U327 ( .A1(n460), .A2(n445), .ZN(n561) );
  XOR2_X1 U328 ( .A(n468), .B(KEYINPUT28), .Z(n527) );
  XNOR2_X1 U329 ( .A(n446), .B(G190GAT), .ZN(n447) );
  XNOR2_X1 U330 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT78), .B(KEYINPUT0), .Z(n290) );
  XNOR2_X1 U332 ( .A(G134GAT), .B(KEYINPUT80), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U334 ( .A(n291), .B(KEYINPUT79), .Z(n293) );
  XNOR2_X1 U335 ( .A(G113GAT), .B(G127GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n343) );
  XOR2_X1 U337 ( .A(G183GAT), .B(G176GAT), .Z(n295) );
  XNOR2_X1 U338 ( .A(G15GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U340 ( .A(n296), .B(G190GAT), .Z(n298) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G71GAT), .Z(n378) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(n378), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U344 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n300) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U347 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n304) );
  XNOR2_X1 U349 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(G169GAT), .B(n305), .Z(n439) );
  XNOR2_X1 U352 ( .A(n439), .B(KEYINPUT83), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n343), .B(n308), .ZN(n460) );
  XOR2_X1 U355 ( .A(G162GAT), .B(KEYINPUT73), .Z(n310) );
  XNOR2_X1 U356 ( .A(G50GAT), .B(G218GAT), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n351) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n311), .B(G211GAT), .ZN(n438) );
  XNOR2_X1 U360 ( .A(n351), .B(n438), .ZN(n326) );
  XOR2_X1 U361 ( .A(G141GAT), .B(G22GAT), .Z(n386) );
  XOR2_X1 U362 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n313) );
  XNOR2_X1 U363 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U365 ( .A(n386), .B(n314), .Z(n316) );
  NAND2_X1 U366 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U368 ( .A(G204GAT), .B(KEYINPUT86), .Z(n318) );
  XNOR2_X1 U369 ( .A(KEYINPUT84), .B(KEYINPUT24), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n320), .B(n319), .Z(n324) );
  XNOR2_X1 U372 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n321), .B(KEYINPUT2), .ZN(n338) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(G78GAT), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n322), .B(G148GAT), .ZN(n366) );
  XNOR2_X1 U376 ( .A(n338), .B(n366), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n468) );
  XOR2_X1 U379 ( .A(G57GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U380 ( .A(G1GAT), .B(G141GAT), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U382 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n330) );
  XNOR2_X1 U383 ( .A(KEYINPUT5), .B(KEYINPUT88), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U385 ( .A(n332), .B(n331), .Z(n337) );
  XOR2_X1 U386 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n334) );
  NAND2_X1 U387 ( .A1(G225GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U389 ( .A(KEYINPUT4), .B(n335), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U391 ( .A(G85GAT), .B(n338), .Z(n340) );
  XNOR2_X1 U392 ( .A(G29GAT), .B(G162GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U394 ( .A(n342), .B(n341), .Z(n345) );
  XNOR2_X1 U395 ( .A(n343), .B(G120GAT), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n518) );
  XOR2_X1 U397 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n347) );
  NAND2_X1 U398 ( .A1(G232GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U400 ( .A(n348), .B(KEYINPUT9), .Z(n353) );
  XOR2_X1 U401 ( .A(G29GAT), .B(G43GAT), .Z(n350) );
  XNOR2_X1 U402 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n394) );
  XNOR2_X1 U404 ( .A(n394), .B(n351), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U406 ( .A(G92GAT), .B(KEYINPUT65), .Z(n355) );
  XNOR2_X1 U407 ( .A(G134GAT), .B(G106GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U409 ( .A(n357), .B(n356), .Z(n359) );
  XOR2_X1 U410 ( .A(G36GAT), .B(G190GAT), .Z(n433) );
  XNOR2_X1 U411 ( .A(G99GAT), .B(G85GAT), .ZN(n379) );
  XOR2_X1 U412 ( .A(n433), .B(n379), .Z(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n551) );
  XOR2_X1 U414 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n361) );
  NAND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n363) );
  INV_X1 U417 ( .A(KEYINPUT31), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n369) );
  INV_X1 U419 ( .A(n369), .ZN(n368) );
  XOR2_X1 U420 ( .A(G176GAT), .B(G204GAT), .Z(n365) );
  XNOR2_X1 U421 ( .A(G64GAT), .B(G92GAT), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n436) );
  XNOR2_X1 U423 ( .A(n366), .B(n436), .ZN(n370) );
  INV_X1 U424 ( .A(n370), .ZN(n367) );
  NAND2_X1 U425 ( .A1(n368), .A2(n367), .ZN(n372) );
  NAND2_X1 U426 ( .A1(n370), .A2(n369), .ZN(n371) );
  NAND2_X1 U427 ( .A1(n372), .A2(n371), .ZN(n376) );
  XOR2_X1 U428 ( .A(G57GAT), .B(KEYINPUT13), .Z(n400) );
  XNOR2_X1 U429 ( .A(n400), .B(KEYINPUT71), .ZN(n374) );
  INV_X1 U430 ( .A(KEYINPUT33), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n380) );
  XOR2_X1 U432 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n382) );
  XNOR2_X1 U433 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n398) );
  XOR2_X1 U435 ( .A(G113GAT), .B(G36GAT), .Z(n384) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(G50GAT), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U438 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U439 ( .A1(G229GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U441 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n390) );
  XNOR2_X1 U442 ( .A(KEYINPUT67), .B(G8GAT), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U444 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U445 ( .A(G15GAT), .B(G1GAT), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n393), .B(KEYINPUT69), .ZN(n403) );
  XNOR2_X1 U447 ( .A(n394), .B(n403), .ZN(n395) );
  XNOR2_X1 U448 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U449 ( .A(n398), .B(n397), .ZN(n567) );
  NAND2_X1 U450 ( .A1(n558), .A2(n567), .ZN(n399) );
  XNOR2_X1 U451 ( .A(n399), .B(KEYINPUT46), .ZN(n418) );
  XOR2_X1 U452 ( .A(G8GAT), .B(G183GAT), .Z(n430) );
  XOR2_X1 U453 ( .A(n430), .B(n400), .Z(n402) );
  XNOR2_X1 U454 ( .A(G211GAT), .B(G155GAT), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n407) );
  XOR2_X1 U456 ( .A(n403), .B(KEYINPUT12), .Z(n405) );
  NAND2_X1 U457 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U459 ( .A(n407), .B(n406), .Z(n409) );
  XNOR2_X1 U460 ( .A(G127GAT), .B(G71GAT), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n409), .B(n408), .ZN(n417) );
  XOR2_X1 U462 ( .A(KEYINPUT76), .B(G64GAT), .Z(n411) );
  XNOR2_X1 U463 ( .A(G22GAT), .B(G78GAT), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U465 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n413) );
  XNOR2_X1 U466 ( .A(KEYINPUT15), .B(KEYINPUT74), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U468 ( .A(n415), .B(n414), .Z(n416) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n489) );
  NAND2_X1 U470 ( .A1(n418), .A2(n489), .ZN(n419) );
  NOR2_X1 U471 ( .A1(n551), .A2(n419), .ZN(n421) );
  XNOR2_X1 U472 ( .A(KEYINPUT47), .B(KEYINPUT107), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n427) );
  XOR2_X1 U474 ( .A(n551), .B(KEYINPUT36), .Z(n581) );
  NOR2_X1 U475 ( .A1(n581), .A2(n489), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n422), .B(KEYINPUT45), .ZN(n423) );
  NAND2_X1 U477 ( .A1(n423), .A2(n572), .ZN(n424) );
  NOR2_X1 U478 ( .A1(n567), .A2(n424), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n425), .B(KEYINPUT108), .ZN(n426) );
  NOR2_X1 U480 ( .A1(n427), .A2(n426), .ZN(n429) );
  XNOR2_X1 U481 ( .A(G218GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U482 ( .A(n431), .B(KEYINPUT91), .ZN(n432) );
  XOR2_X1 U483 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U484 ( .A1(G226GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U486 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U487 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U488 ( .A(n441), .B(n440), .ZN(n463) );
  NOR2_X1 U489 ( .A1(n449), .A2(n463), .ZN(n442) );
  XOR2_X1 U490 ( .A(n442), .B(KEYINPUT54), .Z(n443) );
  NOR2_X1 U491 ( .A1(n518), .A2(n443), .ZN(n565) );
  AND2_X1 U492 ( .A1(n468), .A2(n565), .ZN(n444) );
  XNOR2_X1 U493 ( .A(KEYINPUT55), .B(n444), .ZN(n445) );
  NAND2_X1 U494 ( .A1(n561), .A2(n551), .ZN(n448) );
  XOR2_X1 U495 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n446) );
  XNOR2_X1 U496 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n454) );
  INV_X1 U497 ( .A(n489), .ZN(n575) );
  INV_X1 U498 ( .A(n460), .ZN(n524) );
  XOR2_X1 U499 ( .A(n463), .B(KEYINPUT27), .Z(n470) );
  NAND2_X1 U500 ( .A1(n518), .A2(n470), .ZN(n459) );
  NOR2_X1 U501 ( .A1(n449), .A2(n459), .ZN(n542) );
  NAND2_X1 U502 ( .A1(n524), .A2(n542), .ZN(n450) );
  XOR2_X1 U503 ( .A(KEYINPUT109), .B(n450), .Z(n451) );
  NOR2_X1 U504 ( .A1(n451), .A2(n527), .ZN(n452) );
  XNOR2_X1 U505 ( .A(KEYINPUT110), .B(n452), .ZN(n537) );
  AND2_X1 U506 ( .A1(n575), .A2(n537), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n456) );
  INV_X1 U508 ( .A(G127GAT), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(G1342GAT) );
  XOR2_X1 U510 ( .A(KEYINPUT95), .B(KEYINPUT34), .Z(n479) );
  NAND2_X1 U511 ( .A1(n567), .A2(n572), .ZN(n492) );
  NOR2_X1 U512 ( .A1(n551), .A2(n489), .ZN(n457) );
  XOR2_X1 U513 ( .A(KEYINPUT16), .B(n457), .Z(n458) );
  XNOR2_X1 U514 ( .A(n458), .B(KEYINPUT77), .ZN(n477) );
  NOR2_X1 U515 ( .A1(n527), .A2(n459), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT92), .ZN(n476) );
  INV_X1 U518 ( .A(n463), .ZN(n521) );
  NAND2_X1 U519 ( .A1(n521), .A2(n524), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n464), .A2(n468), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT94), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT25), .B(n466), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n467), .B(KEYINPUT93), .ZN(n472) );
  NOR2_X1 U524 ( .A1(n468), .A2(n524), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT26), .ZN(n564) );
  NAND2_X1 U526 ( .A1(n470), .A2(n564), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n472), .A2(n471), .ZN(n474) );
  INV_X1 U528 ( .A(n518), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n488) );
  NAND2_X1 U531 ( .A1(n477), .A2(n488), .ZN(n505) );
  NOR2_X1 U532 ( .A1(n492), .A2(n505), .ZN(n486) );
  NAND2_X1 U533 ( .A1(n486), .A2(n518), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U536 ( .A1(n521), .A2(n486), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT35), .B(KEYINPUT97), .Z(n483) );
  NAND2_X1 U539 ( .A1(n486), .A2(n524), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n485) );
  XOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT96), .Z(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n486), .A2(n527), .ZN(n487) );
  XNOR2_X1 U544 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT98), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U546 ( .A1(n489), .A2(n488), .ZN(n490) );
  NOR2_X1 U547 ( .A1(n490), .A2(n581), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n491), .B(KEYINPUT37), .ZN(n517) );
  NOR2_X1 U549 ( .A1(n492), .A2(n517), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n493), .B(KEYINPUT38), .ZN(n501) );
  NAND2_X1 U551 ( .A1(n518), .A2(n501), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n501), .A2(n521), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT40), .Z(n499) );
  NAND2_X1 U557 ( .A1(n524), .A2(n501), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n501), .A2(n527), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n502), .B(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n503), .ZN(G1331GAT) );
  INV_X1 U563 ( .A(n567), .ZN(n504) );
  NAND2_X1 U564 ( .A1(n504), .A2(n558), .ZN(n516) );
  NOR2_X1 U565 ( .A1(n516), .A2(n505), .ZN(n506) );
  XOR2_X1 U566 ( .A(KEYINPUT101), .B(n506), .Z(n513) );
  NAND2_X1 U567 ( .A1(n513), .A2(n518), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n507), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n521), .A2(n513), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n511) );
  NAND2_X1 U573 ( .A1(n513), .A2(n524), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U577 ( .A1(n513), .A2(n527), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT104), .ZN(n520) );
  NOR2_X1 U580 ( .A1(n517), .A2(n516), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n518), .A2(n528), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  XOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT105), .Z(n523) );
  NAND2_X1 U584 ( .A1(n528), .A2(n521), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n528), .A2(n524), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n525), .B(KEYINPUT106), .ZN(n526) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n526), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U590 ( .A(n529), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n567), .A2(n537), .ZN(n532) );
  XOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT111), .Z(n531) );
  XNOR2_X1 U594 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n534) );
  NAND2_X1 U596 ( .A1(n558), .A2(n537), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT112), .Z(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U601 ( .A1(n551), .A2(n537), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT116), .Z(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n564), .A2(n542), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n543), .B(KEYINPUT117), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n552), .A2(n567), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U611 ( .A1(n552), .A2(n558), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U615 ( .A1(n552), .A2(n575), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n561), .A2(n567), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n556) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(n557), .Z(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n575), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(n563), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .Z(n569) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT124), .B(n566), .Z(n576) );
  NAND2_X1 U633 ( .A1(n576), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U638 ( .A(n576), .ZN(n580) );
  OR2_X1 U639 ( .A1(n572), .A2(n580), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n579) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1355GAT) );
endmodule

