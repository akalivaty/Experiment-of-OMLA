//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT64), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n453), .A2(G2106), .B1(KEYINPUT65), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  INV_X1    g040(.A(G113), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AND3_X1   g044(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n467), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  OAI221_X1 g057(.A(new_n481), .B1(new_n480), .B2(new_n479), .C1(G112), .C2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n472), .A2(new_n482), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n473), .A2(G136), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n482), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n470), .B2(new_n471), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(new_n494), .C1(new_n470), .C2(new_n471), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  XOR2_X1   g074(.A(KEYINPUT69), .B(KEYINPUT4), .Z(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n464), .A3(new_n494), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n492), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(G543), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n508), .A2(G62), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(G75), .A2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G88), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n514), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND2_X1  g094(.A1(new_n516), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n508), .A2(G89), .A3(new_n509), .A4(new_n514), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n508), .A2(G63), .A3(G651), .A4(new_n509), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n520), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  NAND2_X1  g101(.A1(new_n516), .A2(G52), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n508), .A2(G90), .A3(new_n509), .A4(new_n514), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n508), .A2(G64), .A3(new_n509), .ZN(new_n530));
  AND2_X1   g105(.A1(G77), .A2(G543), .ZN(new_n531));
  OAI21_X1  g106(.A(G651), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND4_X1  g109(.A1(new_n508), .A2(G81), .A3(new_n509), .A4(new_n514), .ZN(new_n535));
  INV_X1    g110(.A(G43), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n514), .A2(G543), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n508), .A2(G56), .A3(new_n509), .ZN(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR3_X1   g120(.A1(new_n538), .A2(new_n542), .A3(new_n544), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n516), .A2(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n513), .A2(new_n514), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G91), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n508), .A2(new_n509), .ZN(new_n560));
  XOR2_X1   g135(.A(KEYINPUT72), .B(G65), .Z(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n562), .A2(KEYINPUT73), .A3(G651), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(KEYINPUT73), .B1(new_n562), .B2(G651), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n556), .B(new_n558), .C1(new_n564), .C2(new_n565), .ZN(G299));
  OAI21_X1  g141(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n513), .A2(G87), .A3(new_n514), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n516), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(new_n557), .A2(G86), .ZN(new_n571));
  INV_X1    g146(.A(G48), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  OAI221_X1 g148(.A(new_n571), .B1(new_n572), .B2(new_n537), .C1(new_n539), .C2(new_n573), .ZN(G305));
  NAND2_X1  g149(.A1(new_n516), .A2(G47), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n513), .A2(new_n514), .ZN(new_n576));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OAI221_X1 g153(.A(new_n575), .B1(new_n576), .B2(new_n577), .C1(new_n578), .C2(new_n539), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n508), .A2(G92), .A3(new_n509), .A4(new_n514), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n516), .A2(G54), .ZN(new_n584));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n560), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(KEYINPUT74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n580), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n580), .B1(new_n593), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n464), .A2(new_n475), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT12), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(G2100), .Z(new_n609));
  NAND2_X1  g184(.A1(new_n484), .A2(G123), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n473), .A2(G135), .ZN(new_n611));
  OR2_X1    g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n612), .B(G2104), .C1(G111), .C2(new_n482), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n609), .A2(new_n615), .ZN(G156));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2430), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2435), .ZN(new_n618));
  XOR2_X1   g193(.A(G2427), .B(G2438), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT14), .ZN(new_n621));
  XOR2_X1   g196(.A(G2443), .B(G2446), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G1341), .B(G1348), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n623), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n627), .B(new_n628), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G14), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(G401));
  XOR2_X1   g206(.A(G2072), .B(G2078), .Z(new_n632));
  XOR2_X1   g207(.A(G2084), .B(G2090), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2067), .B(G2678), .Z(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n632), .B1(new_n636), .B2(KEYINPUT18), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT76), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n639), .A3(KEYINPUT17), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2096), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(G227));
  XOR2_X1   g220(.A(G1956), .B(G2474), .Z(new_n646));
  XOR2_X1   g221(.A(G1961), .B(G1966), .Z(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1971), .B(G1976), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT19), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n652), .B1(KEYINPUT20), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n655), .B(new_n656), .C1(KEYINPUT20), .C2(new_n654), .ZN(new_n657));
  XOR2_X1   g232(.A(G1991), .B(G1996), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT77), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1981), .B(G1986), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(G229));
  INV_X1    g241(.A(G16), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G23), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n669), .B2(new_n667), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT33), .Z(new_n671));
  OR2_X1    g246(.A1(new_n671), .A2(G1976), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(G6), .ZN(new_n673));
  INV_X1    g248(.A(G305), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n674), .B2(new_n667), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT32), .B(G1981), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT80), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(G1976), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n667), .A2(G22), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G166), .B2(new_n667), .ZN(new_n681));
  INV_X1    g256(.A(G1971), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND4_X1  g258(.A1(new_n672), .A2(new_n678), .A3(new_n679), .A4(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n667), .A2(G24), .ZN(new_n686));
  INV_X1    g261(.A(G290), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n667), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1986), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(KEYINPUT78), .A2(G29), .ZN(new_n691));
  NOR2_X1   g266(.A1(KEYINPUT78), .A2(G29), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G25), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n484), .A2(G119), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n473), .A2(G131), .ZN(new_n697));
  OR2_X1    g272(.A1(G95), .A2(G2105), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n698), .B(G2104), .C1(G107), .C2(new_n482), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n695), .B1(new_n701), .B2(new_n694), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT79), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(KEYINPUT81), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n684), .B2(KEYINPUT34), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n690), .B(new_n705), .C1(new_n707), .C2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT36), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n694), .A2(G35), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G162), .B2(new_n694), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT29), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(G2090), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT89), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(G2090), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT90), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(KEYINPUT89), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT24), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(G34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(G34), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n694), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n477), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G2084), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n614), .A2(KEYINPUT87), .A3(new_n694), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT30), .B(G28), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G16), .A2(G21), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G168), .B2(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G1966), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT87), .B1(new_n614), .B2(new_n694), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n728), .A2(new_n731), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(new_n482), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n473), .A2(G139), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n475), .A2(G103), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n738), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G29), .B2(G33), .ZN(new_n745));
  INV_X1    g320(.A(G2072), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G32), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n484), .A2(G129), .B1(G105), .B2(new_n475), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n473), .A2(G141), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n747), .B1(new_n753), .B2(G29), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  OAI22_X1  g330(.A1(new_n745), .A2(new_n746), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n733), .A2(G1966), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n736), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n745), .A2(new_n746), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT86), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n762));
  INV_X1    g337(.A(G26), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n693), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n694), .A2(KEYINPUT28), .A3(G26), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n484), .A2(G128), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n473), .A2(G140), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(new_n482), .B2(G116), .ZN(new_n768));
  INV_X1    g343(.A(G104), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n482), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(KEYINPUT84), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(KEYINPUT84), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n766), .B(new_n767), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n764), .B(new_n765), .C1(new_n774), .C2(new_n725), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n761), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G5), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G171), .B2(G16), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G1961), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n759), .A2(new_n760), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n758), .A2(new_n777), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G164), .A2(new_n694), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G27), .B2(new_n694), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G16), .A2(G19), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n548), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1341), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n720), .A2(new_n782), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n726), .A2(new_n727), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n779), .B2(G1961), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n754), .B2(new_n755), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT88), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n667), .A2(G20), .ZN(new_n795));
  OAI211_X1 g370(.A(KEYINPUT23), .B(new_n795), .C1(new_n597), .C2(new_n667), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(KEYINPUT23), .B2(new_n795), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n717), .A2(KEYINPUT90), .B1(new_n785), .B2(new_n784), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT82), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G4), .B2(G16), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n800), .A2(G4), .A3(G16), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n801), .B(new_n802), .C1(new_n592), .C2(new_n667), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT83), .B(G1348), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n798), .A2(new_n799), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT31), .B(G11), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n790), .A2(new_n794), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT91), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n711), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(G311));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT92), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n711), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(G150));
  NAND2_X1  g390(.A1(new_n516), .A2(G55), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n513), .A2(G93), .A3(new_n514), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n816), .B(new_n817), .C1(new_n818), .C2(new_n539), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G860), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT37), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n592), .A2(new_n600), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n513), .A2(G67), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n539), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n817), .A2(new_n816), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n545), .B2(new_n547), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n538), .A2(new_n542), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n819), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n824), .B(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n821), .B1(new_n834), .B2(G860), .ZN(G145));
  INV_X1    g410(.A(G37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n484), .A2(G130), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n473), .A2(G142), .ZN(new_n838));
  OR2_X1    g413(.A1(G106), .A2(G2105), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n839), .B(G2104), .C1(G118), .C2(new_n482), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n743), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n841), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n738), .A2(new_n739), .A3(new_n742), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n842), .A2(new_n700), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n700), .B1(new_n842), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n773), .A2(G164), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n773), .A2(G164), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n752), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n607), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n499), .A2(new_n501), .ZN(new_n855));
  INV_X1    g430(.A(new_n492), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n774), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n753), .A3(new_n850), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n854), .B1(new_n853), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n849), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n851), .A2(new_n852), .A3(new_n752), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n753), .B1(new_n858), .B2(new_n850), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n607), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n860), .A3(new_n848), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n477), .B(new_n487), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n614), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n868), .A2(KEYINPUT93), .A3(new_n870), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT93), .B1(new_n868), .B2(new_n870), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n836), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT94), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n868), .A2(new_n870), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT93), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n868), .A2(KEYINPUT93), .A3(new_n870), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT94), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n836), .A4(new_n871), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT95), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n602), .B(new_n833), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n562), .A2(G651), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT73), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n890), .A2(new_n563), .B1(G91), .B2(new_n557), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n556), .A3(new_n589), .ZN(new_n892));
  INV_X1    g467(.A(new_n589), .ZN(new_n893));
  NAND2_X1  g468(.A1(G299), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT41), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n887), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n887), .A2(new_n895), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n886), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n886), .B2(new_n900), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n669), .A2(G303), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n515), .A2(new_n517), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(G288), .A3(new_n512), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n906), .A3(G290), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G290), .B1(new_n904), .B2(new_n906), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n909), .A3(G305), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n687), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n674), .B1(new_n912), .B2(new_n907), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT42), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n903), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G868), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(G868), .B2(new_n829), .ZN(G295));
  OAI21_X1  g493(.A(new_n917), .B1(G868), .B2(new_n829), .ZN(G331));
  XNOR2_X1  g494(.A(G301), .B(G168), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n830), .B2(new_n832), .ZN(new_n921));
  XNOR2_X1  g496(.A(G301), .B(G286), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n831), .A2(KEYINPUT71), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n819), .B1(new_n923), .B2(new_n546), .ZN(new_n924));
  INV_X1    g499(.A(new_n832), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n897), .A3(new_n898), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n921), .A2(new_n926), .A3(new_n892), .A4(new_n894), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT98), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n914), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n928), .A2(new_n914), .A3(new_n931), .A4(new_n929), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n928), .A2(new_n914), .A3(new_n929), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT100), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n930), .B1(new_n910), .B2(new_n913), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n936), .A2(new_n937), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n938), .A2(new_n945), .A3(KEYINPUT44), .A4(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT99), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n930), .A2(new_n932), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(new_n836), .A3(new_n935), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n950), .B2(KEYINPUT43), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n941), .A2(new_n943), .A3(new_n934), .A4(new_n942), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n948), .A3(KEYINPUT43), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT97), .B(KEYINPUT44), .Z(new_n957));
  OAI21_X1  g532(.A(new_n947), .B1(new_n956), .B2(new_n957), .ZN(G397));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(G164), .B2(G1384), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n469), .A2(G40), .A3(new_n474), .A4(new_n476), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n773), .B(G2067), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT104), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n966), .B2(new_n753), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT46), .B1(new_n964), .B2(G1996), .ZN(new_n968));
  OR3_X1    g543(.A1(new_n964), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(G1996), .B2(new_n752), .ZN(new_n972));
  INV_X1    g547(.A(new_n964), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n964), .A2(new_n975), .A3(new_n753), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT103), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  OR3_X1    g553(.A1(new_n978), .A2(new_n700), .A3(new_n703), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n773), .A2(G2067), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n964), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n700), .B(new_n703), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT105), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n978), .B1(new_n973), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(G290), .A2(G1986), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(new_n964), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT48), .Z(new_n987));
  AOI211_X1 g562(.A(new_n971), .B(new_n981), .C1(new_n984), .C2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n573), .A2(new_n539), .ZN(new_n989));
  OAI21_X1  g564(.A(G1981), .B1(new_n989), .B2(KEYINPUT109), .ZN(new_n990));
  OR2_X1    g565(.A1(G305), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n992));
  NAND2_X1  g567(.A1(G305), .A2(new_n990), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(KEYINPUT49), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n963), .A2(new_n996), .A3(new_n857), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G8), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(KEYINPUT49), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n998), .B1(G1976), .B2(new_n669), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1002), .B(new_n1003), .C1(G1976), .C2(new_n669), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G303), .A2(G8), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT108), .B(KEYINPUT55), .Z(new_n1008));
  XNOR2_X1  g583(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n857), .A2(KEYINPUT45), .A3(new_n996), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(new_n959), .C1(G164), .C2(G1384), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n962), .B1(new_n960), .B2(KEYINPUT106), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n682), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n963), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n857), .A2(new_n1021), .A3(new_n996), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g599(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT107), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1020), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1011), .B1(new_n1018), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1006), .A2(new_n1010), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1001), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G288), .A2(G1976), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT111), .ZN(new_n1034));
  OAI22_X1  g609(.A1(new_n1032), .A2(new_n1034), .B1(G1981), .B2(G305), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n999), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1020), .A2(G2090), .A3(new_n1025), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n1017), .B2(new_n682), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1009), .B1(new_n1038), .B2(new_n1011), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1030), .A2(new_n1010), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1006), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n857), .A2(new_n996), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n962), .B1(new_n1042), .B2(KEYINPUT50), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1025), .A2(KEYINPUT107), .ZN(new_n1044));
  NOR4_X1   g619(.A1(G164), .A2(new_n1023), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1043), .B(new_n727), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1966), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n960), .B1(new_n1012), .B2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(G164), .A2(new_n959), .A3(G1384), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n963), .B1(new_n1052), .B2(KEYINPUT112), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1055), .A2(KEYINPUT113), .A3(new_n727), .A4(new_n1043), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1048), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(G8), .A3(G168), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT63), .B1(new_n1041), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1006), .A2(new_n1040), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT63), .B1(new_n1030), .B2(new_n1010), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1031), .B(new_n1036), .C1(new_n1060), .C2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1057), .A2(KEYINPUT120), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1048), .A2(new_n1066), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(G168), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1057), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n1071));
  NOR2_X1   g646(.A1(G168), .A2(new_n1011), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1072), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(KEYINPUT121), .A3(new_n1072), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT62), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1027), .A2(G1961), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(KEYINPUT53), .A3(new_n785), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1086), .A3(KEYINPUT122), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(KEYINPUT123), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(KEYINPUT123), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1089), .B(new_n1090), .C1(new_n1017), .C2(G2078), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  NOR4_X1   g667(.A1(new_n1051), .A2(new_n1053), .A3(new_n1088), .A4(G2078), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(new_n1083), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1087), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G171), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT121), .B1(new_n1076), .B2(new_n1072), .ZN(new_n1098));
  AOI211_X1 g673(.A(new_n1078), .B(new_n1073), .C1(new_n1065), .C2(new_n1067), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1082), .A2(new_n1097), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1956), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT114), .B(new_n1105), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT56), .B(G2072), .Z(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT116), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1015), .A2(new_n1016), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g689(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n891), .A2(new_n556), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(G299), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1118), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(new_n1108), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(KEYINPUT61), .A3(new_n1121), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1027), .A2(G1348), .B1(G2067), .B2(new_n997), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n592), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT61), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1016), .A2(new_n975), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1015), .A2(KEYINPUT117), .A3(new_n975), .A4(new_n1016), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n997), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1128), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1135), .ZN(new_n1137));
  AOI211_X1 g712(.A(KEYINPUT118), .B(new_n1137), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n548), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1123), .A2(new_n593), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1123), .A2(new_n593), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT60), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n548), .B(new_n1146), .C1(new_n1136), .C2(new_n1138), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1127), .A2(new_n1142), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1143), .A2(new_n1121), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n1149), .A3(new_n1119), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT53), .B(new_n785), .C1(new_n963), .C2(KEYINPUT124), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(KEYINPUT124), .B2(new_n963), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n960), .A3(new_n1012), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1084), .A2(new_n1091), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G171), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT54), .B(new_n1155), .C1(new_n1095), .C2(G171), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1154), .A2(G171), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT54), .B1(new_n1096), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1150), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1104), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1064), .B1(new_n1163), .B2(new_n1041), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT102), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n985), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(G290), .A2(G1986), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1166), .B(new_n1167), .Z(new_n1168));
  OAI21_X1  g743(.A(new_n984), .B1(new_n964), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n988), .B1(new_n1164), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n630), .A2(new_n665), .A3(new_n664), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1173), .B1(new_n875), .B2(new_n882), .ZN(new_n1174));
  NOR2_X1   g748(.A1(G227), .A2(new_n462), .ZN(new_n1175));
  AND4_X1   g749(.A1(KEYINPUT126), .A2(new_n1174), .A3(new_n955), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1177));
  AOI211_X1 g751(.A(KEYINPUT99), .B(new_n934), .C1(new_n933), .C2(new_n935), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n1178), .A2(new_n951), .ZN(new_n1179));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1179), .B2(new_n953), .ZN(new_n1180));
  AOI21_X1  g754(.A(KEYINPUT126), .B1(new_n1180), .B2(new_n1174), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n1172), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n1174), .A2(new_n955), .A3(new_n1175), .ZN(new_n1183));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g759(.A1(new_n1180), .A2(KEYINPUT126), .A3(new_n1174), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n1185), .A2(KEYINPUT127), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1182), .A2(new_n1187), .ZN(G308));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1186), .ZN(G225));
endmodule


