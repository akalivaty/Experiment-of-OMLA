//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G110), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT69), .B(G128), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n194), .A2(KEYINPUT23), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G128), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n191), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(G146), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n205), .B2(new_n208), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n199), .B1(new_n192), .B2(new_n193), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT24), .B(G110), .Z(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n201), .A2(new_n202), .A3(new_n213), .A4(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n211), .B2(new_n210), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT80), .B1(new_n219), .B2(new_n200), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n204), .A2(new_n207), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT82), .B1(new_n222), .B2(G146), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n204), .A2(new_n207), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n194), .A2(KEYINPUT23), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n197), .A2(new_n196), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n228), .A2(new_n191), .A3(new_n199), .A4(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n198), .A2(KEYINPUT81), .A3(new_n191), .A4(new_n199), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n215), .A2(new_n216), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n209), .B(new_n227), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n221), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(G221), .A3(G234), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(KEYINPUT22), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n242), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n221), .A2(new_n236), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n188), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n243), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n245), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n190), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n243), .A2(new_n245), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n189), .A2(G902), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G472), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT0), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n195), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n225), .A2(G143), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT64), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n257), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n225), .A2(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n260), .A2(G146), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n270), .A2(new_n271), .B1(new_n258), .B2(new_n195), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n272), .A2(KEYINPUT65), .A3(new_n265), .A4(new_n267), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n225), .B2(G143), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n260), .A2(KEYINPUT66), .A3(G146), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n261), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n264), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n241), .A2(KEYINPUT11), .A3(G134), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G137), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n282), .B2(G137), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n241), .A2(G134), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT67), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n285), .ZN(new_n290));
  AOI211_X1 g104(.A(G131), .B(new_n284), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G131), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n290), .ZN(new_n293));
  INV_X1    g107(.A(new_n284), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n274), .B(new_n280), .C1(new_n291), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n193), .A2(G116), .ZN(new_n297));
  INV_X1    g111(.A(G116), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n298), .A2(KEYINPUT71), .A3(G119), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT71), .B1(new_n298), .B2(G119), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT2), .B(G113), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n270), .A2(new_n271), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n195), .A2(KEYINPUT69), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G128), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(G143), .B2(new_n225), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n307), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n278), .A2(new_n312), .A3(G128), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n317), .B(new_n307), .C1(new_n311), .C2(new_n313), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n284), .B1(new_n287), .B2(new_n290), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n321));
  XNOR2_X1  g135(.A(G134), .B(G137), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(new_n292), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n288), .A2(new_n283), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT68), .A3(G131), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n320), .A2(new_n292), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n296), .A2(new_n306), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  INV_X1    g143(.A(G237), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT73), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G237), .ZN(new_n333));
  AOI21_X1  g147(.A(G953), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G210), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT27), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n338), .A3(G210), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n336), .B2(new_n339), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n329), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n342), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(G101), .A3(new_n340), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n328), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n296), .A2(new_n327), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT72), .A3(KEYINPUT30), .ZN(new_n348));
  OR2_X1    g162(.A1(KEYINPUT72), .A2(KEYINPUT30), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT72), .A2(KEYINPUT30), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n296), .A2(new_n327), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n346), .B1(new_n352), .B2(new_n305), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT31), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n256), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n306), .B1(new_n348), .B2(new_n351), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT74), .B(KEYINPUT31), .C1(new_n356), .C2(new_n346), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n352), .A2(new_n305), .ZN(new_n359));
  INV_X1    g173(.A(new_n346), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n328), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n347), .A2(new_n305), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n296), .A2(new_n327), .A3(new_n306), .A4(KEYINPUT28), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n343), .A2(new_n345), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n366), .A2(KEYINPUT75), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT75), .B1(new_n366), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n361), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n255), .B(new_n188), .C1(new_n358), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n366), .A2(new_n367), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(KEYINPUT75), .A3(new_n367), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n378), .A2(new_n355), .A3(new_n361), .A4(new_n357), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n379), .A2(KEYINPUT76), .A3(new_n255), .A4(new_n188), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT32), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n379), .A2(KEYINPUT32), .A3(new_n255), .A4(new_n188), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n328), .A2(KEYINPUT78), .A3(new_n362), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT78), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n363), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n364), .A2(KEYINPUT77), .A3(new_n328), .ZN(new_n388));
  OR3_X1    g202(.A1(new_n347), .A2(KEYINPUT77), .A3(new_n305), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n385), .B(new_n387), .C1(new_n390), .C2(new_n362), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(new_n367), .ZN(new_n393));
  INV_X1    g207(.A(new_n367), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n359), .B2(new_n328), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n392), .B1(new_n366), .B2(new_n367), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n188), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G472), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n384), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n254), .B1(new_n383), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g215(.A(KEYINPUT9), .B(G234), .Z(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G221), .B1(new_n403), .B2(G902), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G140), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n238), .A2(G227), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n313), .A2(new_n195), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n316), .B1(new_n278), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G104), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G107), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n412), .A2(G107), .ZN(new_n415));
  OAI21_X1  g229(.A(G101), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT3), .B1(new_n412), .B2(G107), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT3), .ZN(new_n418));
  INV_X1    g232(.A(G107), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(G104), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n417), .A2(new_n420), .A3(new_n329), .A4(new_n413), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n411), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n319), .B2(new_n423), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n291), .A2(new_n295), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n425), .A2(KEYINPUT12), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT12), .B1(new_n425), .B2(new_n427), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT10), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n269), .A2(new_n273), .B1(new_n279), .B2(new_n278), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n417), .A2(new_n420), .A3(new_n413), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G101), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(G101), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT4), .A3(new_n421), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n433), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n319), .A2(KEYINPUT10), .A3(new_n423), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n432), .A2(new_n439), .A3(new_n426), .A4(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n409), .B1(new_n430), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n432), .A2(new_n439), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n427), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n441), .A3(new_n408), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(KEYINPUT83), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT83), .B1(new_n443), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g263(.A(G469), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G469), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n441), .A2(new_n408), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n430), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n408), .B1(new_n445), .B2(new_n441), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n451), .B(new_n188), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(G469), .A2(G902), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n405), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n334), .A2(G214), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n260), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n334), .A2(G143), .A3(G214), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT18), .A2(G131), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT87), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT87), .B1(new_n204), .B2(new_n207), .ZN(new_n468));
  OAI21_X1  g282(.A(G146), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n227), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n292), .B1(new_n462), .B2(new_n463), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT18), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n222), .A2(KEYINPUT19), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n222), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n466), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n477), .B2(KEYINPUT19), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n210), .B1(new_n478), .B2(new_n225), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n334), .A2(G143), .A3(G214), .ZN(new_n480));
  AOI21_X1  g294(.A(G143), .B1(new_n334), .B2(G214), .ZN(new_n481));
  OAI21_X1  g295(.A(G131), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n462), .A2(new_n292), .A3(new_n463), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n471), .A2(new_n473), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n412), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n460), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n472), .A2(KEYINPUT17), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n212), .C1(new_n484), .C2(KEYINPUT17), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT18), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n470), .B(new_n465), .C1(new_n482), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n479), .A2(new_n484), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n492), .ZN(new_n495));
  INV_X1    g309(.A(new_n487), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(KEYINPUT88), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n488), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G475), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n188), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n499), .A4(new_n188), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n490), .A2(new_n492), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(new_n496), .ZN(new_n507));
  AOI211_X1 g321(.A(KEYINPUT89), .B(new_n487), .C1(new_n490), .C2(new_n492), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n493), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n499), .B1(new_n509), .B2(new_n188), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G952), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(G953), .ZN(new_n513));
  NAND2_X1  g327(.A1(G234), .A2(G237), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT21), .B(G898), .Z(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(G902), .A3(G953), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n195), .A2(G143), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT13), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n523), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n192), .B2(new_n260), .ZN(new_n527));
  OAI211_X1 g341(.A(G134), .B(new_n525), .C1(new_n527), .C2(new_n524), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n282), .B(new_n526), .C1(new_n192), .C2(new_n260), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n298), .A2(G122), .ZN(new_n530));
  INV_X1    g344(.A(G122), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(G116), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n419), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(G116), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n298), .A2(G122), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(G107), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n528), .A2(new_n529), .A3(new_n533), .A4(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n260), .B1(new_n308), .B2(new_n310), .ZN(new_n538));
  OAI21_X1  g352(.A(G134), .B1(new_n538), .B2(new_n523), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n529), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n534), .A2(KEYINPUT14), .A3(G107), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n533), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT14), .A4(G107), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT90), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT90), .B1(new_n547), .B2(new_n540), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n537), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n403), .A2(new_n187), .A3(G953), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n537), .B(new_n550), .C1(new_n546), .C2(new_n548), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT91), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G478), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(KEYINPUT15), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n556), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n511), .A2(new_n522), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G214), .B1(G237), .B2(G902), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n433), .A2(new_n206), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n319), .A2(G125), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT86), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G224), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G953), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT86), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n433), .B2(new_n206), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n565), .B2(new_n570), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(G110), .B(G122), .Z(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n305), .A2(new_n436), .A3(new_n438), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT5), .B(new_n297), .C1(new_n299), .C2(new_n300), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n297), .A2(KEYINPUT5), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(G113), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT84), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n577), .A2(new_n581), .A3(G113), .A4(new_n578), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n580), .A2(new_n303), .A3(new_n423), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT85), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT85), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n576), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n575), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n584), .A2(new_n574), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT6), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n587), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n586), .B1(new_n576), .B2(new_n583), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n574), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT6), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n573), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n580), .A2(new_n303), .A3(new_n422), .A4(new_n582), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n303), .A2(new_n579), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n423), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n574), .B(KEYINPUT8), .Z(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n565), .A2(new_n570), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n568), .A2(KEYINPUT7), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n589), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n603), .B2(new_n604), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n188), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G210), .B1(G237), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n596), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n571), .A2(new_n572), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n594), .B1(new_n593), .B2(new_n607), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n588), .A2(KEYINPUT6), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n603), .ZN(new_n617));
  INV_X1    g431(.A(new_n604), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n589), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n619), .B2(new_n605), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n610), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n562), .B1(new_n612), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n459), .A2(new_n561), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n401), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NAND2_X1  g439(.A1(new_n379), .A2(new_n188), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G472), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n381), .A2(new_n253), .A3(new_n458), .A4(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT92), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n373), .A2(new_n380), .B1(G472), .B2(new_n626), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(KEYINPUT92), .A3(new_n253), .A4(new_n458), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT94), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n553), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n553), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n544), .A2(new_n545), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n547), .A2(KEYINPUT90), .A3(new_n540), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n550), .B1(new_n639), .B2(new_n537), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n635), .B(KEYINPUT33), .C1(new_n636), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n552), .B(new_n553), .C1(new_n634), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(G478), .A3(new_n188), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n557), .A2(KEYINPUT95), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n557), .A2(KEYINPUT95), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n554), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n651), .B(new_n522), .C1(new_n504), .C2(new_n510), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n562), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT93), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n612), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n611), .B1(new_n596), .B2(new_n609), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n616), .A2(new_n610), .A3(new_n620), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT93), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n633), .A2(new_n653), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NAND2_X1  g477(.A1(new_n509), .A2(new_n188), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G475), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n502), .A3(new_n503), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n560), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n660), .A2(new_n522), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n633), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  OAI21_X1  g486(.A(new_n237), .B1(KEYINPUT36), .B2(new_n242), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n242), .A2(KEYINPUT36), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n221), .A2(new_n236), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n673), .A2(new_n252), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT96), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT96), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n673), .A2(new_n678), .A3(new_n252), .A4(new_n675), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n250), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n561), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n631), .A3(new_n683), .A4(new_n458), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT37), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n191), .ZN(G12));
  OR2_X1    g500(.A1(new_n250), .A2(new_n680), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT32), .B1(new_n373), .B2(new_n380), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n458), .B(new_n687), .C1(new_n688), .C2(new_n399), .ZN(new_n689));
  INV_X1    g503(.A(new_n660), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n516), .B1(new_n520), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT97), .B1(new_n667), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT97), .ZN(new_n696));
  NOR4_X1   g510(.A1(new_n666), .A2(new_n696), .A3(new_n560), .A4(new_n693), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  NOR2_X1   g514(.A1(new_n612), .A2(new_n621), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT38), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(KEYINPUT38), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n704), .A2(new_n654), .A3(new_n687), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n693), .B(KEYINPUT39), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n458), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT40), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n511), .A2(new_n560), .ZN(new_n711));
  INV_X1    g525(.A(new_n353), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n390), .B2(new_n394), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(new_n188), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n383), .B(new_n384), .C1(new_n255), .C2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n705), .A2(new_n710), .A3(new_n711), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(new_n689), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n651), .B(new_n694), .C1(new_n504), .C2(new_n510), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT98), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n666), .A2(KEYINPUT98), .A3(new_n651), .A4(new_n694), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n718), .A2(new_n660), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  OAI21_X1  g539(.A(new_n188), .B1(new_n453), .B2(new_n454), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n455), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n405), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n253), .B(new_n729), .C1(new_n688), .C2(new_n399), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n660), .A2(new_n653), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT41), .B(G113), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NOR2_X1   g548(.A1(new_n730), .A2(new_n668), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n298), .ZN(G18));
  AND3_X1   g550(.A1(new_n656), .A2(new_n729), .A3(new_n659), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n682), .B(new_n737), .C1(new_n688), .C2(new_n399), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  AOI22_X1  g553(.A1(new_n391), .A2(new_n367), .B1(new_n354), .B2(new_n353), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n712), .A2(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n255), .A3(new_n188), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n253), .A2(new_n627), .A3(new_n743), .A4(new_n522), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n660), .A3(new_n711), .A4(new_n729), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  AOI21_X1  g560(.A(G472), .B1(new_n740), .B2(new_n741), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n747), .A2(new_n188), .B1(new_n626), .B2(G472), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n721), .A3(new_n687), .A4(new_n722), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n656), .A2(new_n729), .A3(new_n659), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT99), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT99), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n687), .A2(new_n627), .A3(new_n743), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n723), .A2(new_n752), .A3(new_n737), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  OAI21_X1  g570(.A(new_n253), .B1(new_n688), .B2(new_n399), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n657), .A2(new_n658), .A3(new_n562), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT100), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT100), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n657), .A2(new_n658), .A3(new_n760), .A4(new_n562), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n443), .A2(new_n446), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(G469), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n405), .B1(new_n457), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n759), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n721), .A2(new_n767), .A3(new_n722), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n757), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n759), .A2(new_n761), .A3(new_n765), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n371), .A2(new_n382), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n384), .A3(new_n398), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n772), .A2(KEYINPUT101), .A3(new_n253), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT101), .B1(new_n772), .B2(new_n253), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n723), .B(new_n770), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n769), .B1(new_n775), .B2(KEYINPUT42), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  INV_X1    g591(.A(KEYINPUT102), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n695), .B2(new_n697), .ZN(new_n779));
  INV_X1    g593(.A(new_n697), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n502), .A2(new_n503), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n556), .B(new_n558), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n665), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n696), .B1(new_n783), .B2(new_n693), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n784), .A3(KEYINPUT102), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n401), .A2(new_n779), .A3(new_n785), .A4(new_n770), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  INV_X1    g601(.A(new_n455), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n763), .A2(KEYINPUT45), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT83), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n762), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n447), .ZN(new_n792));
  OAI211_X1 g606(.A(G469), .B(new_n789), .C1(new_n792), .C2(KEYINPUT45), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n456), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n788), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(KEYINPUT46), .A3(new_n456), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n405), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n707), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT103), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n759), .A2(new_n761), .ZN(new_n801));
  INV_X1    g615(.A(new_n631), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n511), .A2(new_n651), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n804));
  AOI21_X1  g618(.A(G902), .B1(new_n641), .B2(new_n643), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n649), .B1(new_n805), .B2(G478), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT104), .B1(new_n666), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n802), .A2(new_n687), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT44), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT44), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n801), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n800), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  NAND2_X1  g629(.A1(new_n794), .A2(new_n795), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n816), .A2(new_n455), .A3(new_n797), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT47), .B1(new_n817), .B2(new_n405), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n688), .A2(new_n399), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n798), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n759), .A2(new_n761), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n723), .A2(new_n254), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n818), .A2(new_n819), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  NAND3_X1  g639(.A1(new_n822), .A2(KEYINPUT113), .A3(new_n729), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  INV_X1    g641(.A(new_n729), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n827), .B1(new_n801), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n515), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n804), .A2(new_n809), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n773), .A2(new_n774), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n833), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n835), .A3(new_n836), .A4(new_n831), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(KEYINPUT48), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n715), .A2(new_n254), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(new_n830), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n806), .B1(new_n781), .B2(new_n665), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n513), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT48), .B1(new_n834), .B2(new_n837), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n840), .A2(new_n511), .A3(new_n806), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT114), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n840), .A2(new_n848), .A3(new_n511), .A4(new_n806), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n830), .A2(new_n753), .A3(new_n831), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n804), .A2(new_n809), .A3(new_n516), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n748), .A2(new_n253), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT112), .B1(new_n857), .B2(new_n801), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n855), .A2(new_n859), .A3(new_n856), .A4(new_n822), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n728), .A2(new_n404), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n818), .B2(new_n821), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n853), .B(new_n854), .C1(new_n861), .C2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n857), .A2(new_n828), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n654), .A3(new_n704), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT50), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n850), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n851), .A2(new_n852), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n871), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n850), .A2(new_n865), .A3(new_n869), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n845), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n660), .A2(new_n711), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT109), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n681), .B2(new_n694), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n250), .A2(new_n680), .A3(KEYINPUT109), .A4(new_n693), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n715), .A3(new_n765), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n699), .A2(new_n724), .A3(new_n755), .A4(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT110), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n622), .A2(new_n783), .A3(new_n521), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n630), .A2(new_n632), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n684), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n841), .A2(KEYINPUT106), .A3(new_n522), .A4(new_n683), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT106), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n622), .B2(new_n652), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n630), .A2(new_n632), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n624), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n895), .A2(KEYINPUT107), .A3(new_n624), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n890), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT108), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n749), .B2(new_n766), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n723), .A2(new_n770), .A3(KEYINPUT108), .A4(new_n753), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n666), .A2(new_n782), .A3(new_n693), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n822), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n718), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n904), .A2(new_n907), .A3(new_n786), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT52), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n887), .A2(new_n900), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n745), .B1(new_n731), .B2(new_n730), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n738), .B1(new_n730), .B2(new_n668), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n776), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n691), .B1(new_n698), .B2(new_n723), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n886), .A3(new_n755), .A4(new_n882), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n776), .A3(new_n913), .ZN(new_n919));
  INV_X1    g733(.A(new_n890), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT107), .B1(new_n895), .B2(new_n624), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n895), .A2(KEYINPUT107), .A3(new_n624), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n908), .B(new_n920), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n883), .A2(KEYINPUT52), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n919), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI221_X1 g739(.A(KEYINPUT54), .B1(new_n910), .B2(new_n916), .C1(new_n915), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n866), .A2(new_n660), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n776), .A2(new_n913), .A3(KEYINPUT111), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT111), .B1(new_n776), .B2(new_n913), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n915), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT52), .B1(new_n883), .B2(new_n884), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n923), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n932), .A3(new_n909), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n900), .A2(new_n914), .A3(new_n918), .A4(new_n908), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n915), .B1(new_n934), .B2(new_n924), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT54), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n875), .A2(new_n926), .A3(new_n927), .A4(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(G952), .A2(G953), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT117), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n728), .A2(KEYINPUT49), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n253), .A2(new_n562), .A3(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n943), .A2(new_n803), .A3(new_n405), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT105), .Z(new_n945));
  OAI21_X1  g759(.A(new_n704), .B1(KEYINPUT49), .B2(new_n728), .ZN(new_n946));
  OR3_X1    g760(.A1(new_n945), .A2(new_n715), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n941), .A2(new_n947), .ZN(G75));
  NOR2_X1   g762(.A1(new_n614), .A2(new_n615), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n613), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT55), .Z(new_n951));
  AOI21_X1  g765(.A(new_n188), .B1(new_n933), .B2(new_n935), .ZN(new_n952));
  AOI211_X1 g766(.A(KEYINPUT56), .B(new_n951), .C1(new_n952), .C2(G210), .ZN(new_n953));
  INV_X1    g767(.A(new_n951), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n933), .A2(new_n935), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(G210), .A3(G902), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT56), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n238), .A2(G952), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n953), .A2(new_n958), .A3(new_n959), .ZN(G51));
  XOR2_X1   g774(.A(new_n456), .B(KEYINPUT57), .Z(new_n961));
  AND3_X1   g775(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n936), .B1(new_n933), .B2(new_n935), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n453), .A2(new_n454), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n933), .A2(new_n935), .ZN(new_n967));
  OR3_X1    g781(.A1(new_n967), .A2(new_n188), .A3(new_n793), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n959), .B1(new_n966), .B2(new_n968), .ZN(G54));
  INV_X1    g783(.A(new_n959), .ZN(new_n970));
  NAND2_X1  g784(.A1(KEYINPUT58), .A2(G475), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n188), .B(new_n971), .C1(new_n933), .C2(new_n935), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n972), .B2(new_n498), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n952), .A2(KEYINPUT58), .A3(G475), .A4(new_n498), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT118), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT118), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n972), .A2(new_n976), .A3(new_n498), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n973), .B1(new_n975), .B2(new_n977), .ZN(G60));
  OAI22_X1  g792(.A1(new_n925), .A2(new_n915), .B1(new_n910), .B2(new_n916), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n937), .B1(new_n979), .B2(new_n936), .ZN(new_n980));
  NAND2_X1  g794(.A1(G478), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT59), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n644), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n644), .A2(new_n983), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n955), .A2(KEYINPUT54), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n937), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n984), .A2(new_n959), .A3(new_n987), .ZN(G63));
  XNOR2_X1  g802(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n673), .A2(new_n675), .ZN(new_n991));
  NAND2_X1  g805(.A1(G217), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT119), .Z(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT60), .Z(new_n994));
  NAND3_X1  g808(.A1(new_n955), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n970), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n251), .B(KEYINPUT120), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n955), .B2(new_n994), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n990), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n994), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n997), .B1(new_n967), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(new_n970), .A3(new_n989), .A4(new_n995), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1000), .A2(new_n1003), .ZN(G66));
  NAND2_X1  g818(.A1(new_n900), .A2(new_n913), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n238), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT122), .Z(new_n1007));
  OAI21_X1  g821(.A(G953), .B1(new_n518), .B2(new_n566), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n949), .B1(G898), .B2(new_n238), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G69));
  NOR2_X1   g825(.A1(new_n692), .A2(new_n238), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n352), .B(new_n478), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n833), .A2(new_n876), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n800), .B1(new_n1015), .B2(new_n813), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n917), .A2(new_n755), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n824), .A2(new_n776), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1016), .A2(new_n786), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n1013), .B(new_n1014), .C1(new_n1019), .C2(G953), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT124), .ZN(new_n1021));
  INV_X1    g835(.A(new_n708), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n783), .B1(new_n511), .B2(new_n806), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n401), .A2(new_n1022), .A3(new_n822), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1021), .B1(new_n814), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1024), .ZN(new_n1026));
  AOI211_X1 g840(.A(KEYINPUT124), .B(new_n1026), .C1(new_n800), .C2(new_n813), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n824), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1017), .A2(KEYINPUT62), .A3(new_n716), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n917), .A2(new_n716), .A3(new_n755), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT62), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1029), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(G953), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1014), .B(KEYINPUT123), .Z(new_n1036));
  OAI21_X1  g850(.A(new_n1020), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n238), .B1(G227), .B2(G900), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1038), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n1040), .B(new_n1020), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1039), .A2(new_n1041), .ZN(G72));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  OAI21_X1  g858(.A(new_n1044), .B1(new_n1019), .B2(new_n1005), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n359), .A2(new_n328), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT126), .Z(new_n1047));
  NAND3_X1  g861(.A1(new_n1045), .A2(new_n367), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1044), .B1(new_n395), .B2(new_n353), .ZN(new_n1049));
  XOR2_X1   g863(.A(new_n1049), .B(KEYINPUT127), .Z(new_n1050));
  OAI211_X1 g864(.A(new_n1048), .B(new_n970), .C1(new_n979), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1005), .ZN(new_n1052));
  OAI211_X1 g866(.A(new_n1052), .B(new_n1034), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1053));
  AND3_X1   g867(.A1(new_n1053), .A2(KEYINPUT125), .A3(new_n1044), .ZN(new_n1054));
  AOI21_X1  g868(.A(KEYINPUT125), .B1(new_n1053), .B2(new_n1044), .ZN(new_n1055));
  NOR3_X1   g869(.A1(new_n1054), .A2(new_n1055), .A3(new_n1047), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1051), .B1(new_n1056), .B2(new_n394), .ZN(G57));
endmodule


