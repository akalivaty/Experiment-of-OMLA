//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n205), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n208), .B1(new_n212), .B2(new_n213), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(new_n216), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n215), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT66), .B(G50), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n245), .A2(new_n209), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n244), .A2(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G68), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n209), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR3_X1   g0056(.A1(KEYINPUT70), .A2(G20), .A3(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G77), .ZN(new_n263));
  INV_X1    g0063(.A(G20), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G68), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n254), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT11), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n249), .B1(new_n251), .B2(new_n253), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n266), .A2(new_n267), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT76), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  AND2_X1   g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n209), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n276), .A2(KEYINPUT67), .A3(G1), .A4(G13), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G41), .A2(G45), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G1), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n275), .A2(G274), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n278), .B2(G1), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n244), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n275), .A2(new_n282), .A3(new_n277), .A4(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G238), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n288), .A2(new_n290), .A3(G232), .A4(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT73), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n294), .A2(KEYINPUT73), .A3(G232), .A4(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G97), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(G226), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n293), .A2(new_n295), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n274), .A2(new_n209), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n299), .A2(KEYINPUT74), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT74), .B1(new_n299), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n287), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT13), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT13), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n305), .B(new_n287), .C1(new_n301), .C2(new_n302), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(G179), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n306), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n308), .A3(new_n312), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n272), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n307), .A2(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n317));
  INV_X1    g0117(.A(new_n312), .ZN(new_n318));
  AOI211_X1 g0118(.A(KEYINPUT14), .B(new_n318), .C1(new_n304), .C2(new_n306), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n317), .A2(KEYINPUT76), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n271), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n270), .B1(new_n310), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n304), .B2(new_n306), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G226), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n280), .B1(new_n284), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT69), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n294), .A2(G222), .A3(new_n297), .ZN(new_n333));
  INV_X1    g0133(.A(G77), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n294), .A2(G1698), .ZN(new_n335));
  INV_X1    g0135(.A(G223), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n333), .B1(new_n334), .B2(new_n294), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n300), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(new_n331), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n332), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n340), .A2(G179), .ZN(new_n341));
  INV_X1    g0141(.A(new_n251), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n259), .B1(new_n244), .B2(G20), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n342), .A2(new_n343), .B1(new_n259), .B2(new_n246), .ZN(new_n344));
  INV_X1    g0144(.A(new_n258), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT8), .B(G58), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n345), .A2(G150), .B1(new_n262), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n264), .B1(new_n201), .B2(new_n259), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT71), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n254), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n344), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n340), .A2(new_n311), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n341), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n353), .B(KEYINPUT9), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n340), .A2(G200), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n356), .B(new_n357), .C1(new_n322), .C2(new_n340), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT18), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n289), .A2(KEYINPUT77), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT3), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n365), .A3(G33), .ZN(new_n366));
  AOI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n288), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n247), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n288), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(G33), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT7), .B1(new_n372), .B2(G20), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n215), .A2(new_n247), .ZN(new_n375));
  OAI21_X1  g0175(.A(G20), .B1(new_n375), .B2(new_n201), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n258), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(KEYINPUT16), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n368), .A2(G20), .ZN(new_n382));
  AOI21_X1  g0182(.A(G33), .B1(new_n363), .B2(new_n365), .ZN(new_n383));
  INV_X1    g0183(.A(new_n290), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n368), .B1(new_n294), .B2(G20), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n247), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n381), .B1(new_n387), .B2(new_n378), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n380), .A2(new_n254), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT78), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n346), .A2(new_n246), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n347), .A2(new_n252), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n390), .B(new_n391), .C1(new_n392), .C2(new_n251), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n342), .A2(new_n252), .A3(new_n347), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n390), .B1(new_n395), .B2(new_n391), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT79), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n391), .B1(new_n392), .B2(new_n251), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT78), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n393), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n389), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n280), .B1(new_n284), .B2(new_n216), .ZN(new_n404));
  INV_X1    g0204(.A(new_n300), .ZN(new_n405));
  NOR2_X1   g0205(.A1(G223), .A2(G1698), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n329), .B2(G1698), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n366), .A3(new_n288), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G169), .ZN(new_n412));
  INV_X1    g0212(.A(G179), .ZN(new_n413));
  OR3_X1    g0213(.A1(new_n404), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n362), .B1(new_n403), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n403), .A2(new_n362), .A3(new_n415), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n404), .A2(new_n410), .A3(new_n322), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(G200), .B2(new_n411), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(new_n389), .A3(new_n402), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n378), .B1(new_n369), .B2(new_n373), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n352), .B1(new_n424), .B2(KEYINPUT16), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n388), .B1(new_n397), .B2(new_n401), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n420), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n417), .A2(new_n418), .A3(new_n423), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n335), .A2(new_n285), .B1(new_n217), .B2(new_n294), .ZN(new_n430));
  INV_X1    g0230(.A(new_n294), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n431), .A2(new_n216), .A3(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n300), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G244), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n284), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n280), .A3(new_n435), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n436), .A2(KEYINPUT72), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G190), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n252), .A2(G77), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n251), .A2(new_n441), .B1(G77), .B2(new_n245), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n345), .A2(new_n347), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n442), .B1(new_n447), .B2(new_n254), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n440), .B(new_n448), .C1(new_n324), .C2(new_n439), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n439), .B2(new_n413), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n437), .A2(new_n311), .A3(new_n438), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n361), .A2(new_n429), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n217), .B1(new_n385), .B2(new_n386), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT6), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n455), .A2(new_n456), .A3(G107), .ZN(new_n457));
  XNOR2_X1  g0257(.A(G97), .B(G107), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n459), .A2(new_n264), .B1(new_n334), .B2(new_n258), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n254), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n246), .A2(new_n456), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  OR3_X1    g0263(.A1(new_n261), .A2(KEYINPUT80), .A3(G1), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT80), .B1(new_n261), .B2(G1), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n342), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n465), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT81), .B1(new_n467), .B2(new_n251), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n468), .A3(G97), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n461), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n366), .A2(G244), .A3(new_n297), .A4(new_n288), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT4), .A2(G244), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n288), .A2(new_n290), .A3(new_n475), .A4(new_n297), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n288), .A2(new_n290), .A3(G250), .A4(G1698), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n275), .A2(new_n277), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n244), .A2(G45), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(G41), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n481), .A2(new_n300), .B1(new_n489), .B2(G257), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n488), .A2(G274), .A3(new_n275), .A4(new_n277), .ZN(new_n491));
  AOI21_X1  g0291(.A(G200), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(G257), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n479), .B1(new_n473), .B2(new_n472), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n491), .C1(new_n494), .C2(new_n405), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G190), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n471), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n490), .A2(new_n322), .A3(new_n491), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n324), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n502), .A3(new_n471), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n495), .A2(new_n311), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n481), .A2(new_n300), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(new_n413), .A3(new_n493), .A4(new_n491), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n505), .A2(new_n507), .A3(new_n470), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(G238), .A2(G1698), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n434), .B2(G1698), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(new_n366), .A3(new_n288), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n512), .B2(new_n514), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n516), .A2(new_n517), .A3(new_n405), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT83), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n483), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n244), .A2(KEYINPUT83), .A3(G45), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n520), .A2(G250), .A3(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(KEYINPUT84), .A3(new_n275), .A4(new_n277), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT84), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(G250), .A3(new_n521), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n482), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n275), .A2(G274), .A3(new_n277), .ZN(new_n528));
  INV_X1    g0328(.A(G45), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(G1), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(G200), .B1(new_n518), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n517), .A2(new_n405), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n515), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n523), .A2(new_n526), .B1(new_n530), .B2(new_n528), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(G190), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n262), .A2(new_n538), .A3(G97), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  INV_X1    g0340(.A(G87), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n540), .A2(new_n541), .B1(new_n296), .B2(new_n264), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n539), .B1(new_n542), .B2(new_n538), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n366), .A2(new_n264), .A3(G68), .A4(new_n288), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n254), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n444), .A2(new_n246), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n466), .A2(new_n468), .A3(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT87), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n466), .A2(new_n468), .A3(new_n551), .A4(G87), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n533), .A2(new_n537), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n311), .B1(new_n518), .B2(new_n532), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n535), .A2(new_n413), .A3(new_n536), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n444), .B(KEYINPUT86), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n468), .A3(new_n466), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n546), .A3(new_n547), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n504), .A2(new_n509), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n487), .ZN(new_n564));
  NOR2_X1   g0364(.A1(KEYINPUT5), .A2(G41), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n530), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n566), .A2(new_n275), .A3(G270), .A4(new_n277), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n491), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT88), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT88), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n491), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n218), .A2(new_n297), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n366), .A2(new_n288), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT89), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n431), .A2(G303), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n366), .A2(G257), .A3(new_n297), .A4(new_n288), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n366), .A2(KEYINPUT89), .A3(new_n288), .A4(new_n573), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n300), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n572), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT90), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n572), .A2(new_n581), .A3(KEYINPUT90), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n342), .A2(G116), .A3(new_n464), .A4(new_n465), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n586), .B(KEYINPUT91), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n478), .B(new_n264), .C1(G33), .C2(new_n456), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n254), .C1(new_n264), .C2(G116), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT92), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n245), .B2(G116), .ZN(new_n594));
  INV_X1    g0394(.A(G116), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n246), .A2(KEYINPUT92), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n591), .A2(new_n592), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n311), .B1(new_n587), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n584), .A2(new_n585), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n584), .A2(new_n601), .A3(new_n585), .A4(new_n598), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT23), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n604), .A2(new_n264), .A3(G107), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT23), .B1(new_n217), .B2(G20), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n605), .A2(new_n606), .B1(G20), .B2(new_n514), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n541), .A2(G20), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT22), .B1(new_n294), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT24), .ZN(new_n611));
  AND2_X1   g0411(.A1(KEYINPUT22), .A2(G87), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n372), .A2(new_n264), .A3(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n610), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n254), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n466), .A2(new_n468), .A3(G107), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n246), .A2(new_n217), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT25), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n566), .A2(new_n275), .A3(G264), .A4(new_n277), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n491), .A2(new_n622), .ZN(new_n623));
  MUX2_X1   g0423(.A(G250), .B(G257), .S(G1698), .Z(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n366), .A3(new_n288), .ZN(new_n625));
  NAND2_X1  g0425(.A1(G33), .A2(G294), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n300), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT93), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n405), .B1(new_n625), .B2(new_n626), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT93), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n311), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n631), .A2(new_n623), .A3(new_n413), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n621), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n617), .A2(new_n620), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n616), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n630), .A2(new_n322), .A3(new_n632), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n324), .B1(new_n631), .B2(new_n623), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n585), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT90), .B1(new_n572), .B2(new_n581), .ZN(new_n644));
  OAI21_X1  g0444(.A(G190), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n584), .A2(G200), .A3(new_n585), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n587), .A2(new_n597), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n582), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n647), .A3(G179), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n603), .A2(new_n642), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n328), .A2(new_n453), .A3(new_n563), .A4(new_n652), .ZN(G372));
  NAND2_X1  g0453(.A1(new_n359), .A2(new_n360), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n423), .A2(new_n427), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n326), .A2(new_n452), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n321), .B2(new_n657), .ZN(new_n658));
  AOI221_X4 g0458(.A(KEYINPUT18), .B1(new_n412), .B2(new_n414), .C1(new_n389), .C2(new_n402), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n416), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n654), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n355), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n453), .A2(new_n328), .ZN(new_n665));
  INV_X1    g0465(.A(new_n561), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n562), .A2(KEYINPUT26), .A3(new_n508), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n508), .A2(new_n554), .A3(new_n561), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT94), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n633), .A2(new_n634), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n637), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n621), .B(KEYINPUT94), .C1(new_n633), .C2(new_n634), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n676), .A2(new_n603), .A3(new_n651), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n508), .B1(new_n498), .B2(new_n503), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n562), .A3(new_n641), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n671), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n665), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n664), .A2(new_n681), .ZN(G369));
  AND2_X1   g0482(.A1(new_n603), .A2(new_n651), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n244), .A2(new_n264), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(G213), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OR3_X1    g0490(.A1(new_n683), .A2(new_n648), .A3(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n603), .A2(new_n651), .A3(new_n649), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n648), .B2(new_n690), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n642), .B1(new_n637), .B2(new_n690), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n635), .A2(new_n690), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n683), .A2(new_n689), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n702), .A2(new_n642), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n676), .A2(new_n689), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n206), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n540), .A2(new_n541), .A3(new_n595), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n213), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n680), .A2(new_n690), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n603), .A2(new_n635), .A3(new_n651), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n678), .A3(new_n562), .A4(new_n641), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT95), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n668), .A2(new_n720), .A3(new_n669), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n668), .B2(new_n669), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n667), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n723), .A3(new_n561), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n717), .B1(new_n724), .B2(new_n690), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n554), .A2(new_n561), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n508), .B(new_n727), .C1(new_n498), .C2(new_n503), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(new_n692), .A3(new_n642), .A4(new_n690), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n490), .A2(new_n634), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n518), .A2(new_n532), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n650), .A3(KEYINPUT30), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n413), .B1(new_n631), .B2(new_n623), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n535), .B2(new_n536), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n584), .A2(new_n735), .A3(new_n495), .A4(new_n585), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n535), .A2(new_n572), .A3(new_n536), .A4(new_n581), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n738), .B2(new_n730), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n733), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n689), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n726), .B1(new_n729), .B2(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n716), .A2(new_n725), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT96), .Z(new_n749));
  OAI21_X1  g0549(.A(new_n714), .B1(new_n749), .B2(G1), .ZN(G364));
  XNOR2_X1  g0550(.A(new_n695), .B(KEYINPUT97), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n264), .A2(G13), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n244), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n708), .ZN(new_n756));
  INV_X1    g0556(.A(new_n694), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(new_n726), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n264), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT103), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n294), .A2(new_n206), .ZN(new_n765));
  INV_X1    g0565(.A(G355), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n766), .B1(G116), .B2(new_n206), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n239), .A2(new_n529), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n372), .A2(new_n707), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n213), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n529), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n767), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n209), .B1(G20), .B2(new_n311), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n761), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n756), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n264), .A2(new_n413), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT99), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n322), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G58), .A2(new_n783), .B1(new_n786), .B2(G77), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n778), .A2(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G190), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n322), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n789), .A2(G68), .B1(new_n790), .B2(G50), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n264), .A2(G179), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n784), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n377), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n264), .B1(new_n781), .B2(new_n413), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n796), .A2(new_n456), .B1(new_n797), .B2(new_n541), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n792), .A2(new_n322), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n217), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n798), .A2(new_n431), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n787), .A2(new_n791), .A3(new_n795), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n785), .A2(new_n803), .B1(new_n804), .B2(new_n796), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n790), .B(KEYINPUT100), .Z(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(new_n807), .B2(G326), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT101), .ZN(new_n809));
  INV_X1    g0609(.A(new_n793), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n294), .B1(new_n810), .B2(G329), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  INV_X1    g0612(.A(new_n789), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT33), .B(G317), .Z(new_n814));
  OAI221_X1 g0614(.A(new_n811), .B1(new_n812), .B2(new_n799), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n783), .B2(G322), .ZN(new_n816));
  INV_X1    g0616(.A(G303), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n797), .B(KEYINPUT102), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n816), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n802), .B1(new_n809), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n777), .B1(new_n821), .B2(new_n774), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n752), .A2(new_n758), .B1(new_n764), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  NOR2_X1   g0624(.A1(new_n452), .A2(new_n689), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n449), .B1(new_n448), .B2(new_n690), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(new_n826), .B2(new_n452), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n715), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n680), .A2(new_n690), .A3(new_n827), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n747), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n756), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n829), .A2(new_n747), .A3(new_n830), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n759), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n775), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n756), .B1(new_n836), .B2(G77), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT104), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n789), .A2(G150), .B1(new_n790), .B2(G137), .ZN(new_n839));
  INV_X1    g0639(.A(G143), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n785), .B2(new_n377), .C1(new_n840), .C2(new_n782), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT34), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n796), .A2(new_n215), .B1(new_n799), .B2(new_n247), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n372), .B1(new_n844), .B2(new_n793), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n843), .B(new_n845), .C1(G50), .C2(new_n818), .ZN(new_n846));
  INV_X1    g0646(.A(new_n796), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(G97), .B1(new_n810), .B2(G311), .ZN(new_n848));
  INV_X1    g0648(.A(new_n790), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n541), .B2(new_n799), .C1(new_n817), .C2(new_n849), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n595), .A2(new_n785), .B1(new_n782), .B2(new_n804), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n813), .A2(KEYINPUT105), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n813), .A2(KEYINPUT105), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n850), .B(new_n851), .C1(G283), .C2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n294), .B1(new_n818), .B2(G107), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT106), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n842), .A2(new_n846), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n838), .B1(new_n775), .B2(new_n859), .C1(new_n827), .C2(new_n835), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n834), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G384));
  NOR3_X1   g0662(.A1(new_n652), .A2(new_n563), .A3(new_n689), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT110), .B1(new_n863), .B2(new_n745), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT110), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n729), .A2(new_n746), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n271), .A2(new_n689), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT107), .Z(new_n869));
  NAND3_X1  g0669(.A1(new_n321), .A2(new_n327), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n869), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT76), .B1(new_n317), .B2(new_n319), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n314), .A2(new_n272), .A3(new_n315), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n270), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n871), .B1(new_n874), .B2(new_n326), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n828), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n403), .A2(new_n415), .ZN(new_n878));
  INV_X1    g0678(.A(new_n687), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n403), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n421), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT109), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n394), .A2(new_n396), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n424), .A2(KEYINPUT16), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n425), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n884), .B1(new_n888), .B2(new_n687), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n380), .A2(new_n254), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n424), .A2(KEYINPUT16), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n885), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(KEYINPUT109), .A3(new_n879), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n415), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n889), .A2(new_n893), .A3(new_n421), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n883), .B1(KEYINPUT37), .B2(new_n895), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n655), .A2(new_n660), .B1(new_n889), .B2(new_n893), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n877), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n882), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n889), .A2(new_n893), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n428), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n867), .A2(new_n876), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n412), .A2(new_n414), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n421), .B1(new_n426), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n426), .A2(new_n687), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n911), .A2(new_n882), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n880), .B1(new_n655), .B2(new_n660), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n877), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT111), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n903), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n903), .B2(new_n914), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n918), .A2(KEYINPUT40), .A3(new_n867), .A4(new_n876), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n907), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n867), .A2(new_n665), .ZN(new_n921));
  OAI21_X1  g0721(.A(G330), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n898), .A2(new_n903), .A3(KEYINPUT39), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n896), .A2(new_n897), .A3(new_n877), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n428), .A2(new_n910), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n911), .A2(new_n882), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n924), .B1(new_n929), .B2(KEYINPUT39), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n874), .A2(new_n690), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n930), .A2(new_n931), .B1(new_n660), .B2(new_n879), .ZN(new_n932));
  INV_X1    g0732(.A(new_n825), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n870), .A2(new_n875), .B1(new_n830), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT108), .ZN(new_n936));
  INV_X1    g0736(.A(new_n904), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n935), .B2(KEYINPUT108), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n932), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n665), .B1(new_n716), .B2(new_n725), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n664), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n923), .A2(new_n942), .B1(new_n244), .B2(new_n753), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n942), .B2(new_n923), .ZN(new_n944));
  INV_X1    g0744(.A(new_n459), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n945), .A2(KEYINPUT35), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(KEYINPUT35), .ZN(new_n947));
  NOR4_X1   g0747(.A1(new_n946), .A2(new_n947), .A3(new_n212), .A4(new_n595), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n213), .A2(new_n334), .A3(new_n375), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n259), .A2(G68), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n244), .B(G13), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n944), .A2(new_n949), .A3(new_n952), .ZN(G367));
  AOI21_X1  g0753(.A(new_n776), .B1(new_n707), .B2(new_n445), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n234), .B2(new_n770), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n756), .ZN(new_n956));
  INV_X1    g0756(.A(new_n797), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT46), .B1(new_n957), .B2(G116), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n818), .A2(KEYINPUT46), .A3(G116), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n854), .B2(new_n804), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n372), .B1(G317), .B2(new_n810), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n799), .A2(new_n456), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G107), .B2(new_n847), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n961), .B(new_n963), .C1(new_n806), .C2(new_n803), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n812), .A2(new_n785), .B1(new_n782), .B2(new_n817), .ZN(new_n965));
  OR4_X1    g0765(.A1(new_n958), .A2(new_n960), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n855), .A2(G159), .B1(G50), .B2(new_n786), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT114), .ZN(new_n968));
  INV_X1    g0768(.A(G137), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n294), .B1(new_n793), .B2(new_n969), .C1(new_n796), .C2(new_n247), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n215), .A2(new_n797), .B1(new_n799), .B2(new_n334), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(new_n783), .C2(G150), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n968), .B(new_n972), .C1(new_n840), .C2(new_n806), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n967), .A2(KEYINPUT114), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n966), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n956), .B1(new_n976), .B2(new_n774), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n553), .A2(new_n690), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n727), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n666), .A2(new_n978), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n763), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n678), .B1(new_n471), .B2(new_n690), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n508), .A2(new_n689), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n703), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT112), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n509), .B1(new_n983), .B2(new_n635), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n986), .A2(KEYINPUT42), .B1(new_n690), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n979), .A2(new_n980), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n988), .A2(new_n990), .B1(KEYINPUT43), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n992), .B(new_n993), .Z(new_n994));
  INV_X1    g0794(.A(new_n985), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n701), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n994), .B(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n705), .A2(new_n985), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT44), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n703), .A2(new_n704), .A3(new_n995), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(new_n701), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n702), .A2(new_n698), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n703), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT113), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n695), .B(new_n1006), .C1(KEYINPUT97), .C2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n751), .A2(KEYINPUT113), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n1009), .B2(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n749), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n749), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n708), .B(KEYINPUT41), .Z(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n755), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n982), .B1(new_n998), .B2(new_n1017), .ZN(G387));
  NAND2_X1  g0818(.A1(new_n699), .A2(new_n763), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n765), .A2(new_n711), .B1(G107), .B2(new_n206), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n231), .A2(new_n529), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n346), .A2(G50), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT50), .ZN(new_n1023));
  AOI211_X1 g0823(.A(G45), .B(new_n710), .C1(G68), .C2(G77), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n770), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1020), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n756), .B1(new_n1026), .B2(new_n776), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G50), .A2(new_n783), .B1(new_n786), .B2(G68), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n377), .A2(new_n849), .B1(new_n813), .B2(new_n346), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n797), .A2(new_n334), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1029), .A2(new_n962), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n558), .A2(new_n847), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n372), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G150), .B2(new_n810), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n372), .B1(G326), .B2(new_n810), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n796), .A2(new_n812), .B1(new_n797), .B2(new_n804), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n807), .A2(G322), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G317), .A2(new_n783), .B1(new_n786), .B2(G303), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n803), .C2(new_n854), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1036), .B1(new_n595), .B2(new_n799), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1035), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1027), .B1(new_n1047), .B2(new_n774), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1010), .A2(new_n755), .B1(new_n1019), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1011), .A2(new_n708), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1010), .A2(new_n749), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n1004), .A2(new_n755), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n776), .B1(G97), .B2(new_n707), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n242), .A2(new_n769), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n708), .B(new_n755), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n799), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n847), .A2(G77), .B1(new_n1057), .B2(G87), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n247), .B2(new_n797), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n372), .B1(new_n840), .B2(new_n793), .C1(new_n785), .C2(new_n346), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G50), .C2(new_n855), .ZN(new_n1061));
  INV_X1    g0861(.A(G150), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n782), .A2(new_n377), .B1(new_n1062), .B2(new_n849), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n783), .A2(G311), .B1(G317), .B2(new_n790), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1066));
  XNOR2_X1  g0866(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n294), .B(new_n800), .C1(G322), .C2(new_n810), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n847), .A2(G116), .B1(new_n957), .B2(G283), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n804), .C2(new_n785), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G303), .B2(new_n855), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1061), .A2(new_n1064), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1056), .B1(new_n775), .B2(new_n1072), .C1(new_n985), .C2(new_n761), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1053), .A2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n709), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1075), .A2(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G390));
  NAND2_X1  g0880(.A1(new_n826), .A2(new_n452), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n724), .A2(new_n690), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n933), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n870), .A2(new_n875), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n864), .A2(new_n866), .A3(G330), .A4(new_n827), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AND4_X1   g0887(.A1(KEYINPUT118), .A2(new_n1084), .A3(new_n747), .A4(new_n827), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT118), .B1(new_n876), .B2(new_n747), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(G330), .B(new_n827), .C1(new_n863), .C2(new_n745), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n870), .A3(new_n875), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1084), .A2(new_n827), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n864), .A2(new_n866), .A3(G330), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n830), .A2(new_n933), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n867), .A2(G330), .A3(new_n665), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n664), .A2(new_n940), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n931), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n874), .A2(KEYINPUT117), .A3(new_n690), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1103), .A2(new_n918), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n931), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n930), .B1(new_n934), .B2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1108), .B(new_n1110), .C1(new_n1089), .C2(new_n1088), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1096), .B2(new_n1084), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT39), .B1(new_n903), .B2(new_n914), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n937), .B2(KEYINPUT39), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT111), .B1(new_n925), .B2(new_n928), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n903), .A2(new_n914), .A3(new_n915), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1115), .A2(new_n1116), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1082), .A2(new_n933), .B1(new_n870), .B2(new_n875), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1112), .A2(new_n1114), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1111), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1102), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1098), .A2(new_n1101), .A3(new_n1111), .A4(new_n1121), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n708), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1111), .A2(new_n1121), .A3(new_n755), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n756), .B1(new_n836), .B2(new_n347), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  AOI22_X1  g0928(.A1(new_n855), .A2(G137), .B1(new_n786), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT119), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n783), .A2(G132), .B1(G128), .B2(new_n790), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT120), .Z(new_n1132));
  AOI21_X1  g0932(.A(new_n431), .B1(new_n810), .B2(G125), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n259), .B2(new_n799), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n957), .A2(G150), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G159), .C2(new_n847), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1130), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n854), .A2(new_n217), .B1(new_n456), .B2(new_n785), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT121), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n431), .B1(new_n793), .B2(new_n804), .C1(new_n247), .C2(new_n799), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n849), .A2(new_n812), .B1(new_n334), .B2(new_n796), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n783), .C2(G116), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n541), .B2(new_n819), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1138), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1127), .B1(new_n1145), .B2(new_n774), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1114), .B2(new_n835), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1126), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1148), .A2(KEYINPUT122), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(KEYINPUT122), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1125), .B1(new_n1149), .B2(new_n1150), .ZN(G378));
  XNOR2_X1  g0951(.A(new_n1100), .B(KEYINPUT123), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1124), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n907), .A2(G330), .A3(new_n919), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n353), .A2(new_n879), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n361), .B(new_n1155), .Z(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1158), .A2(G330), .A3(new_n907), .A4(new_n919), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1160), .A2(new_n939), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n939), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1153), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT57), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n709), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1153), .B(KEYINPUT57), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT124), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n939), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1160), .A2(new_n939), .A3(new_n1161), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT124), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(KEYINPUT57), .A4(new_n1153), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1166), .A2(new_n1168), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1159), .A2(new_n759), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n756), .B1(new_n836), .B2(G50), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n796), .A2(new_n247), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n485), .B1(new_n793), .B2(new_n812), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1179), .A2(new_n1180), .A3(new_n1030), .A4(new_n372), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n785), .B2(new_n557), .C1(new_n217), .C2(new_n782), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n799), .A2(new_n215), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n813), .A2(new_n456), .B1(new_n849), .B2(new_n595), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n485), .B1(new_n371), .B2(new_n261), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n259), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G128), .A2(new_n783), .B1(new_n786), .B2(G137), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n790), .A2(G125), .B1(new_n847), .B2(G150), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n789), .A2(G132), .B1(new_n957), .B2(new_n1128), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1057), .A2(G159), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n810), .C2(G124), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1189), .B1(KEYINPUT58), .B2(new_n1185), .C1(new_n1194), .C2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1178), .B1(new_n1199), .B2(new_n774), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1173), .A2(new_n755), .B1(new_n1177), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1176), .A2(new_n1201), .ZN(G375));
  NAND3_X1  g1002(.A1(new_n1090), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1015), .B(KEYINPUT125), .Z(new_n1204));
  NAND3_X1  g1004(.A1(new_n1102), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1085), .A2(new_n759), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n756), .B1(new_n836), .B2(G68), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n855), .A2(new_n1128), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n818), .A2(G159), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n790), .A2(G132), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1183), .B1(G50), .B2(new_n847), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1033), .B1(G128), .B2(new_n810), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n785), .B2(new_n1062), .C1(new_n969), .C2(new_n782), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n799), .A2(new_n334), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n431), .B1(new_n793), .B2(new_n817), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G294), .C2(new_n790), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n456), .B2(new_n819), .C1(new_n854), .C2(new_n595), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1032), .B1(new_n785), .B2(new_n217), .C1(new_n812), .C2(new_n782), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n1212), .A2(new_n1214), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1207), .B1(new_n1220), .B2(new_n774), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1098), .A2(new_n755), .B1(new_n1206), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1205), .A2(new_n1222), .ZN(G381));
  NAND2_X1  g1023(.A1(new_n1079), .A2(new_n861), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1224), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1125), .A2(new_n1148), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(G387), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n1201), .A3(new_n1176), .A4(new_n1227), .ZN(G407));
  INV_X1    g1028(.A(new_n1226), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n688), .A2(G213), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G375), .C2(new_n1232), .ZN(G409));
  XNOR2_X1  g1033(.A(G393), .B(G396), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT127), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G387), .A2(new_n1079), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(new_n1079), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1236), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1239), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(new_n1237), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1234), .B(KEYINPUT127), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT61), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1203), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1090), .A2(new_n1097), .A3(new_n1100), .A4(KEYINPUT60), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n708), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1222), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n861), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(G384), .A3(new_n1222), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1231), .A2(G2897), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1253), .B(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1173), .A2(new_n1153), .A3(new_n1204), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1226), .B1(new_n1201), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1176), .A2(G378), .A3(new_n1201), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1176), .A2(KEYINPUT126), .A3(G378), .A4(new_n1201), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1257), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1255), .B1(new_n1262), .B2(new_n1231), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1262), .A2(new_n1231), .A3(new_n1253), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1245), .B(new_n1263), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1257), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1253), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1230), .A3(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT62), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1244), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1263), .A2(new_n1245), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1235), .B1(new_n1241), .B2(new_n1237), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1264), .A2(KEYINPUT63), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1274), .A2(new_n1276), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1273), .A2(new_n1281), .ZN(G405));
  NAND2_X1  g1082(.A1(G375), .A2(new_n1229), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1267), .A2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1253), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1279), .ZN(G402));
endmodule


