//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226,
    new_n1227, new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(KEYINPUT68), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(KEYINPUT68), .B2(new_n459), .ZN(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(KEYINPUT69), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n473), .C1(new_n466), .C2(new_n467), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(G101), .A3(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT70), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n466), .A2(new_n467), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n483), .B2(new_n473), .ZN(new_n489));
  OAI211_X1 g064(.A(KEYINPUT72), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  OR2_X1    g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n487), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n496), .A2(KEYINPUT73), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(KEYINPUT73), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n464), .A2(new_n468), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(G138), .B(new_n473), .C1(new_n466), .C2(new_n467), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT74), .B(G114), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT75), .B1(new_n511), .B2(G2105), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT74), .A2(G114), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT74), .A2(G114), .ZN(new_n514));
  OAI211_X1 g089(.A(KEYINPUT75), .B(G2105), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n510), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  OAI211_X1 g104(.A(G50), .B(G543), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  AND2_X1   g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n532), .B1(new_n528), .B2(new_n529), .ZN(new_n533));
  INV_X1    g108(.A(G88), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g112(.A(KEYINPUT76), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n527), .B1(new_n537), .B2(new_n538), .ZN(G166));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT77), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT7), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  OR2_X1    g118(.A1(KEYINPUT6), .A2(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(KEYINPUT6), .A2(G651), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n521), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G51), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n548));
  INV_X1    g123(.A(G89), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n533), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n543), .A2(new_n550), .ZN(G168));
  AOI22_X1  g126(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n526), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI21_X1  g129(.A(G543), .B1(new_n528), .B2(new_n529), .ZN(new_n555));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n533), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(G171));
  AOI22_X1  g133(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n526), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  INV_X1    g136(.A(G43), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n533), .A2(new_n561), .B1(new_n555), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n546), .A2(G53), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n524), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n573), .A2(new_n526), .B1(new_n574), .B2(new_n533), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  NAND2_X1  g154(.A1(new_n537), .A2(new_n538), .ZN(new_n580));
  INV_X1    g155(.A(new_n527), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G303));
  NAND2_X1  g157(.A1(new_n546), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n533), .ZN(G288));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n522), .B2(new_n523), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT78), .B(G651), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n544), .A2(new_n545), .B1(new_n522), .B2(new_n523), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G86), .B1(new_n546), .B2(G48), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n594), .A2(G85), .B1(new_n546), .B2(G47), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n526), .B2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n546), .A2(G54), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n524), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n526), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT79), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n594), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT10), .Z(new_n606));
  AND2_X1   g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n600), .B1(new_n607), .B2(G868), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G286), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n576), .B(KEYINPUT80), .Z(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n610), .ZN(G297));
  AOI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n610), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G860), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT81), .Z(G148));
  NAND2_X1  g192(.A1(new_n607), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND4_X1  g196(.A1(new_n464), .A2(new_n468), .A3(G2104), .A4(new_n473), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT13), .Z(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n492), .A2(G123), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(KEYINPUT82), .ZN(new_n630));
  INV_X1    g205(.A(G111), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n629), .A2(KEYINPUT82), .B1(new_n631), .B2(G2105), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n484), .A2(G135), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n626), .A2(new_n627), .A3(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n641), .B(new_n647), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n625), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n635), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  MUX2_X1   g250(.A(new_n675), .B(new_n674), .S(new_n667), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(G229));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n497), .B2(new_n498), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(G35), .ZN(new_n692));
  OR3_X1    g267(.A1(new_n691), .A2(KEYINPUT29), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G2090), .ZN(new_n694));
  OAI21_X1  g269(.A(KEYINPUT29), .B1(new_n691), .B2(new_n692), .ZN(new_n695));
  AND3_X1   g270(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n690), .A2(G32), .ZN(new_n699));
  INV_X1    g274(.A(G129), .ZN(new_n700));
  OR3_X1    g275(.A1(new_n491), .A2(KEYINPUT91), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(KEYINPUT91), .B1(new_n491), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g278(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT26), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n704), .B(new_n706), .C1(G141), .C2(new_n484), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n699), .B1(new_n709), .B2(new_n690), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(KEYINPUT92), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(KEYINPUT92), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n634), .A2(new_n690), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT94), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n564), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G16), .B2(G19), .ZN(new_n719));
  INV_X1    g294(.A(G1341), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT93), .ZN(new_n723));
  INV_X1    g298(.A(G28), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n724), .B2(KEYINPUT30), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(KEYINPUT30), .B2(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n721), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n717), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(G286), .A2(G16), .ZN(new_n729));
  INV_X1    g304(.A(G21), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(G16), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G1966), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n729), .B(G1966), .C1(G16), .C2(new_n730), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  NAND2_X1  g310(.A1(G164), .A2(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G27), .B2(G29), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n481), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT90), .B(G2084), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n746), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1961), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n719), .A2(new_n720), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n728), .A2(new_n738), .A3(new_n745), .A4(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n713), .B1(new_n711), .B2(new_n714), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n690), .A2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n484), .A2(G139), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n464), .A2(new_n468), .A3(G127), .ZN(new_n760));
  NAND2_X1  g335(.A1(G115), .A2(G2104), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n756), .B(new_n759), .C1(new_n762), .C2(new_n473), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT89), .Z(new_n764));
  OAI21_X1  g339(.A(new_n755), .B1(new_n764), .B2(new_n690), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G2072), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n746), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n576), .B2(new_n746), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n737), .A2(new_n735), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2072), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(new_n755), .C1(new_n764), .C2(new_n690), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n690), .A2(G26), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT28), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n492), .A2(G128), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(G116), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(G2105), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n484), .B2(G140), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2067), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n766), .A2(new_n772), .A3(new_n774), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n604), .A2(new_n606), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n746), .A2(G4), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT88), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(KEYINPUT88), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G1348), .ZN(new_n793));
  INV_X1    g368(.A(G1348), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n790), .A2(new_n794), .A3(new_n791), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n785), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n698), .A2(new_n715), .A3(new_n754), .A4(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(G6), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G305), .B2(new_n746), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1981), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n746), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n746), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1971), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT87), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G23), .ZN(new_n806));
  XNOR2_X1  g381(.A(G288), .B(KEYINPUT86), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n806), .B1(new_n808), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT33), .B(G1976), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n804), .A2(KEYINPUT87), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n801), .A2(new_n805), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n815));
  NOR2_X1   g390(.A1(G25), .A2(G29), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n484), .A2(G131), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT84), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n492), .A2(G119), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n816), .B1(new_n823), .B2(G29), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n824), .A2(new_n826), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n746), .A2(G24), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT85), .Z(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G290), .B2(G16), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(G1986), .Z(new_n832));
  NOR3_X1   g407(.A1(new_n827), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n814), .A2(new_n815), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n814), .A2(new_n815), .A3(new_n836), .A4(new_n833), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n797), .B1(new_n835), .B2(new_n837), .ZN(G311));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n839));
  XNOR2_X1  g414(.A(G311), .B(new_n839), .ZN(G150));
  AOI22_X1  g415(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n526), .ZN(new_n842));
  INV_X1    g417(.A(G93), .ZN(new_n843));
  INV_X1    g418(.A(G55), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n533), .A2(new_n843), .B1(new_n555), .B2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(KEYINPUT96), .ZN(new_n850));
  OR3_X1    g425(.A1(new_n842), .A2(KEYINPUT96), .A3(new_n845), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n564), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n846), .B(KEYINPUT96), .C1(new_n560), .C2(new_n563), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n607), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT97), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n857), .B2(new_n858), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n849), .B1(new_n863), .B2(new_n864), .ZN(G145));
  NAND2_X1  g440(.A1(new_n709), .A2(new_n782), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n518), .A2(KEYINPUT100), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n508), .A2(new_n517), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n782), .B1(new_n703), .B2(new_n707), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n866), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n782), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n708), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n870), .B1(new_n876), .B2(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n763), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n877), .A3(new_n764), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(KEYINPUT101), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n880), .A2(KEYINPUT101), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n489), .A2(G130), .A3(new_n490), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT102), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(KEYINPUT102), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  INV_X1    g464(.A(G118), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(G2105), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n484), .ZN(new_n893));
  INV_X1    g468(.A(G142), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n887), .A2(new_n888), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n888), .B1(new_n887), .B2(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n623), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(new_n623), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n823), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n883), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n904), .B(new_n822), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n881), .A3(new_n882), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(G162), .A2(new_n481), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n499), .A2(G160), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n910), .A2(new_n634), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n634), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n907), .A2(KEYINPUT104), .A3(new_n881), .A4(new_n882), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n906), .A4(new_n914), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(KEYINPUT40), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT40), .B1(new_n916), .B2(new_n920), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G395));
  XNOR2_X1  g498(.A(G303), .B(KEYINPUT107), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(G305), .ZN(new_n925));
  XNOR2_X1  g500(.A(G166), .B(KEYINPUT107), .ZN(new_n926));
  OAI211_X1 g501(.A(G48), .B(G543), .C1(new_n528), .C2(new_n529), .ZN(new_n927));
  INV_X1    g502(.A(G86), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n533), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n591), .B2(new_n590), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n593), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n807), .B(G290), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n925), .A2(new_n933), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(KEYINPUT108), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n937), .A2(KEYINPUT42), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(KEYINPUT109), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n618), .B(KEYINPUT105), .ZN(new_n946));
  INV_X1    g521(.A(new_n854), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n618), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n854), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n607), .A2(new_n576), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n786), .A2(G299), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(KEYINPUT41), .ZN(new_n958));
  XNOR2_X1  g533(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n953), .B2(new_n954), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n957), .B1(new_n952), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n939), .B2(new_n940), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n965), .B2(new_n943), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n945), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n962), .B1(new_n966), .B2(new_n945), .ZN(new_n968));
  OAI21_X1  g543(.A(G868), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n846), .A2(new_n610), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(G295));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n970), .ZN(G331));
  XNOR2_X1  g547(.A(G168), .B(G171), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n854), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n854), .A2(new_n973), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n956), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n955), .A2(KEYINPUT41), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n953), .A2(new_n954), .A3(new_n959), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n975), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n953), .A2(KEYINPUT110), .A3(new_n954), .A4(new_n959), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n976), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(new_n940), .A3(new_n939), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n981), .B1(new_n958), .B2(new_n960), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n976), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G37), .B1(new_n941), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n984), .A2(KEYINPUT111), .A3(new_n940), .A4(new_n939), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n987), .A2(new_n991), .A3(new_n992), .A4(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n941), .A2(new_n990), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(new_n939), .A3(new_n940), .ZN(new_n995));
  INV_X1    g570(.A(G37), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT44), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n987), .A2(new_n991), .A3(new_n992), .A4(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1001), .A2(new_n1006), .ZN(G397));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n592), .A2(new_n1008), .A3(new_n595), .A4(new_n593), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT116), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n930), .A2(new_n1011), .A3(new_n1008), .A4(new_n593), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(G305), .B2(G1981), .ZN(new_n1019));
  AND3_X1   g594(.A1(G305), .A2(new_n1018), .A3(G1981), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1014), .B(new_n1017), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n474), .A2(new_n478), .A3(new_n475), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n478), .B1(new_n474), .B2(new_n475), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n473), .B1(new_n469), .B2(new_n470), .ZN(new_n1026));
  INV_X1    g601(.A(G40), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n508), .B2(new_n517), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1022), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1021), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1019), .ZN(new_n1032));
  NAND3_X1  g607(.A1(G305), .A2(new_n1018), .A3(G1981), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1017), .B1(new_n1034), .B2(new_n1014), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT119), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1020), .A2(new_n1019), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1015), .B(new_n1016), .C1(new_n1037), .C2(new_n1013), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1030), .A4(new_n1021), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G288), .A2(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1013), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1030), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n807), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT52), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1030), .B(new_n1048), .C1(new_n1045), .C2(new_n807), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G1384), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n867), .A2(new_n869), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1384), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n518), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1053), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1058), .A3(new_n1028), .ZN(new_n1059));
  INV_X1    g634(.A(G1971), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1057), .A2(KEYINPUT50), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n472), .A2(new_n480), .A3(G40), .ZN(new_n1063));
  NOR2_X1   g638(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n508), .B2(new_n517), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1061), .B1(G2090), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G166), .A2(new_n1022), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT115), .B1(new_n1070), .B2(KEYINPUT55), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1072), .B(new_n1073), .C1(G166), .C2(new_n1022), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT114), .B1(new_n1070), .B2(KEYINPUT55), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n1076));
  NOR4_X1   g651(.A1(G166), .A2(new_n1076), .A3(new_n1073), .A4(new_n1022), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1071), .B(new_n1074), .C1(new_n1075), .C2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1069), .A2(G8), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1043), .A2(new_n1044), .B1(new_n1052), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1050), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n518), .A2(new_n1064), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1028), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n518), .B2(new_n1056), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1060), .A2(new_n1059), .B1(new_n1087), .B2(new_n694), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1082), .B1(new_n1088), .B2(new_n1022), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1041), .A2(new_n1081), .A3(new_n1079), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1054), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n508), .B2(new_n517), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1063), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1966), .B1(new_n1058), .B2(new_n1093), .ZN(new_n1094));
  NOR4_X1   g669(.A1(new_n1086), .A2(new_n1063), .A3(G2084), .A4(new_n1066), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1096), .A2(G286), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT120), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT63), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT63), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT120), .B(new_n1100), .C1(new_n1090), .C2(new_n1097), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1080), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT125), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n518), .A2(new_n1054), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1028), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1029), .A2(KEYINPUT45), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n732), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n1108));
  INV_X1    g683(.A(G2084), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1062), .A2(new_n1067), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(G286), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(new_n1022), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT126), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1108), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1118));
  OAI21_X1  g693(.A(G168), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1114), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1096), .B(new_n1113), .C1(new_n1022), .C2(G168), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1116), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G168), .A2(new_n1022), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1103), .A2(new_n1124), .A3(new_n1111), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT62), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(new_n1128), .A3(new_n1125), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1059), .B2(G2078), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT127), .B(G1961), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n1068), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1130), .A2(G2078), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1058), .A2(new_n1093), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1090), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1127), .A2(new_n1129), .A3(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1055), .A2(new_n1058), .A3(new_n1028), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1956), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n576), .B(KEYINPUT57), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1141), .A2(new_n1145), .A3(new_n1143), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT61), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1028), .A2(new_n1151), .A3(new_n1029), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT58), .B(G1341), .ZN(new_n1154));
  OAI22_X1  g729(.A1(G1996), .A2(new_n1059), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n564), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1158), .A3(new_n564), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1149), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1144), .A2(new_n1162), .A3(new_n1146), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1161), .A2(KEYINPUT61), .A3(new_n1148), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(G2067), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1166), .A2(new_n1167), .B1(new_n794), .B2(new_n1068), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1153), .A2(KEYINPUT122), .A3(new_n1165), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(KEYINPUT60), .A3(new_n607), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1168), .A2(new_n1169), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1160), .A2(new_n1164), .A3(new_n1171), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n786), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1148), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g755(.A(KEYINPUT124), .B(new_n1148), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1175), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT45), .B1(new_n871), .B2(new_n1056), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1055), .A2(new_n1028), .A3(new_n1134), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(G171), .B(KEYINPUT54), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1133), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1186), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1188), .A2(new_n1131), .B1(new_n1136), .B2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1190), .A2(new_n1051), .A3(new_n1079), .A4(new_n1089), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1125), .B2(new_n1123), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1182), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1102), .A2(new_n1139), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1183), .A2(new_n1028), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(G290), .A2(G1986), .ZN(new_n1197));
  AND2_X1   g772(.A1(G290), .A2(G1986), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n782), .B(new_n1165), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT112), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1201), .A2(new_n1195), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT113), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n823), .A2(new_n825), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n822), .A2(new_n826), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1196), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n708), .B(G1996), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1196), .A2(new_n1207), .ZN(new_n1208));
  AND4_X1   g783(.A1(new_n1199), .A2(new_n1203), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1194), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1203), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n875), .A2(new_n1165), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1195), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1195), .B1(new_n1201), .B2(new_n709), .ZN(new_n1214));
  OAI21_X1  g789(.A(KEYINPUT46), .B1(new_n1195), .B2(G1996), .ZN(new_n1215));
  OR3_X1    g790(.A1(new_n1195), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT47), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT48), .ZN(new_n1220));
  AND4_X1   g795(.A1(new_n1206), .A2(new_n1203), .A3(new_n1208), .A4(new_n1220), .ZN(new_n1221));
  NOR3_X1   g796(.A1(new_n1213), .A2(new_n1218), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1210), .A2(new_n1222), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g798(.A1(new_n916), .A2(new_n920), .ZN(new_n1225));
  INV_X1    g799(.A(G227), .ZN(new_n1226));
  OAI211_X1 g800(.A(G319), .B(new_n1226), .C1(new_n652), .C2(new_n651), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n685), .B2(new_n688), .ZN(new_n1228));
  AND3_X1   g802(.A1(new_n1225), .A2(new_n1004), .A3(new_n1228), .ZN(G308));
  NAND3_X1  g803(.A1(new_n1225), .A2(new_n1004), .A3(new_n1228), .ZN(G225));
endmodule


