//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n457), .A2(G2106), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(KEYINPUT67), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(G567), .B2(new_n459), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G137), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AND3_X1   g047(.A1(new_n472), .A2(KEYINPUT69), .A3(G101), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT69), .B1(new_n472), .B2(G101), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g050(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(G125), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n469), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n475), .A2(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g060(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT71), .Z(new_n488));
  NOR2_X1   g063(.A1(new_n479), .A2(new_n480), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(new_n469), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(G124), .A2(new_n490), .B1(new_n491), .B2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT72), .ZN(G162));
  OAI211_X1 g069(.A(G138), .B(new_n469), .C1(new_n479), .C2(new_n480), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .A4(new_n469), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT73), .A2(G114), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT73), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n497), .A2(new_n498), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n516), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT74), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n520), .A2(G543), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n520), .A2(new_n521), .A3(new_n512), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n515), .A2(new_n523), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n522), .A2(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n512), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n514), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n522), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n524), .A2(G90), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n514), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n522), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n524), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND4_X1  g128(.A1(new_n520), .A2(G53), .A3(G543), .A4(new_n521), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n512), .A2(G65), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n514), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(G91), .B2(new_n524), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G299));
  NAND2_X1  g135(.A1(new_n522), .A2(G49), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n524), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n510), .B2(new_n511), .ZN(new_n566));
  AND2_X1   g141(.A1(G73), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n521), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n520), .A2(G86), .A3(new_n521), .A4(new_n512), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G305));
  XOR2_X1   g146(.A(KEYINPUT75), .B(G85), .Z(new_n572));
  AOI22_X1  g147(.A1(G47), .A2(new_n522), .B1(new_n524), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT76), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n514), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G290));
  INV_X1    g152(.A(G868), .ZN(new_n578));
  NOR2_X1   g153(.A1(G301), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G54), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n520), .A2(G543), .A3(new_n521), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(KEYINPUT77), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n582), .B1(KEYINPUT77), .B2(new_n581), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n520), .A2(new_n521), .A3(new_n512), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n514), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n583), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n579), .B1(new_n594), .B2(new_n578), .ZN(G284));
  AOI21_X1  g170(.A(new_n579), .B1(new_n594), .B2(new_n578), .ZN(G321));
  NAND2_X1  g171(.A1(G299), .A2(new_n578), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n578), .B2(G168), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n578), .B2(G168), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n594), .B1(new_n600), .B2(G860), .ZN(G148));
  NOR2_X1   g176(.A1(new_n548), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n594), .A2(new_n600), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n468), .A2(new_n472), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n491), .A2(G135), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n490), .A2(G123), .ZN(new_n614));
  OR2_X1    g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n615), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND3_X1  g193(.A1(new_n611), .A2(new_n612), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n628), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT82), .ZN(new_n636));
  OAI21_X1  g211(.A(G14), .B1(new_n632), .B2(new_n634), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT83), .ZN(new_n641));
  NOR2_X1   g216(.A1(G2072), .A2(G2078), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n444), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(KEYINPUT17), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT84), .Z(new_n647));
  OAI211_X1 g222(.A(new_n639), .B(new_n640), .C1(new_n444), .C2(new_n642), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n641), .A2(new_n639), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n649), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n658), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  MUX2_X1   g239(.A(new_n664), .B(new_n663), .S(new_n656), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G22), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G166), .B2(new_n673), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(G1971), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(G1971), .ZN(new_n678));
  MUX2_X1   g253(.A(G6), .B(G305), .S(G16), .Z(new_n679));
  XOR2_X1   g254(.A(KEYINPUT32), .B(G1981), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(G23), .ZN(new_n682));
  INV_X1    g257(.A(G288), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n673), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT33), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n677), .A2(new_n678), .A3(new_n681), .A4(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G25), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n491), .A2(G131), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n490), .A2(G119), .ZN(new_n693));
  OR2_X1    g268(.A1(G95), .A2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n694), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n691), .B1(new_n697), .B2(new_n690), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n673), .A2(G24), .ZN(new_n701));
  INV_X1    g276(.A(G290), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(KEYINPUT85), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(G16), .B1(new_n702), .B2(KEYINPUT85), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(G1986), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G1986), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n689), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT36), .ZN(new_n710));
  NAND2_X1  g285(.A1(G160), .A2(G29), .ZN(new_n711));
  INV_X1    g286(.A(G34), .ZN(new_n712));
  AOI21_X1  g287(.A(G29), .B1(new_n712), .B2(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(KEYINPUT24), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G2084), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n673), .A2(G5), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G171), .B2(new_n673), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT94), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n690), .A2(G32), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n491), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n490), .A2(G129), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n721), .B1(new_n731), .B2(new_n690), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT92), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n717), .B1(G1961), .B2(new_n720), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G29), .A2(G35), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G162), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT29), .B(G2090), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n733), .A2(new_n734), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n690), .A2(KEYINPUT28), .A3(G26), .ZN(new_n743));
  AOI21_X1  g318(.A(KEYINPUT28), .B1(new_n690), .B2(G26), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G116), .B2(new_n469), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT87), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n491), .A2(G140), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n490), .A2(G128), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n743), .B(new_n744), .C1(new_n753), .C2(G29), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT88), .B(G2067), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  INV_X1    g333(.A(G28), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT30), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(KEYINPUT30), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n756), .B(new_n762), .C1(new_n690), .C2(new_n617), .ZN(new_n763));
  NOR2_X1   g338(.A1(G168), .A2(new_n673), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n673), .B2(G21), .ZN(new_n765));
  INV_X1    g340(.A(G1966), .ZN(new_n766));
  NOR2_X1   g341(.A1(G27), .A2(G29), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G164), .B2(G29), .ZN(new_n768));
  OAI22_X1  g343(.A1(new_n765), .A2(new_n766), .B1(new_n768), .B2(G2078), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n715), .A2(new_n716), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT90), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n754), .A2(new_n755), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n763), .A2(new_n769), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n737), .A2(new_n741), .A3(new_n742), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(G115), .A2(G2104), .ZN(new_n775));
  INV_X1    g350(.A(G127), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n489), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n469), .B1(new_n777), .B2(KEYINPUT89), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(KEYINPUT89), .B2(new_n777), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT25), .ZN(new_n780));
  NAND2_X1  g355(.A1(G103), .A2(G2104), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(G2105), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n469), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n491), .A2(G139), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G33), .B(new_n785), .S(G29), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(new_n442), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n673), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n548), .B2(new_n673), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1341), .Z(new_n790));
  AOI22_X1  g365(.A1(new_n765), .A2(new_n766), .B1(new_n768), .B2(G2078), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n787), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G1961), .B2(new_n720), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n673), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n594), .B2(new_n673), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G1348), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(G1348), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n793), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n673), .A2(G20), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT23), .Z(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G299), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1956), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n735), .B2(new_n736), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n774), .A2(new_n798), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n710), .A2(new_n805), .ZN(G311));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n807));
  XNOR2_X1  g382(.A(G311), .B(new_n807), .ZN(G150));
  NAND2_X1  g383(.A1(new_n594), .A2(G559), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n522), .A2(G55), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT98), .B(G93), .Z(new_n813));
  OAI221_X1 g388(.A(new_n811), .B1(new_n514), .B2(new_n812), .C1(new_n586), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(new_n547), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n810), .B(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT39), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(KEYINPUT39), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n818), .A2(new_n819), .A3(G860), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n814), .A2(G860), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n820), .A2(new_n822), .ZN(G145));
  NAND2_X1  g398(.A1(new_n491), .A2(G142), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n827));
  INV_X1    g402(.A(G118), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(G2105), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n490), .B2(G130), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n608), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n753), .B(new_n785), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n730), .B(G164), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n696), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(G162), .B(new_n617), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G160), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT101), .B(G37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g420(.A1(new_n814), .A2(new_n578), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n592), .B(G299), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT41), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n603), .B(new_n815), .ZN(new_n849));
  MUX2_X1   g424(.A(new_n848), .B(new_n847), .S(new_n849), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT42), .ZN(new_n851));
  XNOR2_X1  g426(.A(G290), .B(G305), .ZN(new_n852));
  XNOR2_X1  g427(.A(G303), .B(G288), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n851), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n846), .B1(new_n856), .B2(new_n578), .ZN(G295));
  OAI21_X1  g432(.A(new_n846), .B1(new_n856), .B2(new_n578), .ZN(G331));
  XNOR2_X1  g433(.A(new_n815), .B(G301), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n859), .A2(G168), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(G168), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n848), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n847), .B1(new_n860), .B2(new_n861), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n863), .A2(new_n854), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n854), .B1(new_n863), .B2(new_n864), .ZN(new_n866));
  OAI211_X1 g441(.A(KEYINPUT43), .B(new_n843), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n864), .ZN(new_n868));
  INV_X1    g443(.A(new_n854), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n863), .A2(new_n854), .A3(new_n864), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n867), .B1(new_n872), .B2(KEYINPUT43), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT44), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(new_n843), .C1(new_n865), .C2(new_n866), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n872), .B2(new_n875), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n874), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n874), .B2(new_n879), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(G397));
  INV_X1    g458(.A(G1384), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n506), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT45), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n482), .ZN(new_n888));
  INV_X1    g463(.A(new_n474), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n472), .A2(KEYINPUT69), .A3(G101), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n888), .A2(G40), .A3(new_n891), .A4(new_n470), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G1996), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n730), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n752), .B(G2067), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n697), .A2(new_n699), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n697), .A2(new_n699), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(G1986), .B2(G290), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G1986), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n702), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT104), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n893), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n506), .A2(KEYINPUT105), .A3(new_n884), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT105), .B1(new_n506), .B2(new_n884), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n907), .A2(new_n908), .A3(new_n892), .ZN(new_n909));
  INV_X1    g484(.A(G8), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT113), .Z(new_n912));
  INV_X1    g487(.A(G1981), .ZN(new_n913));
  INV_X1    g488(.A(new_n568), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n569), .A2(new_n570), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT108), .ZN(new_n918));
  AOI211_X1 g493(.A(KEYINPUT109), .B(new_n913), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n913), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT109), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n915), .A2(new_n916), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n568), .A3(new_n918), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(G1981), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT110), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT49), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n927), .A3(G1981), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n928), .B(new_n929), .C1(new_n930), .C2(new_n921), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(new_n926), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n928), .B1(new_n930), .B2(new_n921), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT49), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n933), .B2(KEYINPUT49), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n932), .B(new_n911), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(G288), .A2(G1976), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT114), .Z(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n920), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n912), .B1(new_n941), .B2(KEYINPUT115), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT115), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n943), .A3(new_n920), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n683), .A2(G1976), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n885), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G40), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n475), .A2(new_n482), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n506), .A2(KEYINPUT105), .A3(new_n884), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n951), .A3(G8), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n683), .A2(G1976), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n952), .A2(KEYINPUT52), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(KEYINPUT52), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n937), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n937), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n884), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n961), .A2(new_n949), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n887), .ZN(new_n963));
  INV_X1    g538(.A(G1971), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n947), .A2(new_n966), .A3(new_n950), .ZN(new_n967));
  INV_X1    g542(.A(G2090), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n892), .B1(KEYINPUT50), .B2(new_n885), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n910), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  NAND2_X1  g547(.A1(G303), .A2(G8), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT106), .B(KEYINPUT55), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n971), .B2(new_n975), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n942), .A2(new_n944), .B1(new_n960), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n949), .B1(new_n885), .B2(KEYINPUT50), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n947), .A2(new_n950), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(KEYINPUT50), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n968), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n965), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G8), .ZN(new_n986));
  INV_X1    g561(.A(new_n975), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n977), .B2(new_n978), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n956), .A2(KEYINPUT116), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n937), .A2(new_n955), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n967), .A2(new_n716), .A3(new_n969), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n886), .B1(new_n907), .B2(new_n908), .ZN(new_n996));
  AOI21_X1  g571(.A(G1966), .B1(new_n996), .B2(new_n962), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n998), .A2(new_n910), .A3(G286), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT63), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(KEYINPUT63), .ZN(new_n1001));
  INV_X1    g576(.A(new_n971), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(new_n987), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n960), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n980), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT62), .ZN(new_n1007));
  OAI21_X1  g582(.A(G286), .B1(new_n995), .B2(new_n997), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n961), .A2(new_n949), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n982), .B2(new_n886), .ZN(new_n1010));
  OAI211_X1 g585(.A(G168), .B(new_n994), .C1(new_n1010), .C2(G1966), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1008), .A2(KEYINPUT51), .A3(new_n1011), .A4(G8), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(G8), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT123), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1007), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT123), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(KEYINPUT62), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n963), .B2(G2078), .ZN(new_n1025));
  INV_X1    g600(.A(G1961), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT50), .ZN(new_n1027));
  INV_X1    g602(.A(new_n885), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n949), .B1(new_n1028), .B2(new_n966), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1032));
  AOI21_X1  g607(.A(G301), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1019), .A2(new_n1023), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1956), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n966), .B1(new_n947), .B2(new_n950), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n981), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n555), .B2(new_n559), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1042), .B(new_n442), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n887), .A2(new_n949), .A3(new_n961), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT119), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n962), .A2(new_n1046), .A3(new_n887), .A4(new_n1043), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1037), .A2(new_n1041), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1045), .B(new_n1047), .C1(new_n983), .C2(G1956), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1041), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1051), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2067), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n909), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1348), .B1(new_n967), .B2(new_n969), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n594), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1049), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n506), .B2(new_n884), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1009), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT58), .B(G1341), .Z(new_n1066));
  AOI22_X1  g641(.A1(new_n1065), .A2(new_n894), .B1(new_n951), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1063), .B1(new_n1067), .B2(new_n547), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1066), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n963), .A2(G1996), .B1(new_n909), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT59), .A3(new_n548), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n1073));
  INV_X1    g648(.A(G1348), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1075), .B2(new_n1058), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1061), .B1(new_n1076), .B2(new_n594), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1072), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT120), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1048), .A2(KEYINPUT61), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1053), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1061), .B(new_n1078), .C1(new_n1076), .C2(new_n594), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1080), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1048), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT121), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1091), .A3(new_n1088), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1062), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1031), .A2(G301), .A3(new_n1032), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1065), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1025), .A2(new_n1030), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1098), .A2(KEYINPUT125), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(KEYINPUT125), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT54), .B(new_n1095), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1097), .A2(G171), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n1033), .B2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1101), .A2(new_n1021), .A3(new_n1022), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1034), .B1(new_n1094), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n990), .A2(new_n992), .ZN(new_n1107));
  INV_X1    g682(.A(new_n978), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1108), .A2(new_n976), .B1(new_n987), .B2(new_n986), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT124), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n937), .A2(new_n955), .A3(new_n991), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n991), .B1(new_n937), .B2(new_n955), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT124), .B(new_n1109), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1005), .A2(new_n1006), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n980), .B(KEYINPUT117), .C1(new_n1000), .C2(new_n1004), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n906), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n904), .A2(KEYINPUT48), .A3(new_n893), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n899), .A2(new_n893), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT48), .B1(new_n904), .B2(new_n893), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n893), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n731), .B2(new_n896), .ZN(new_n1125));
  OR3_X1    g700(.A1(new_n1124), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT46), .B1(new_n1124), .B2(G1996), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT47), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n895), .A2(new_n896), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1130), .A2(new_n897), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1057), .B2(new_n752), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1129), .B1(new_n1124), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1123), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT126), .B1(new_n1118), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1106), .A2(new_n1115), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n942), .A2(new_n944), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n960), .A2(new_n979), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1109), .B(new_n999), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1141), .A2(new_n1142), .B1(new_n960), .B2(new_n1003), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1006), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1137), .A2(new_n1144), .A3(new_n1117), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n905), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n1147), .A3(new_n1134), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1136), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g724(.A1(G229), .A2(new_n466), .A3(G227), .ZN(new_n1151));
  OAI21_X1  g725(.A(new_n1151), .B1(new_n636), .B2(new_n637), .ZN(new_n1152));
  AOI21_X1  g726(.A(new_n1152), .B1(new_n842), .B2(new_n843), .ZN(new_n1153));
  AND3_X1   g727(.A1(new_n1153), .A2(KEYINPUT127), .A3(new_n877), .ZN(new_n1154));
  AOI21_X1  g728(.A(KEYINPUT127), .B1(new_n1153), .B2(new_n877), .ZN(new_n1155));
  NOR2_X1   g729(.A1(new_n1154), .A2(new_n1155), .ZN(G308));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n877), .ZN(G225));
endmodule


