//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n212), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT64), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT65), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  AND2_X1   g0052(.A1(KEYINPUT66), .A2(G41), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT66), .A2(G41), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n253), .A2(new_n254), .A3(G45), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT67), .B1(new_n255), .B2(G1), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT66), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT66), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT67), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n263), .A3(new_n209), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n256), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G226), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G77), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  OAI211_X1 g0081(.A(G222), .B(new_n281), .C1(new_n277), .C2(new_n278), .ZN(new_n282));
  OAI211_X1 g0082(.A(G223), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT69), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n287), .A2(new_n288), .A3(new_n219), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT69), .B1(new_n266), .B2(new_n267), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n282), .A4(new_n283), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n286), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n276), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G50), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n219), .C1(G1), .C2(new_n210), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n298), .B1(new_n301), .B2(G50), .ZN(new_n302));
  AND2_X1   g0102(.A1(KEYINPUT70), .A2(G58), .ZN(new_n303));
  NOR2_X1   g0103(.A1(KEYINPUT70), .A2(G58), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT8), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT8), .A2(G58), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n305), .A2(new_n210), .A3(G33), .A4(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G20), .A2(G33), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n299), .A2(new_n219), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n302), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n296), .B(new_n314), .C1(G179), .C2(new_n294), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT3), .ZN(new_n316));
  INV_X1    g0116(.A(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(G232), .A3(new_n281), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(G238), .A3(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n279), .A2(G107), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n291), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n273), .A2(G244), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n269), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G200), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n325), .A2(G190), .A3(new_n269), .A4(new_n326), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n330), .A2(G20), .A3(new_n317), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n210), .A2(new_n317), .ZN(new_n333));
  INV_X1    g0133(.A(G77), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n332), .A2(new_n333), .B1(new_n210), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n312), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n297), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(KEYINPUT71), .A3(new_n334), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT71), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n297), .B2(G77), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n338), .A2(new_n340), .B1(new_n301), .B2(G77), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n328), .A2(new_n329), .A3(new_n342), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n327), .A2(G179), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n327), .B2(new_n295), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n315), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  INV_X1    g0148(.A(G159), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n333), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT70), .B(G58), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n201), .B1(new_n352), .B2(G68), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(new_n210), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n318), .A2(new_n210), .A3(new_n319), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n318), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n319), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n223), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n348), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT7), .B1(new_n279), .B2(new_n210), .ZN(new_n361));
  INV_X1    g0161(.A(new_n358), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n303), .B2(new_n304), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n216), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n350), .B1(new_n365), .B2(G20), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n366), .A3(KEYINPUT16), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n360), .A2(new_n312), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n306), .B1(new_n352), .B2(KEYINPUT8), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n300), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(KEYINPUT75), .C1(new_n337), .C2(new_n369), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT75), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n305), .A2(new_n300), .A3(new_n307), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n337), .B1(new_n305), .B2(new_n307), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n378));
  INV_X1    g0178(.A(G226), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G1698), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(G223), .B2(G1698), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n381), .A2(new_n279), .B1(new_n317), .B2(new_n225), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n378), .B1(new_n382), .B2(new_n291), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n269), .A2(new_n383), .A3(G179), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n269), .A2(new_n383), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n295), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT18), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n377), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n269), .A2(new_n383), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(G200), .B1(new_n269), .B2(new_n383), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n368), .B(new_n376), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n371), .A2(new_n375), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n363), .A2(new_n366), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n313), .B1(new_n398), .B2(new_n348), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n397), .B1(new_n399), .B2(new_n367), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n269), .A2(new_n383), .A3(new_n391), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n385), .B2(G200), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n388), .A2(new_n390), .A3(new_n396), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n293), .ZN(new_n405));
  OAI21_X1  g0205(.A(G200), .B1(new_n405), .B2(new_n275), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT9), .B(new_n302), .C1(new_n311), .C2(new_n313), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT9), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n313), .B1(new_n308), .B2(new_n310), .ZN(new_n409));
  INV_X1    g0209(.A(new_n302), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n276), .A2(G190), .A3(new_n293), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n406), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT10), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n407), .A2(new_n411), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n294), .B2(G200), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT10), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n413), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n347), .B(new_n404), .C1(new_n415), .C2(new_n419), .ZN(new_n420));
  OR3_X1    g0220(.A1(new_n297), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT12), .B1(new_n297), .B2(G68), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n421), .A2(new_n422), .B1(new_n301), .B2(G68), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n210), .A2(G33), .A3(G77), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n223), .A2(G20), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n424), .B(new_n425), .C1(new_n333), .C2(new_n202), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n312), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT11), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(KEYINPUT11), .A3(new_n312), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n423), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n423), .A2(new_n429), .A3(KEYINPUT73), .A4(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n262), .A2(new_n263), .A3(new_n209), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n263), .B1(new_n262), .B2(new_n209), .ZN(new_n438));
  INV_X1    g0238(.A(new_n268), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(G226), .A2(G1698), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n235), .B2(G1698), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n320), .B1(G33), .B2(G97), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n270), .A2(new_n288), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n266), .A2(KEYINPUT69), .A3(new_n267), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n443), .A2(new_n446), .B1(new_n224), .B2(new_n272), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT13), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n270), .A2(G238), .A3(new_n271), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n379), .A2(new_n281), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n235), .A2(G1698), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n277), .C2(new_n278), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G97), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n449), .B1(new_n291), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT13), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n269), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n448), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G169), .ZN(new_n459));
  INV_X1    g0259(.A(G179), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n459), .A2(KEYINPUT14), .B1(new_n460), .B2(new_n458), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n459), .A2(KEYINPUT14), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n436), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT74), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n448), .A2(G190), .A3(new_n457), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n435), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n269), .A2(new_n455), .A3(new_n456), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n456), .B1(new_n269), .B2(new_n455), .ZN(new_n468));
  OAI21_X1  g0268(.A(G200), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT72), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT72), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n458), .A2(new_n471), .A3(G200), .ZN(new_n472));
  AOI211_X1 g0272(.A(new_n464), .B(new_n466), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n472), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n465), .A2(new_n435), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT74), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n463), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n420), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n209), .A2(G33), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n297), .A2(new_n480), .A3(new_n219), .A4(new_n299), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G97), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n337), .A2(new_n205), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(G97), .B(G107), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT6), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n487), .A2(new_n205), .A3(G107), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n309), .ZN(new_n492));
  OAI21_X1  g0292(.A(G107), .B1(new_n361), .B2(new_n362), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n485), .B1(new_n494), .B2(new_n312), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT5), .B1(new_n259), .B2(new_n261), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT5), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n209), .B(G45), .C1(new_n497), .C2(G41), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(new_n270), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n498), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n497), .B1(new_n253), .B2(new_n254), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(new_n268), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(new_n281), .C1(new_n277), .C2(new_n278), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n320), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n320), .A2(G250), .A3(G1698), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n506), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n503), .B1(new_n291), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G190), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT76), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n499), .A2(new_n502), .A3(KEYINPUT76), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n514), .A2(new_n515), .B1(new_n291), .B2(new_n510), .ZN(new_n516));
  INV_X1    g0316(.A(G200), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n495), .B(new_n512), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n510), .A2(new_n291), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n295), .B1(new_n519), .B2(new_n503), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n489), .B1(new_n487), .B2(new_n486), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n521), .A2(new_n210), .B1(new_n334), .B2(new_n333), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n206), .B1(new_n357), .B2(new_n358), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n312), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(new_n483), .A3(new_n484), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n510), .A2(new_n291), .ZN(new_n526));
  INV_X1    g0326(.A(new_n515), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT76), .B1(new_n499), .B2(new_n502), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n460), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n520), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n320), .A2(new_n210), .A3(G68), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n210), .B1(new_n453), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G87), .B2(new_n207), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n535), .A2(KEYINPUT79), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT79), .B1(new_n535), .B2(new_n532), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n531), .B(new_n534), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n312), .ZN(new_n539));
  INV_X1    g0339(.A(new_n330), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n297), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n482), .A2(new_n540), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI22_X1  g0344(.A1(KEYINPUT77), .A2(new_n226), .B1(new_n260), .B2(G1), .ZN(new_n545));
  NAND2_X1  g0345(.A1(KEYINPUT77), .A2(G250), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(new_n209), .A3(G45), .A4(new_n265), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n547), .A3(new_n270), .ZN(new_n548));
  INV_X1    g0348(.A(G116), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n317), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G238), .A2(G1698), .ZN(new_n551));
  INV_X1    g0351(.A(G244), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(G1698), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n553), .B2(new_n320), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT78), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n291), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(G1698), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G238), .B2(G1698), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n558), .A2(new_n279), .B1(new_n317), .B2(new_n549), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(KEYINPUT78), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n460), .B(new_n548), .C1(new_n556), .C2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n548), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n446), .B1(new_n559), .B2(KEYINPUT78), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n554), .A2(new_n555), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n544), .B(new_n561), .C1(G169), .C2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n481), .A2(new_n225), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n541), .B(new_n567), .C1(new_n538), .C2(new_n312), .ZN(new_n568));
  OAI211_X1 g0368(.A(G190), .B(new_n548), .C1(new_n556), .C2(new_n560), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n565), .C2(new_n517), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n518), .A2(new_n530), .A3(new_n566), .A4(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n481), .A2(G116), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n337), .A2(G116), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n299), .A2(new_n219), .B1(G20), .B2(new_n549), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n508), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT20), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n572), .A2(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n287), .A2(new_n219), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n500), .B2(new_n501), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n259), .A2(new_n261), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n498), .B1(new_n581), .B2(new_n497), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n580), .A2(G270), .B1(new_n582), .B2(new_n268), .ZN(new_n583));
  OAI211_X1 g0383(.A(G264), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n584));
  OAI211_X1 g0384(.A(G257), .B(new_n281), .C1(new_n277), .C2(new_n278), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n318), .A2(G303), .A3(new_n319), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n291), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n578), .A2(G179), .A3(new_n583), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n587), .A2(new_n291), .ZN(new_n591));
  OAI211_X1 g0391(.A(G270), .B(new_n270), .C1(new_n496), .C2(new_n498), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n502), .ZN(new_n593));
  OAI21_X1  g0393(.A(G169), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n589), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n295), .B1(new_n583), .B2(new_n588), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT21), .B1(new_n596), .B2(new_n578), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n583), .A2(new_n588), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n578), .B1(new_n599), .B2(G200), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n391), .B2(new_n599), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT81), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G250), .A2(G1698), .ZN(new_n604));
  INV_X1    g0404(.A(G257), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(G1698), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(new_n320), .B1(G33), .B2(G294), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n603), .B1(new_n607), .B2(new_n446), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G250), .B2(G1698), .ZN(new_n610));
  INV_X1    g0410(.A(G294), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n610), .A2(new_n279), .B1(new_n317), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n291), .A3(KEYINPUT81), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G264), .B(new_n270), .C1(new_n496), .C2(new_n498), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n615), .A2(new_n502), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n391), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n291), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(new_n502), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n517), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT23), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n210), .B2(G107), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(new_n550), .B2(new_n210), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n210), .B(G87), .C1(new_n277), .C2(new_n278), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(KEYINPUT22), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(KEYINPUT22), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(KEYINPUT24), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT24), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n626), .B(KEYINPUT22), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n625), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n312), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT25), .ZN(new_n635));
  AOI211_X1 g0435(.A(G107), .B(new_n297), .C1(KEYINPUT80), .C2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(KEYINPUT80), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n482), .B2(G107), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n621), .A2(new_n634), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n629), .A2(KEYINPUT24), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n632), .A2(new_n631), .A3(new_n625), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n313), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(new_n639), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n482), .A2(G107), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n295), .B1(new_n614), .B2(new_n616), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n619), .A2(new_n460), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n644), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n641), .A2(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n479), .A2(new_n571), .A3(new_n602), .A4(new_n651), .ZN(G372));
  INV_X1    g0452(.A(KEYINPUT82), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n418), .B1(new_n417), .B2(new_n413), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n414), .A2(KEYINPUT10), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n419), .A2(new_n415), .A3(KEYINPUT82), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n396), .A2(new_n403), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n471), .B1(new_n458), .B2(G200), .ZN(new_n660));
  AOI211_X1 g0460(.A(KEYINPUT72), .B(new_n517), .C1(new_n448), .C2(new_n457), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n475), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n464), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n474), .A2(KEYINPUT74), .A3(new_n475), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n346), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n659), .B1(new_n667), .B2(new_n463), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n388), .A2(new_n390), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n658), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n670), .A2(new_n315), .ZN(new_n671));
  INV_X1    g0471(.A(new_n566), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n644), .A2(new_n647), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n598), .A2(new_n650), .B1(new_n673), .B2(new_n621), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n672), .B1(new_n571), .B2(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n520), .A2(new_n525), .A3(new_n529), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(KEYINPUT26), .A3(new_n566), .A4(new_n570), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n570), .A2(new_n566), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n530), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n479), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n671), .A2(new_n683), .ZN(G369));
  INV_X1    g0484(.A(new_n578), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT27), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n209), .A3(new_n210), .A4(G13), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n687), .A2(G213), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G343), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT83), .Z(new_n692));
  OAI211_X1 g0492(.A(new_n598), .B(new_n601), .C1(new_n685), .C2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT21), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n594), .B2(new_n685), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n695), .B(new_n589), .C1(new_n594), .C2(new_n590), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n691), .B(KEYINPUT83), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n578), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n651), .B1(new_n673), .B2(new_n692), .ZN(new_n702));
  INV_X1    g0502(.A(new_n648), .ZN(new_n703));
  INV_X1    g0503(.A(new_n649), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n703), .A2(new_n704), .B1(new_n634), .B2(new_n640), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(new_n692), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n651), .A2(new_n696), .A3(new_n692), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n581), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n213), .A2(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G1), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n217), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n588), .A2(G179), .A3(new_n592), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n618), .A2(new_n502), .A3(new_n615), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n565), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(KEYINPUT84), .A3(KEYINPUT30), .A4(new_n511), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT84), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n511), .A2(new_n565), .A3(new_n718), .A4(new_n719), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n565), .A2(new_n719), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n460), .A3(new_n728), .A4(new_n599), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n721), .A2(new_n725), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n730), .B2(new_n697), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT85), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n697), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT85), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n571), .A2(new_n602), .A3(new_n651), .A4(new_n692), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n733), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n682), .B2(new_n692), .ZN(new_n744));
  AOI211_X1 g0544(.A(KEYINPUT29), .B(new_n697), .C1(new_n675), .C2(new_n681), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n717), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(new_n699), .A2(G330), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT86), .Z(new_n751));
  INV_X1    g0551(.A(G13), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n209), .B1(new_n753), .B2(G45), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n713), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT87), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(new_n700), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n219), .B1(G20), .B2(new_n295), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n210), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(new_n391), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n206), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G159), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT32), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n210), .A2(new_n460), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n391), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n763), .B(new_n768), .C1(G50), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n352), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n769), .A2(G190), .A3(new_n517), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n320), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n770), .A2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n391), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n210), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n777), .A2(new_n223), .B1(new_n205), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n769), .A2(new_n764), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n775), .B(new_n780), .C1(G77), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT90), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n772), .B(new_n783), .C1(new_n225), .C2(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n777), .A2(new_n790), .B1(new_n774), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT92), .Z(new_n793));
  INV_X1    g0593(.A(G329), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n279), .B1(new_n765), .B2(new_n794), .C1(new_n781), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n771), .ZN(new_n797));
  INV_X1    g0597(.A(G326), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n797), .A2(new_n798), .B1(new_n762), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n779), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n796), .B(new_n800), .C1(G294), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n788), .B(KEYINPUT91), .Z(new_n804));
  OAI211_X1 g0604(.A(new_n793), .B(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n760), .B1(new_n789), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n756), .B(KEYINPUT88), .Z(new_n807));
  NAND3_X1  g0607(.A1(new_n752), .A2(new_n317), .A3(KEYINPUT89), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT89), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(G13), .B2(G33), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n759), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n213), .A2(new_n320), .ZN(new_n816));
  INV_X1    g0616(.A(G355), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n817), .B1(G116), .B2(new_n213), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n251), .A2(G45), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n213), .A2(new_n279), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n260), .B2(new_n218), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n807), .B1(new_n815), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n806), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n813), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n699), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n758), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  AOI21_X1  g0628(.A(new_n697), .B1(new_n675), .B2(new_n681), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT93), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n344), .A2(new_n345), .A3(new_n692), .ZN(new_n831));
  INV_X1    g0631(.A(new_n342), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n697), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n343), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n830), .B(new_n831), .C1(new_n834), .C2(new_n666), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n343), .A2(new_n833), .B1(new_n344), .B2(new_n345), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n344), .A2(new_n345), .A3(new_n692), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT93), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n829), .B(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n756), .B1(new_n742), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n742), .B2(new_n840), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n812), .A2(new_n760), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n807), .B1(G77), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n762), .A2(new_n225), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G303), .B2(new_n771), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n205), .B2(new_n779), .C1(new_n799), .C2(new_n777), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n279), .B1(new_n781), .B2(new_n549), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n774), .A2(new_n611), .B1(new_n765), .B2(new_n795), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n206), .B2(new_n804), .ZN(new_n851));
  INV_X1    g0651(.A(new_n774), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(G143), .B1(new_n782), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(G150), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n777), .B2(new_n854), .C1(new_n855), .C2(new_n797), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n762), .A2(new_n223), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n320), .B1(new_n860), .B2(new_n765), .C1(new_n779), .C2(new_n773), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n857), .B2(new_n856), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n804), .A2(new_n202), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n844), .B1(new_n865), .B2(new_n759), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n812), .B2(new_n839), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(new_n867), .ZN(G384));
  OR2_X1    g0668(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n869), .A2(G116), .A3(new_n220), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT36), .Z(new_n872));
  NAND3_X1  g0672(.A1(new_n218), .A2(G77), .A3(new_n364), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n202), .A2(G68), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n209), .B(G13), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n690), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n669), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n641), .B1(new_n705), .B2(new_n696), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n518), .A2(new_n530), .A3(new_n566), .A4(new_n570), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n566), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n677), .A2(new_n680), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n839), .B(new_n692), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n831), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n435), .A2(new_n692), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n477), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n885), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n665), .A2(new_n463), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n370), .B1(new_n337), .B2(new_n369), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n368), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n386), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n690), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n394), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n295), .B1(new_n269), .B2(new_n383), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(G179), .B2(new_n385), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT94), .B1(new_n400), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT37), .B1(new_n400), .B2(new_n402), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT94), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n377), .A2(new_n901), .A3(new_n386), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT95), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n377), .B2(new_n690), .ZN(new_n905));
  AOI211_X1 g0705(.A(KEYINPUT95), .B(new_n877), .C1(new_n368), .C2(new_n376), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n896), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n894), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n404), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n878), .B1(new_n890), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT96), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT39), .B1(new_n911), .B2(new_n912), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n917));
  XOR2_X1   g0717(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n918));
  NOR2_X1   g0718(.A1(new_n392), .A2(new_n393), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT97), .B1(new_n377), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT97), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n402), .A2(new_n921), .A3(new_n368), .A4(new_n376), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n387), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT37), .B1(new_n907), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT95), .B1(new_n400), .B2(new_n877), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n377), .A2(new_n904), .A3(new_n690), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n927), .A2(new_n902), .A3(new_n899), .A4(new_n900), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n924), .A2(new_n928), .B1(new_n404), .B2(new_n907), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n917), .B(new_n918), .C1(new_n929), .C2(KEYINPUT38), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n916), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n463), .A2(new_n697), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n915), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n914), .A2(KEYINPUT96), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n479), .B1(new_n744), .B2(new_n745), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n671), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n839), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n886), .B2(new_n888), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n917), .B1(new_n929), .B2(KEYINPUT38), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n736), .A2(new_n738), .A3(new_n740), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT40), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n911), .A2(new_n912), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(new_n944), .A4(new_n942), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n479), .A2(new_n944), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  INV_X1    g0753(.A(G330), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n940), .A2(new_n955), .B1(new_n209), .B2(new_n753), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n940), .A2(new_n955), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n876), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT99), .ZN(G367));
  OAI221_X1 g0759(.A(new_n814), .B1(new_n213), .B2(new_n330), .C1(new_n241), .C2(new_n820), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n762), .A2(new_n205), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n797), .A2(new_n795), .B1(new_n206), .B2(new_n779), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n961), .B(new_n962), .C1(G294), .C2(new_n776), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT46), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n788), .B2(new_n549), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n320), .B1(new_n782), .B2(G283), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n852), .A2(G303), .B1(new_n766), .B2(G317), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n963), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n804), .A2(new_n964), .A3(new_n549), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n776), .A2(G159), .B1(new_n782), .B2(G50), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT106), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n762), .A2(new_n334), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n779), .A2(new_n223), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(G143), .C2(new_n771), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n320), .B1(new_n774), .B2(new_n854), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G137), .B2(new_n766), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(new_n773), .C2(new_n788), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n968), .A2(new_n969), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  OAI211_X1 g0779(.A(new_n807), .B(new_n960), .C1(new_n979), .C2(new_n760), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n692), .A2(new_n568), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT100), .Z(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(new_n679), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n679), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n825), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n754), .ZN(new_n988));
  INV_X1    g0788(.A(new_n708), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n696), .A2(new_n692), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n641), .A2(new_n650), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n709), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n676), .A2(new_n697), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n525), .A2(new_n697), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n518), .A2(new_n530), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n990), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n996), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n710), .A2(KEYINPUT45), .A3(new_n999), .A4(new_n709), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n993), .A2(new_n997), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n993), .A2(new_n997), .A3(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n989), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n998), .A2(new_n1000), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n708), .A2(new_n1009), .A3(new_n1006), .A4(new_n1005), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n702), .A2(new_n706), .A3(new_n991), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n710), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n701), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n700), .A3(new_n710), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n742), .A2(new_n746), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1011), .B1(new_n1017), .B2(KEYINPUT104), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT104), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n742), .A2(new_n1016), .A3(new_n746), .A4(new_n1019), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n1018), .A2(KEYINPUT105), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT105), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n748), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n713), .B(KEYINPUT41), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n988), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n996), .A2(new_n650), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(new_n530), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n697), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n710), .A2(new_n997), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT42), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(KEYINPUT42), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n983), .A2(new_n984), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT43), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n983), .A2(KEYINPUT43), .A3(new_n984), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1034), .A2(new_n1039), .A3(KEYINPUT102), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT102), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n1033), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1033), .A2(new_n1036), .A3(new_n1035), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(KEYINPUT101), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT101), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1040), .A2(new_n1047), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n708), .A2(new_n997), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1046), .A2(new_n1050), .A3(new_n1048), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n987), .B1(new_n1026), .B2(new_n1054), .ZN(G387));
  NAND3_X1  g0855(.A1(new_n702), .A2(new_n706), .A3(new_n813), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n816), .A2(new_n714), .B1(G107), .B2(new_n213), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n238), .A2(new_n260), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n714), .ZN(new_n1059));
  AOI211_X1 g0859(.A(G45), .B(new_n1059), .C1(G68), .C2(G77), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n332), .A2(G50), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT50), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n820), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1057), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n807), .B1(new_n1064), .B2(new_n815), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n774), .A2(new_n202), .B1(new_n765), .B2(new_n854), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n279), .B(new_n1066), .C1(G68), .C2(new_n782), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n779), .A2(new_n330), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n961), .B(new_n1068), .C1(G159), .C2(new_n771), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n788), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(G77), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n776), .A2(new_n369), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n788), .A2(new_n611), .B1(new_n799), .B2(new_n779), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n852), .A2(G317), .B1(new_n782), .B2(G303), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n777), .B2(new_n795), .C1(new_n791), .C2(new_n797), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT49), .Z(new_n1080));
  OAI221_X1 g0880(.A(new_n279), .B1(new_n765), .B2(new_n798), .C1(new_n762), .C2(new_n549), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1073), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1065), .B1(new_n1082), .B2(new_n759), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1016), .A2(new_n988), .B1(new_n1056), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n748), .A2(new_n1016), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n713), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1017), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1085), .B2(new_n1087), .ZN(G393));
  AOI21_X1  g0888(.A(new_n713), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1011), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n988), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n814), .B1(new_n205), .B2(new_n213), .C1(new_n246), .C2(new_n820), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT107), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n807), .A2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n797), .A2(new_n854), .B1(new_n349), .B2(new_n774), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n779), .A2(new_n334), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n845), .B(new_n1098), .C1(G50), .C2(new_n776), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1070), .A2(G68), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n320), .B1(new_n781), .B2(new_n332), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G143), .B2(new_n766), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1097), .A2(new_n1099), .A3(new_n1100), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G317), .A2(new_n771), .B1(new_n852), .B2(G311), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT108), .B(KEYINPUT52), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n763), .B1(G116), .B2(new_n801), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n803), .B2(new_n777), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n279), .B1(new_n765), .B2(new_n791), .C1(new_n781), .C2(new_n611), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1106), .B(new_n1110), .C1(new_n799), .C2(new_n788), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n760), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1093), .A2(KEYINPUT107), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1095), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n825), .B2(new_n999), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1090), .A2(new_n1092), .A3(new_n1115), .ZN(G390));
  INV_X1    g0916(.A(new_n944), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n954), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n942), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n890), .A2(new_n932), .A3(new_n943), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n477), .A2(new_n885), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n887), .B1(new_n665), .B2(new_n463), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n837), .B1(new_n829), .B2(new_n839), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n932), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n931), .B1(new_n1126), .B2(KEYINPUT109), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT109), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1128), .B(new_n932), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1121), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1119), .B1(new_n1130), .B2(KEYINPUT110), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n883), .A2(new_n831), .B1(new_n886), .B2(new_n888), .ZN(new_n1132));
  OAI21_X1  g0932(.A(KEYINPUT109), .B1(new_n1132), .B2(new_n933), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n916), .A2(new_n930), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n1129), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1120), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT110), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n741), .A2(G330), .A3(new_n839), .A4(new_n889), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1135), .A2(new_n1120), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT111), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1135), .A2(KEYINPUT111), .A3(new_n1120), .A4(new_n1139), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1131), .A2(new_n1138), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1134), .A2(new_n811), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n807), .B1(new_n369), .B2(new_n843), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n279), .B1(new_n804), .B2(new_n225), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT113), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n206), .A2(new_n777), .B1(new_n797), .B2(new_n799), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1149), .A2(new_n859), .A3(new_n1098), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G97), .A2(new_n782), .B1(new_n766), .B2(G294), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n549), .C2(new_n774), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n788), .A2(KEYINPUT53), .A3(new_n854), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n279), .B1(new_n766), .B2(G125), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n860), .B2(new_n774), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT112), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1155), .B1(new_n782), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G159), .A2(new_n801), .B1(new_n776), .B2(G137), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT53), .B1(new_n788), .B2(new_n854), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n762), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n771), .A2(G128), .B1(new_n1161), .B2(G50), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1148), .A2(new_n1152), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1146), .B1(new_n1164), .B2(new_n759), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1144), .A2(new_n988), .B1(new_n1145), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1118), .A2(new_n479), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n671), .A2(new_n938), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1124), .B1(new_n742), .B2(new_n941), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1119), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n884), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1117), .A2(new_n954), .A3(new_n941), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1139), .B(new_n1125), .C1(new_n889), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1168), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1086), .B1(new_n1144), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1119), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1135), .A2(KEYINPUT110), .A3(new_n1120), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1138), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(new_n1174), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1166), .B1(new_n1175), .B2(new_n1181), .ZN(G378));
  NAND2_X1  g0982(.A1(new_n950), .A2(G330), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n419), .A2(new_n415), .A3(KEYINPUT82), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT82), .B1(new_n419), .B2(new_n415), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n315), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n314), .A2(new_n690), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT55), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n1191));
  NAND3_X1  g0991(.A1(new_n658), .A2(new_n315), .A3(new_n1188), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1191), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1183), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1195), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n950), .A2(G330), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT116), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n935), .A2(new_n936), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n954), .B(new_n1195), .C1(new_n946), .C2(new_n949), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1197), .B1(new_n950), .B2(G330), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1200), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n937), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1202), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1195), .A2(new_n811), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n756), .B1(G50), .B2(new_n843), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n205), .A2(new_n777), .B1(new_n797), .B2(new_n549), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n973), .B(new_n1210), .C1(new_n352), .C2(new_n1161), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n712), .A2(new_n279), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G283), .B2(new_n766), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n852), .A2(G107), .B1(new_n782), .B2(new_n540), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1071), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1212), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1070), .A2(new_n1157), .ZN(new_n1220));
  INV_X1    g1020(.A(G128), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n774), .A2(new_n1221), .B1(new_n781), .B2(new_n855), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G132), .B2(new_n776), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G150), .A2(new_n801), .B1(new_n771), .B2(G125), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1220), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT59), .Z(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT114), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1161), .A2(G159), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1227), .A2(KEYINPUT114), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1219), .B1(new_n1216), .B2(new_n1215), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1209), .B1(new_n1233), .B2(new_n759), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1207), .A2(new_n988), .B1(new_n1208), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1168), .B1(new_n1144), .B2(new_n1174), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n937), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n937), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1086), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1168), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1180), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT57), .B1(new_n1243), .B2(new_n1207), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1235), .B1(new_n1241), .B2(new_n1244), .ZN(G375));
  NAND2_X1  g1045(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1242), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1171), .A2(new_n1168), .A3(new_n1173), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1025), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1124), .A2(new_n811), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n807), .B1(G68), .B2(new_n843), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n771), .A2(G294), .B1(new_n782), .B2(G107), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n549), .B2(new_n777), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT117), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n279), .B1(new_n765), .B2(new_n803), .C1(new_n774), .C2(new_n799), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1255), .A2(new_n972), .A3(new_n1068), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(new_n205), .C2(new_n804), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n797), .A2(new_n860), .B1(new_n773), .B2(new_n762), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G50), .B2(new_n801), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n320), .B1(new_n765), .B2(new_n1221), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n774), .A2(new_n855), .B1(new_n781), .B2(new_n854), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n776), .C2(new_n1157), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1259), .B(new_n1262), .C1(new_n804), .C2(new_n349), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n760), .B1(new_n1257), .B2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1251), .A2(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1246), .A2(new_n988), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(new_n1266), .ZN(G381));
  NAND2_X1  g1067(.A1(new_n1017), .A2(KEYINPUT104), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(new_n1020), .A3(new_n1091), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT105), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1018), .A2(KEYINPUT105), .A3(new_n1020), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n747), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n754), .B1(new_n1273), .B2(new_n1024), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1046), .A2(new_n1050), .A3(new_n1048), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1050), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n986), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(G390), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OR4_X1    g1080(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1281));
  OR4_X1    g1081(.A1(G378), .A2(G375), .A3(new_n1280), .A4(new_n1281), .ZN(G407));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G343), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(G375), .A2(G378), .A3(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(KEYINPUT118), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G213), .A3(G407), .ZN(G409));
  OAI211_X1 g1088(.A(G378), .B(new_n1235), .C1(new_n1241), .C2(new_n1244), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1145), .A2(new_n1165), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1291), .B2(new_n754), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n713), .B1(new_n1291), .B2(new_n1247), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1180), .B2(new_n1293), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1243), .A2(new_n1025), .A3(new_n1207), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n988), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1208), .A2(new_n1234), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1294), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1289), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(G384), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(KEYINPUT119), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1248), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1171), .A2(KEYINPUT60), .A3(new_n1168), .A4(new_n1173), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(new_n1247), .A3(new_n1086), .A4(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1302), .B1(new_n1306), .B2(new_n1266), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT119), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(G384), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1306), .A2(KEYINPUT119), .A3(new_n1301), .A4(new_n1266), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1300), .A2(new_n1285), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT62), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1300), .A2(new_n1285), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1284), .A2(G2897), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1284), .A2(KEYINPUT122), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1313), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1317), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1318), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1320), .B(new_n1321), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1319), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1316), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1300), .A2(new_n1326), .A3(new_n1285), .A4(new_n1313), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1315), .A2(new_n1324), .A3(new_n1325), .A4(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT124), .ZN(new_n1329));
  OAI21_X1  g1129(.A(G390), .B1(new_n1278), .B2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(G387), .A2(KEYINPUT124), .A3(new_n1279), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(G393), .B(new_n827), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1330), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G387), .A2(G390), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(KEYINPUT123), .ZN(new_n1336));
  OR2_X1    g1136(.A1(new_n1333), .A2(KEYINPUT123), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1335), .A2(new_n1280), .A3(new_n1336), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1334), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1328), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1316), .A2(KEYINPUT121), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT121), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1300), .A2(new_n1343), .A3(new_n1285), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1342), .A2(new_n1323), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1339), .A2(new_n1325), .ZN(new_n1346));
  AOI211_X1 g1146(.A(new_n1302), .B(new_n1309), .C1(new_n1306), .C2(new_n1266), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1312), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AOI211_X1 g1149(.A(new_n1284), .B(new_n1349), .C1(new_n1289), .C2(new_n1299), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1346), .B1(new_n1350), .B2(KEYINPUT63), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT120), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1350), .B2(KEYINPUT63), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT63), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1314), .A2(KEYINPUT120), .A3(new_n1354), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1345), .A2(new_n1351), .A3(new_n1353), .A4(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1341), .A2(new_n1356), .ZN(G405));
  NAND2_X1  g1157(.A1(G375), .A2(new_n1294), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT125), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1358), .A2(new_n1359), .A3(new_n1289), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(G375), .A2(KEYINPUT125), .A3(new_n1294), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT127), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT126), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1362), .B1(new_n1349), .B2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1365));
  AOI22_X1  g1165(.A1(new_n1360), .A2(new_n1361), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1360), .A2(new_n1364), .A3(new_n1361), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1367), .A2(new_n1339), .A3(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1368), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1340), .B1(new_n1370), .B2(new_n1366), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1369), .A2(new_n1371), .ZN(G402));
endmodule


