//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  AOI21_X1  g002(.A(G1gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(KEYINPUT97), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(KEYINPUT97), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n204), .A3(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n216), .B1(new_n213), .B2(KEYINPUT15), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT96), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT96), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n214), .A2(new_n217), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT15), .B(new_n213), .C1(new_n223), .C2(new_n216), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n212), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n206), .A2(new_n204), .A3(new_n208), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(new_n209), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(new_n229), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n234), .B(new_n235), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n237), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n232), .A2(KEYINPUT18), .A3(new_n236), .A4(new_n237), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT11), .B(G169gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G197gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n249), .B(KEYINPUT12), .Z(new_n250));
  OR2_X1    g049(.A1(new_n250), .A2(KEYINPUT95), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(KEYINPUT95), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n245), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n240), .A2(new_n243), .A3(new_n250), .A4(new_n244), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n254), .A2(KEYINPUT98), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(KEYINPUT98), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT77), .ZN(new_n259));
  INV_X1    g058(.A(G148gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(G141gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(G141gat), .ZN(new_n262));
  INV_X1    g061(.A(G141gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT2), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n268));
  AND2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(KEYINPUT78), .A3(new_n266), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n265), .A2(new_n267), .A3(new_n271), .A4(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G141gat), .B(G148gat), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n266), .B(new_n274), .C1(new_n277), .C2(KEYINPUT2), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT79), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n276), .A2(KEYINPUT79), .A3(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT22), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G211gat), .A2(G218gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(KEYINPUT75), .A2(KEYINPUT22), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G211gat), .B(G218gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n284), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G228gat), .ZN(new_n299));
  INV_X1    g098(.A(G233gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n276), .A2(new_n296), .A3(new_n278), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n284), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n290), .A2(new_n292), .ZN(new_n304));
  INV_X1    g103(.A(new_n291), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n306), .B2(new_n307), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n279), .B1(new_n312), .B2(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n301), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT83), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n295), .A2(new_n296), .B1(new_n278), .B2(new_n276), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n308), .B1(new_n302), .B2(new_n284), .ZN(new_n318));
  OAI211_X1 g117(.A(KEYINPUT83), .B(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n311), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT86), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n319), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT86), .A3(new_n311), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(G22gat), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT87), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(G50gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(G78gat), .ZN(new_n333));
  INV_X1    g132(.A(G106gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n323), .A2(new_n336), .A3(G22gat), .A4(new_n328), .ZN(new_n337));
  XOR2_X1   g136(.A(KEYINPUT84), .B(G22gat), .Z(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n327), .A2(new_n311), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n330), .A2(new_n335), .A3(new_n337), .A4(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n335), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n339), .B1(new_n327), .B2(new_n311), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT85), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT85), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n347), .B(new_n343), .C1(new_n340), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n342), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  INV_X1    g150(.A(G169gat), .ZN(new_n352));
  INV_X1    g151(.A(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n354), .A2(KEYINPUT26), .ZN(new_n355));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(KEYINPUT26), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359));
  INV_X1    g158(.A(G183gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT27), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT27), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(G183gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(G183gat), .ZN(new_n365));
  AOI21_X1  g164(.A(G190gat), .B1(new_n365), .B2(KEYINPUT69), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT28), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n360), .A2(KEYINPUT27), .ZN(new_n368));
  INV_X1    g167(.A(G190gat), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT28), .A4(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n351), .B(new_n358), .C1(new_n367), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT64), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n360), .A3(new_n369), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n351), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n374), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n356), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(KEYINPUT23), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT65), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(KEYINPUT25), .ZN(new_n385));
  AND2_X1   g184(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n386));
  NOR2_X1   g185(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n354), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT25), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n383), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT67), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n360), .A3(new_n369), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n376), .A3(new_n377), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT68), .ZN(new_n398));
  AND3_X1   g197(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n396), .A4(new_n395), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n393), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n392), .B1(new_n404), .B2(new_n356), .ZN(new_n405));
  INV_X1    g204(.A(G134gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G127gat), .ZN(new_n407));
  INV_X1    g206(.A(G127gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(G134gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n409), .A3(KEYINPUT70), .ZN(new_n410));
  XNOR2_X1  g209(.A(G113gat), .B(G120gat), .ZN(new_n411));
  OAI221_X1 g210(.A(new_n410), .B1(KEYINPUT70), .B2(new_n407), .C1(KEYINPUT1), .C2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n407), .A2(new_n409), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n414));
  INV_X1    g213(.A(G120gat), .ZN(new_n415));
  OR2_X1    g214(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n415), .A2(G113gat), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n413), .B(new_n414), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n391), .A2(new_n405), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n412), .A2(new_n420), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n382), .A2(new_n389), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT28), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT69), .B1(new_n365), .B2(new_n368), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT69), .B1(new_n360), .B2(KEYINPUT27), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n369), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n429), .A2(new_n370), .B1(G183gat), .B2(G190gat), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n424), .B1(new_n430), .B2(new_n358), .ZN(new_n431));
  INV_X1    g230(.A(new_n393), .ZN(new_n432));
  INV_X1    g231(.A(new_n396), .ZN(new_n433));
  NOR3_X1   g232(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n402), .B1(new_n435), .B2(new_n401), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n397), .A2(KEYINPUT68), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n356), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT25), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n423), .B1(new_n431), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n422), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  OAI22_X1  g242(.A1(new_n441), .A2(new_n442), .B1(KEYINPUT32), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G15gat), .B(G43gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(G71gat), .ZN(new_n446));
  INV_X1    g245(.A(G99gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT73), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT32), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n421), .B1(new_n391), .B2(new_n405), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n431), .A2(new_n439), .A3(new_n423), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n442), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(KEYINPUT33), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n450), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n442), .B1(new_n452), .B2(new_n453), .ZN(new_n459));
  INV_X1    g258(.A(new_n457), .ZN(new_n460));
  NOR4_X1   g259(.A1(new_n459), .A2(KEYINPUT73), .A3(new_n451), .A4(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n449), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT34), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n454), .A2(new_n455), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT34), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n449), .B(new_n465), .C1(new_n458), .C2(new_n461), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n464), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT32), .B(new_n457), .C1(new_n441), .C2(new_n442), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT73), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n456), .A2(new_n450), .A3(new_n457), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n465), .B1(new_n472), .B2(new_n449), .ZN(new_n473));
  INV_X1    g272(.A(new_n466), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n350), .A2(new_n467), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n477));
  INV_X1    g276(.A(G226gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n300), .ZN(new_n479));
  INV_X1    g278(.A(new_n356), .ZN(new_n480));
  AOI211_X1 g279(.A(new_n480), .B(new_n393), .C1(new_n398), .C2(new_n403), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n372), .B(new_n390), .C1(new_n481), .C2(new_n392), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n479), .B1(new_n482), .B2(new_n284), .ZN(new_n483));
  INV_X1    g282(.A(new_n479), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n431), .B2(new_n439), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n309), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G64gat), .B(G92gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G36gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT76), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(new_n207), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(new_n479), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT29), .B1(new_n431), .B2(new_n439), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(new_n308), .C1(new_n493), .C2(new_n479), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n486), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n486), .B2(new_n494), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT30), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n486), .A2(new_n494), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n499), .A2(KEYINPUT30), .A3(new_n490), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n477), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G1gat), .B(G29gat), .Z(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G57gat), .B(G85gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n504), .B(new_n505), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n421), .A2(new_n302), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n283), .B2(KEYINPUT3), .ZN(new_n508));
  INV_X1    g307(.A(new_n279), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n423), .A2(new_n509), .A3(KEYINPUT4), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT4), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n421), .B2(new_n279), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G225gat), .A2(G233gat), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n508), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT5), .ZN(new_n517));
  INV_X1    g316(.A(new_n282), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT79), .B1(new_n276), .B2(new_n278), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n421), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n421), .A2(new_n279), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n514), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n517), .B1(new_n523), .B2(KEYINPUT80), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT80), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n423), .B1(new_n281), .B2(new_n282), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(new_n521), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n527), .B2(new_n514), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n516), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n506), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n508), .A2(new_n513), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n514), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT80), .B(new_n515), .C1(new_n526), .C2(new_n521), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT5), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n523), .A2(KEYINPUT80), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n506), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n530), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n532), .A2(new_n533), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n539), .A2(new_n530), .A3(KEYINPUT6), .A4(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n499), .A2(new_n490), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n486), .A2(new_n491), .A3(new_n494), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT30), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT89), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n501), .A2(new_n544), .A3(new_n545), .A4(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT94), .B1(new_n476), .B2(new_n551), .ZN(new_n552));
  AND4_X1   g351(.A1(new_n545), .A2(new_n501), .A3(new_n544), .A4(new_n550), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n553), .A2(new_n556), .A3(new_n557), .A4(new_n350), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n542), .A2(new_n543), .B1(new_n549), .B2(new_n548), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n350), .A2(new_n475), .A3(new_n467), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT35), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n534), .A2(KEYINPUT39), .A3(new_n514), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(new_n540), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n527), .A2(new_n514), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n566), .B(KEYINPUT39), .C1(new_n534), .C2(new_n514), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n568), .A2(KEYINPUT40), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n565), .A2(KEYINPUT40), .A3(new_n567), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n570), .A2(new_n541), .ZN(new_n571));
  INV_X1    g370(.A(new_n550), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT89), .B1(new_n548), .B2(new_n549), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n569), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n486), .A2(new_n575), .A3(new_n494), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n499), .A2(KEYINPUT37), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n580), .A2(KEYINPUT90), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(KEYINPUT90), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n490), .B(new_n579), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT92), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n580), .B(KEYINPUT90), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n585), .A2(new_n586), .A3(new_n490), .A4(new_n579), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n544), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n575), .B1(new_n486), .B2(new_n494), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT93), .B1(new_n590), .B2(new_n491), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n576), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n590), .A2(KEYINPUT93), .A3(new_n491), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n577), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(new_n594), .A3(new_n547), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n350), .B(new_n574), .C1(new_n588), .C2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n560), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n350), .A2(KEYINPUT88), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT88), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n342), .B2(new_n349), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n597), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n556), .A2(KEYINPUT74), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n475), .A2(new_n467), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(KEYINPUT74), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n602), .A2(KEYINPUT74), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n596), .A2(new_n601), .A3(new_n603), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n258), .B1(new_n563), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  NAND3_X1  g414(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G99gat), .B(G106gat), .Z(new_n618));
  AND2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT103), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n617), .B(new_n618), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n231), .B2(new_n230), .ZN(new_n627));
  AND2_X1   g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n622), .A2(new_n625), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n235), .ZN(new_n632));
  XOR2_X1   g431(.A(G190gat), .B(G218gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT104), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(KEYINPUT104), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n637), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n630), .A2(new_n632), .A3(new_n635), .A4(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n638), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n638), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G71gat), .B(G78gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT99), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT9), .ZN(new_n654));
  INV_X1    g453(.A(G71gat), .ZN(new_n655));
  INV_X1    g454(.A(G78gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G57gat), .A2(G64gat), .ZN(new_n658));
  INV_X1    g457(.A(G57gat), .ZN(new_n659));
  INV_X1    g458(.A(G64gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n653), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n660), .B1(new_n664), .B2(new_n659), .ZN(new_n665));
  NAND3_X1  g464(.A1(KEYINPUT100), .A2(G57gat), .A3(G64gat), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n652), .A2(new_n657), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n234), .B1(new_n668), .B2(KEYINPUT21), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n360), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n669), .A2(new_n360), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n651), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n670), .A3(new_n650), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n649), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n668), .A2(KEYINPUT21), .ZN(new_n678));
  XNOR2_X1  g477(.A(G127gat), .B(G155gat), .ZN(new_n679));
  INV_X1    g478(.A(G211gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(G231gat), .A2(G233gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n678), .B(new_n683), .Z(new_n684));
  NAND3_X1  g483(.A1(new_n673), .A2(new_n675), .A3(new_n649), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n677), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n684), .ZN(new_n687));
  INV_X1    g486(.A(new_n685), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n676), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(G230gat), .A2(G233gat), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n663), .A2(new_n667), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n623), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n621), .A2(new_n663), .A3(new_n667), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT10), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n622), .A2(new_n668), .A3(new_n625), .A4(KEYINPUT10), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n692), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n695), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n692), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(G120gat), .B(G148gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G204gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT105), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G176gat), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n697), .A2(new_n698), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n691), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n700), .A2(new_n692), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n705), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n647), .A2(new_n690), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n609), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n589), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g516(.A1(new_n572), .A2(new_n573), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n203), .A2(new_n207), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n724), .B(new_n725), .C1(new_n207), .C2(new_n719), .ZN(G1325gat));
  INV_X1    g525(.A(G15gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n603), .A2(new_n607), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n556), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n727), .B2(new_n731), .ZN(G1326gat));
  OR2_X1    g531(.A1(new_n598), .A2(new_n600), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n714), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT43), .B(G22gat), .Z(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1327gat));
  AOI21_X1  g536(.A(new_n647), .B1(new_n563), .B2(new_n608), .ZN(new_n738));
  INV_X1    g537(.A(new_n690), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n712), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n258), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n738), .A2(new_n218), .A3(new_n589), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT45), .ZN(new_n743));
  AOI221_X4 g542(.A(KEYINPUT107), .B1(KEYINPUT35), .B2(new_n561), .C1(new_n552), .C2(new_n558), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n559), .B2(new_n562), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n608), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT44), .B1(new_n747), .B2(new_n646), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n738), .A2(KEYINPUT44), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n257), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n254), .B(KEYINPUT98), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(KEYINPUT106), .A3(new_n253), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR4_X1   g556(.A1(new_n748), .A2(new_n749), .A3(new_n544), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n743), .B1(new_n758), .B2(new_n218), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1328gat));
  NAND2_X1  g560(.A1(new_n747), .A2(new_n646), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n749), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n756), .ZN(new_n765));
  OAI21_X1  g564(.A(G36gat), .B1(new_n765), .B2(new_n718), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n738), .A2(new_n741), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n767), .A2(G36gat), .A3(new_n718), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1329gat));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771));
  INV_X1    g570(.A(new_n608), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n563), .A2(KEYINPUT107), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n559), .A2(new_n745), .A3(new_n562), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n763), .B1(new_n775), .B2(new_n647), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n738), .A2(KEYINPUT44), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n776), .A2(new_n728), .A3(new_n756), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(G43gat), .ZN(new_n779));
  INV_X1    g578(.A(G43gat), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n738), .A2(new_n780), .A3(new_n556), .A4(new_n741), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT109), .Z(new_n782));
  OAI21_X1  g581(.A(new_n771), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n764), .A2(KEYINPUT110), .A3(new_n728), .A4(new_n756), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n785), .A2(new_n786), .A3(G43gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(KEYINPUT47), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(G1330gat));
  OAI21_X1  g588(.A(G50gat), .B1(new_n765), .B2(new_n350), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n767), .A2(G50gat), .A3(new_n734), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT48), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n764), .A2(new_n733), .A3(new_n756), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n794), .B2(G50gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(KEYINPUT48), .B2(new_n795), .ZN(G1331gat));
  NOR3_X1   g595(.A1(new_n775), .A2(new_n739), .A3(new_n646), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n754), .A2(new_n712), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n544), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(new_n659), .ZN(G1332gat));
  XOR2_X1   g600(.A(new_n718), .B(KEYINPUT111), .Z(new_n802));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  AND2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n803), .B2(new_n804), .ZN(G1333gat));
  OAI21_X1  g606(.A(G71gat), .B1(new_n799), .B2(new_n729), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n797), .A2(new_n655), .A3(new_n556), .A4(new_n798), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n808), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(G1334gat));
  NOR2_X1   g612(.A1(new_n799), .A2(new_n734), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(new_n656), .ZN(G1335gat));
  NOR2_X1   g614(.A1(new_n754), .A2(new_n690), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n776), .A2(new_n711), .A3(new_n777), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n611), .A3(new_n544), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n747), .A2(new_n646), .A3(new_n816), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT51), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n747), .A2(new_n821), .A3(new_n646), .A4(new_n816), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n820), .A2(new_n589), .A3(new_n711), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n818), .B1(new_n611), .B2(new_n823), .ZN(G1336gat));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(G92gat), .C1(new_n817), .C2(new_n802), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n802), .A2(G92gat), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n820), .A2(new_n711), .A3(new_n822), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT52), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n828), .ZN(new_n832));
  INV_X1    g631(.A(new_n718), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n764), .A2(new_n833), .A3(new_n711), .A4(new_n816), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n832), .A2(new_n829), .B1(new_n834), .B2(G92gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n831), .B1(new_n835), .B2(new_n825), .ZN(G1337gat));
  OAI21_X1  g635(.A(G99gat), .B1(new_n817), .B2(new_n729), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n820), .A2(new_n447), .A3(new_n711), .A4(new_n822), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n604), .B2(new_n838), .ZN(G1338gat));
  INV_X1    g638(.A(new_n816), .ZN(new_n840));
  NOR4_X1   g639(.A1(new_n748), .A2(new_n749), .A3(new_n712), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n334), .B1(new_n841), .B2(new_n733), .ZN(new_n842));
  INV_X1    g641(.A(new_n350), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n820), .A2(new_n843), .A3(new_n711), .A4(new_n822), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(G106gat), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT53), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G106gat), .B1(new_n817), .B2(new_n350), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n847), .B(new_n848), .C1(G106gat), .C2(new_n844), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(G1339gat));
  NAND3_X1  g649(.A1(new_n697), .A2(new_n698), .A3(new_n692), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n708), .A2(new_n851), .A3(KEYINPUT54), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n705), .B1(new_n699), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(KEYINPUT55), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(KEYINPUT113), .A3(new_n710), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n854), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT113), .B1(new_n855), .B2(new_n710), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n249), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n241), .A2(new_n242), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n237), .B1(new_n232), .B2(new_n236), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n752), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n752), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n862), .A2(new_n868), .A3(new_n646), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n711), .A2(new_n752), .A3(new_n866), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n754), .B2(new_n862), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n874), .B2(new_n646), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n739), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n713), .A2(new_n755), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n556), .A3(new_n734), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n802), .A2(new_n589), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT115), .Z(new_n882));
  OAI21_X1  g681(.A(G113gat), .B1(new_n882), .B2(new_n258), .ZN(new_n883));
  INV_X1    g682(.A(new_n877), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n875), .B2(new_n739), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n544), .ZN(new_n886));
  INV_X1    g685(.A(new_n476), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n802), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n416), .A2(new_n417), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(new_n754), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n883), .A2(new_n892), .ZN(G1340gat));
  OAI21_X1  g692(.A(G120gat), .B1(new_n882), .B2(new_n712), .ZN(new_n894));
  INV_X1    g693(.A(new_n890), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n711), .A2(new_n415), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT116), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(G1341gat));
  OAI21_X1  g697(.A(new_n408), .B1(new_n895), .B2(new_n739), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n690), .A2(G127gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n882), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT117), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n899), .B(new_n903), .C1(new_n882), .C2(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1342gat));
  OAI21_X1  g704(.A(G134gat), .B1(new_n882), .B2(new_n647), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n833), .A2(new_n647), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n886), .A2(new_n406), .A3(new_n887), .A4(new_n907), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT56), .Z(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n909), .ZN(G1343gat));
  NAND4_X1  g709(.A1(new_n878), .A2(new_n589), .A3(new_n843), .A4(new_n729), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n802), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(G141gat), .A3(new_n258), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(KEYINPUT58), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n350), .B1(new_n876), .B2(new_n877), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(KEYINPUT57), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  OAI211_X1 g718(.A(KEYINPUT118), .B(new_n919), .C1(new_n885), .C2(new_n350), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n257), .A2(new_n710), .A3(new_n855), .A4(new_n859), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n646), .B1(new_n921), .B2(new_n872), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n690), .B1(new_n924), .B2(new_n871), .ZN(new_n925));
  OAI211_X1 g724(.A(KEYINPUT57), .B(new_n733), .C1(new_n925), .C2(new_n884), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n918), .A2(new_n920), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n880), .A2(new_n728), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G141gat), .B1(new_n929), .B2(new_n258), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n754), .A3(new_n928), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n932), .A2(new_n933), .A3(G141gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n932), .B2(G141gat), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n934), .A2(new_n935), .A3(new_n914), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(G1344gat));
  INV_X1    g737(.A(new_n929), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT59), .B(new_n260), .C1(new_n939), .C2(new_n711), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT57), .B1(new_n885), .B2(new_n350), .ZN(new_n942));
  INV_X1    g741(.A(new_n922), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n690), .B1(new_n943), .B2(new_n871), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n713), .A2(new_n258), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n919), .B(new_n733), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n711), .A3(new_n928), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n941), .B1(new_n948), .B2(G148gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n711), .A2(new_n260), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n940), .A2(new_n949), .B1(new_n913), .B2(new_n950), .ZN(G1345gat));
  OAI21_X1  g750(.A(new_n272), .B1(new_n913), .B2(new_n739), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n690), .A2(G155gat), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT121), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n929), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT122), .Z(G1346gat));
  OAI21_X1  g755(.A(G162gat), .B1(new_n929), .B2(new_n647), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n912), .A2(new_n273), .A3(new_n907), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n718), .A2(new_n589), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n879), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(G169gat), .B1(new_n963), .B2(new_n258), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n878), .A2(new_n544), .A3(new_n889), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n476), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n352), .A3(new_n754), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n964), .A2(new_n967), .ZN(G1348gat));
  AOI21_X1  g767(.A(G176gat), .B1(new_n966), .B2(new_n711), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n963), .A2(new_n712), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(G176gat), .ZN(G1349gat));
  AOI21_X1  g770(.A(new_n360), .B1(new_n962), .B2(new_n690), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n739), .A2(new_n361), .A3(new_n363), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n966), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n974), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT60), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n976), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n978));
  AOI22_X1  g777(.A1(new_n975), .A2(new_n977), .B1(new_n974), .B2(new_n978), .ZN(G1350gat));
  AOI21_X1  g778(.A(new_n369), .B1(new_n962), .B2(new_n646), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT61), .Z(new_n981));
  NAND3_X1  g780(.A1(new_n966), .A2(new_n369), .A3(new_n646), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1351gat));
  NOR2_X1   g782(.A1(new_n728), .A2(new_n961), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n984), .B(new_n946), .C1(new_n917), .C2(new_n919), .ZN(new_n985));
  OR3_X1    g784(.A1(new_n985), .A2(KEYINPUT125), .A3(new_n258), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT125), .B1(new_n985), .B2(new_n258), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(G197gat), .A3(new_n987), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n965), .A2(new_n350), .A3(new_n728), .ZN(new_n989));
  INV_X1    g788(.A(G197gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(new_n990), .A3(new_n754), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT126), .ZN(G1352gat));
  INV_X1    g792(.A(G204gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n989), .A2(new_n994), .A3(new_n711), .ZN(new_n995));
  XOR2_X1   g794(.A(new_n995), .B(KEYINPUT62), .Z(new_n996));
  INV_X1    g795(.A(new_n985), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n997), .A2(KEYINPUT127), .A3(new_n711), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n999), .B1(new_n985), .B2(new_n712), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n998), .A2(G204gat), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n996), .A2(new_n1001), .ZN(G1353gat));
  NAND3_X1  g801(.A1(new_n989), .A2(new_n680), .A3(new_n690), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n997), .A2(new_n690), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  INV_X1    g806(.A(G218gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n989), .A2(new_n1008), .A3(new_n646), .ZN(new_n1009));
  OAI21_X1  g808(.A(G218gat), .B1(new_n985), .B2(new_n647), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1355gat));
endmodule


