

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776;

  BUF_X1 U377 ( .A(G119), .Z(n353) );
  INV_X1 U378 ( .A(KEYINPUT72), .ZN(n447) );
  XNOR2_X2 U379 ( .A(n628), .B(n560), .ZN(n616) );
  XNOR2_X2 U380 ( .A(n763), .B(G146), .ZN(n487) );
  INV_X2 U381 ( .A(G953), .ZN(n561) );
  AND2_X2 U382 ( .A1(n408), .A2(KEYINPUT64), .ZN(n368) );
  AND2_X2 U383 ( .A1(n442), .A2(n440), .ZN(n439) );
  NAND2_X2 U384 ( .A1(n410), .A2(n414), .ZN(n369) );
  XNOR2_X2 U385 ( .A(n497), .B(n496), .ZN(n371) );
  XNOR2_X2 U386 ( .A(n447), .B(G131), .ZN(n516) );
  NOR2_X1 U387 ( .A1(n729), .A2(n619), .ZN(n614) );
  AND2_X1 U388 ( .A1(n431), .A2(n429), .ZN(n428) );
  INV_X1 U389 ( .A(n595), .ZN(n584) );
  INV_X1 U390 ( .A(KEYINPUT48), .ZN(n373) );
  AND2_X1 U391 ( .A1(n423), .A2(n420), .ZN(n409) );
  OR2_X1 U392 ( .A1(n748), .A2(n768), .ZN(n356) );
  XNOR2_X1 U393 ( .A(n374), .B(n373), .ZN(n637) );
  NAND2_X1 U394 ( .A1(n428), .A2(n424), .ZN(n354) );
  NOR2_X1 U395 ( .A1(n622), .A2(n605), .ZN(n515) );
  NOR2_X1 U396 ( .A1(n597), .A2(n551), .ZN(n494) );
  OR2_X1 U397 ( .A1(n583), .A2(n582), .ZN(n698) );
  XNOR2_X2 U398 ( .A(n550), .B(n549), .ZN(n577) );
  XNOR2_X1 U399 ( .A(n531), .B(n530), .ZN(n583) );
  XNOR2_X1 U400 ( .A(n449), .B(n538), .ZN(n763) );
  XNOR2_X1 U401 ( .A(n516), .B(n448), .ZN(n449) );
  XNOR2_X1 U402 ( .A(n505), .B(G134), .ZN(n538) );
  XNOR2_X1 U403 ( .A(KEYINPUT16), .B(G122), .ZN(n496) );
  NAND2_X1 U404 ( .A1(n354), .A2(n776), .ZN(n591) );
  XNOR2_X1 U405 ( .A(n354), .B(G110), .ZN(G12) );
  XNOR2_X1 U406 ( .A(n754), .B(n508), .ZN(n355) );
  BUF_X1 U407 ( .A(n774), .Z(n357) );
  INV_X1 U408 ( .A(n594), .ZN(n358) );
  XNOR2_X2 U409 ( .A(n580), .B(n579), .ZN(n703) );
  BUF_X1 U410 ( .A(n581), .Z(n601) );
  XNOR2_X2 U411 ( .A(n402), .B(n419), .ZN(n748) );
  NOR2_X1 U412 ( .A1(n619), .A2(n384), .ZN(n380) );
  NAND2_X1 U413 ( .A1(n617), .A2(n385), .ZN(n384) );
  NAND2_X1 U414 ( .A1(n383), .A2(KEYINPUT47), .ZN(n381) );
  NAND2_X1 U415 ( .A1(n617), .A2(n620), .ZN(n383) );
  XNOR2_X1 U416 ( .A(G146), .B(G125), .ZN(n504) );
  INV_X1 U417 ( .A(KEYINPUT65), .ZN(n432) );
  AND2_X1 U418 ( .A1(n436), .A2(n391), .ZN(n435) );
  OR2_X1 U419 ( .A1(n574), .A2(KEYINPUT65), .ZN(n436) );
  AND2_X1 U420 ( .A1(n640), .A2(n421), .ZN(n420) );
  NAND2_X1 U421 ( .A1(n509), .A2(n422), .ZN(n421) );
  NOR2_X1 U422 ( .A1(n775), .A2(n615), .ZN(n378) );
  NOR2_X1 U423 ( .A1(n626), .A2(n681), .ZN(n627) );
  NAND2_X1 U424 ( .A1(n362), .A2(n379), .ZN(n626) );
  INV_X1 U425 ( .A(KEYINPUT8), .ZN(n462) );
  INV_X1 U426 ( .A(G237), .ZN(n457) );
  NOR2_X1 U427 ( .A1(G953), .A2(G237), .ZN(n522) );
  INV_X1 U428 ( .A(KEYINPUT86), .ZN(n394) );
  XNOR2_X1 U429 ( .A(G143), .B(G104), .ZN(n518) );
  NAND2_X1 U430 ( .A1(n513), .A2(n638), .ZN(n444) );
  NAND2_X1 U431 ( .A1(n391), .A2(n389), .ZN(n608) );
  AND2_X1 U432 ( .A1(n708), .A2(n390), .ZN(n389) );
  INV_X1 U433 ( .A(n551), .ZN(n390) );
  XNOR2_X1 U434 ( .A(n392), .B(n569), .ZN(n581) );
  XNOR2_X1 U435 ( .A(KEYINPUT10), .B(G140), .ZN(n460) );
  XNOR2_X1 U436 ( .A(n387), .B(n386), .ZN(n470) );
  XNOR2_X1 U437 ( .A(G128), .B(G137), .ZN(n386) );
  XNOR2_X1 U438 ( .A(n388), .B(KEYINPUT23), .ZN(n387) );
  XNOR2_X1 U439 ( .A(KEYINPUT81), .B(KEYINPUT24), .ZN(n388) );
  XNOR2_X1 U440 ( .A(n468), .B(n467), .ZN(n540) );
  XNOR2_X1 U441 ( .A(n466), .B(n465), .ZN(n468) );
  INV_X1 U442 ( .A(KEYINPUT71), .ZN(n465) );
  NAND2_X1 U443 ( .A1(n368), .A2(n409), .ZN(n404) );
  XNOR2_X1 U444 ( .A(G110), .B(G107), .ZN(n483) );
  INV_X1 U445 ( .A(G101), .ZN(n482) );
  XOR2_X1 U446 ( .A(G140), .B(KEYINPUT92), .Z(n481) );
  BUF_X1 U447 ( .A(n641), .Z(n694) );
  OR2_X1 U448 ( .A1(n585), .A2(n358), .ZN(n372) );
  AND2_X1 U449 ( .A1(n426), .A2(KEYINPUT103), .ZN(n425) );
  XNOR2_X1 U450 ( .A(n529), .B(n643), .ZN(n530) );
  OR2_X1 U451 ( .A1(n665), .A2(G902), .ZN(n456) );
  XNOR2_X1 U452 ( .A(n609), .B(KEYINPUT6), .ZN(n595) );
  XNOR2_X1 U453 ( .A(G113), .B(G122), .ZN(n517) );
  XOR2_X1 U454 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n519) );
  AND2_X1 U455 ( .A1(n574), .A2(KEYINPUT65), .ZN(n438) );
  NAND2_X1 U456 ( .A1(n377), .A2(n375), .ZN(n374) );
  AND2_X1 U457 ( .A1(n376), .A2(n633), .ZN(n375) );
  XNOR2_X1 U458 ( .A(n378), .B(KEYINPUT46), .ZN(n377) );
  NAND2_X1 U459 ( .A1(n464), .A2(n463), .ZN(n466) );
  INV_X1 U460 ( .A(KEYINPUT82), .ZN(n422) );
  XNOR2_X1 U461 ( .A(G101), .B(KEYINPUT5), .ZN(n450) );
  INV_X1 U462 ( .A(KEYINPUT45), .ZN(n419) );
  XNOR2_X1 U463 ( .A(G116), .B(G122), .ZN(n532) );
  XOR2_X1 U464 ( .A(KEYINPUT100), .B(G107), .Z(n533) );
  XNOR2_X1 U465 ( .A(KEYINPUT102), .B(KEYINPUT7), .ZN(n534) );
  XOR2_X1 U466 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n535) );
  XNOR2_X1 U467 ( .A(n528), .B(n527), .ZN(n644) );
  XNOR2_X1 U468 ( .A(n526), .B(n525), .ZN(n528) );
  INV_X1 U469 ( .A(KEYINPUT33), .ZN(n579) );
  NOR2_X1 U470 ( .A1(n441), .A2(n558), .ZN(n440) );
  NOR2_X1 U471 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U472 ( .A(n370), .B(n761), .ZN(n472) );
  NOR2_X2 U473 ( .A1(n407), .A2(n406), .ZN(n405) );
  NOR2_X1 U474 ( .A1(n409), .A2(KEYINPUT64), .ZN(n407) );
  XNOR2_X1 U475 ( .A(n487), .B(n486), .ZN(n738) );
  XNOR2_X1 U476 ( .A(n648), .B(KEYINPUT88), .ZN(n668) );
  NOR2_X1 U477 ( .A1(n698), .A2(n699), .ZN(n607) );
  XNOR2_X1 U478 ( .A(n372), .B(KEYINPUT78), .ZN(n587) );
  NAND2_X1 U479 ( .A1(n425), .A2(n427), .ZN(n424) );
  NOR2_X1 U480 ( .A1(n586), .A2(n364), .ZN(n401) );
  XNOR2_X1 U481 ( .A(n476), .B(n475), .ZN(n709) );
  AND2_X1 U482 ( .A1(n621), .A2(n603), .ZN(n359) );
  OR2_X1 U483 ( .A1(n774), .A2(KEYINPUT44), .ZN(n360) );
  AND2_X1 U484 ( .A1(n442), .A2(n444), .ZN(n361) );
  AND2_X1 U485 ( .A1(n382), .A2(n381), .ZN(n362) );
  XOR2_X1 U486 ( .A(n624), .B(KEYINPUT76), .Z(n363) );
  OR2_X1 U487 ( .A1(n594), .A2(n595), .ZN(n364) );
  OR2_X1 U488 ( .A1(n601), .A2(KEYINPUT34), .ZN(n365) );
  XOR2_X1 U489 ( .A(n572), .B(KEYINPUT22), .Z(n366) );
  INV_X1 U490 ( .A(KEYINPUT34), .ZN(n416) );
  AND2_X1 U491 ( .A1(n638), .A2(KEYINPUT82), .ZN(n367) );
  XNOR2_X1 U492 ( .A(n589), .B(n588), .ZN(n776) );
  XNOR2_X1 U493 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X2 U494 ( .A(n369), .B(KEYINPUT35), .ZN(n774) );
  NAND2_X1 U495 ( .A1(n540), .A2(G221), .ZN(n370) );
  BUF_X2 U496 ( .A(n433), .Z(n586) );
  NOR2_X2 U497 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X2 U498 ( .A(n371), .B(n498), .ZN(n754) );
  INV_X1 U499 ( .A(n433), .ZN(n575) );
  XNOR2_X2 U500 ( .A(n573), .B(n366), .ZN(n433) );
  NAND2_X1 U501 ( .A1(n616), .A2(n567), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n627), .B(KEYINPUT74), .ZN(n376) );
  NAND2_X1 U503 ( .A1(n621), .A2(n380), .ZN(n379) );
  NAND2_X1 U504 ( .A1(n619), .A2(KEYINPUT47), .ZN(n382) );
  NOR2_X1 U505 ( .A1(n619), .A2(n618), .ZN(n683) );
  INV_X1 U506 ( .A(KEYINPUT47), .ZN(n385) );
  INV_X1 U507 ( .A(n709), .ZN(n391) );
  NOR2_X1 U508 ( .A1(n734), .A2(n643), .ZN(n646) );
  NOR2_X1 U509 ( .A1(n734), .A2(n664), .ZN(n667) );
  NOR2_X1 U510 ( .A1(n734), .A2(n656), .ZN(n660) );
  NAND2_X2 U511 ( .A1(n405), .A2(n403), .ZN(n734) );
  NAND2_X2 U512 ( .A1(n439), .A2(n445), .ZN(n628) );
  NAND2_X1 U513 ( .A1(n397), .A2(n393), .ZN(n402) );
  NAND2_X1 U514 ( .A1(n396), .A2(n604), .ZN(n395) );
  NOR2_X1 U515 ( .A1(n671), .A2(n359), .ZN(n396) );
  NAND2_X1 U516 ( .A1(n399), .A2(n398), .ZN(n397) );
  NAND2_X1 U517 ( .A1(n593), .A2(n592), .ZN(n398) );
  NAND2_X1 U518 ( .A1(n400), .A2(n360), .ZN(n399) );
  INV_X1 U519 ( .A(n593), .ZN(n400) );
  XNOR2_X1 U520 ( .A(n401), .B(KEYINPUT85), .ZN(n596) );
  NAND2_X1 U521 ( .A1(n356), .A2(n422), .ZN(n408) );
  AND2_X2 U522 ( .A1(n642), .A2(n404), .ZN(n403) );
  NOR2_X1 U523 ( .A1(n408), .A2(KEYINPUT64), .ZN(n406) );
  NAND2_X1 U524 ( .A1(n412), .A2(n411), .ZN(n410) );
  NAND2_X1 U525 ( .A1(n703), .A2(n416), .ZN(n411) );
  NAND2_X1 U526 ( .A1(n413), .A2(n365), .ZN(n412) );
  INV_X1 U527 ( .A(n703), .ZN(n413) );
  AND2_X1 U528 ( .A1(n415), .A2(n363), .ZN(n414) );
  NAND2_X1 U529 ( .A1(n601), .A2(KEYINPUT34), .ZN(n415) );
  XNOR2_X2 U530 ( .A(n418), .B(n417), .ZN(n497) );
  XNOR2_X2 U531 ( .A(KEYINPUT3), .B(G119), .ZN(n417) );
  XNOR2_X2 U532 ( .A(G116), .B(G113), .ZN(n418) );
  NAND2_X1 U533 ( .A1(n641), .A2(n367), .ZN(n423) );
  NAND2_X1 U534 ( .A1(n433), .A2(n432), .ZN(n426) );
  INV_X1 U535 ( .A(n434), .ZN(n427) );
  NAND2_X1 U536 ( .A1(n586), .A2(n430), .ZN(n429) );
  AND2_X1 U537 ( .A1(n576), .A2(n432), .ZN(n430) );
  NAND2_X1 U538 ( .A1(n434), .A2(n576), .ZN(n431) );
  NAND2_X1 U539 ( .A1(n437), .A2(n435), .ZN(n434) );
  NAND2_X1 U540 ( .A1(n575), .A2(n438), .ZN(n437) );
  NAND2_X1 U541 ( .A1(n361), .A2(n445), .ZN(n559) );
  INV_X1 U542 ( .A(n444), .ZN(n441) );
  OR2_X2 U543 ( .A1(n657), .A2(n443), .ZN(n442) );
  OR2_X1 U544 ( .A1(n513), .A2(n638), .ZN(n443) );
  NAND2_X1 U545 ( .A1(n355), .A2(n513), .ZN(n445) );
  XNOR2_X1 U546 ( .A(n516), .B(n517), .ZN(n521) );
  NOR2_X2 U547 ( .A1(n581), .A2(n571), .ZN(n573) );
  AND2_X1 U548 ( .A1(G217), .A2(n477), .ZN(n446) );
  INV_X1 U549 ( .A(n761), .ZN(n527) );
  XNOR2_X1 U550 ( .A(KEYINPUT4), .B(G137), .ZN(n448) );
  XNOR2_X2 U551 ( .A(G143), .B(G128), .ZN(n505) );
  NAND2_X1 U552 ( .A1(n522), .A2(G210), .ZN(n451) );
  XNOR2_X1 U553 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U554 ( .A(KEYINPUT75), .B(KEYINPUT96), .ZN(n452) );
  XNOR2_X1 U555 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U556 ( .A(n497), .B(n454), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n487), .B(n455), .ZN(n665) );
  INV_X1 U558 ( .A(G472), .ZN(n664) );
  XNOR2_X2 U559 ( .A(n456), .B(n664), .ZN(n609) );
  INV_X1 U560 ( .A(G902), .ZN(n543) );
  NAND2_X1 U561 ( .A1(n543), .A2(n457), .ZN(n510) );
  AND2_X1 U562 ( .A1(n510), .A2(G214), .ZN(n558) );
  NOR2_X1 U563 ( .A1(n609), .A2(n558), .ZN(n459) );
  XNOR2_X1 U564 ( .A(KEYINPUT106), .B(KEYINPUT30), .ZN(n458) );
  XNOR2_X1 U565 ( .A(n459), .B(n458), .ZN(n495) );
  XNOR2_X1 U566 ( .A(n504), .B(n460), .ZN(n761) );
  INV_X1 U567 ( .A(KEYINPUT70), .ZN(n461) );
  NAND2_X1 U568 ( .A1(n461), .A2(KEYINPUT8), .ZN(n464) );
  NAND2_X1 U569 ( .A1(n462), .A2(KEYINPUT70), .ZN(n463) );
  NAND2_X1 U570 ( .A1(G234), .A2(n561), .ZN(n467) );
  XNOR2_X1 U571 ( .A(n353), .B(G110), .ZN(n469) );
  XNOR2_X1 U572 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n472), .B(n471), .ZN(n652) );
  NAND2_X1 U574 ( .A1(n652), .A2(n543), .ZN(n476) );
  XOR2_X1 U575 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n474) );
  XNOR2_X1 U576 ( .A(G902), .B(KEYINPUT15), .ZN(n509) );
  NAND2_X1 U577 ( .A1(n509), .A2(G234), .ZN(n473) );
  XNOR2_X1 U578 ( .A(n473), .B(KEYINPUT20), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n474), .B(n446), .ZN(n475) );
  AND2_X1 U580 ( .A1(n477), .A2(G221), .ZN(n479) );
  XNOR2_X1 U581 ( .A(KEYINPUT94), .B(KEYINPUT21), .ZN(n478) );
  XNOR2_X1 U582 ( .A(n479), .B(n478), .ZN(n708) );
  NAND2_X1 U583 ( .A1(n709), .A2(n708), .ZN(n706) );
  NAND2_X1 U584 ( .A1(G227), .A2(n561), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n481), .B(n480), .ZN(n485) );
  XNOR2_X1 U586 ( .A(n482), .B(G104), .ZN(n484) );
  XNOR2_X1 U587 ( .A(n484), .B(n483), .ZN(n498) );
  XNOR2_X1 U588 ( .A(n485), .B(n498), .ZN(n486) );
  OR2_X2 U589 ( .A1(n738), .A2(G902), .ZN(n488) );
  INV_X1 U590 ( .A(G469), .ZN(n733) );
  XNOR2_X2 U591 ( .A(n488), .B(n733), .ZN(n550) );
  OR2_X1 U592 ( .A1(n706), .A2(n550), .ZN(n597) );
  NAND2_X1 U593 ( .A1(G237), .A2(G234), .ZN(n490) );
  INV_X1 U594 ( .A(KEYINPUT14), .ZN(n489) );
  XNOR2_X1 U595 ( .A(n490), .B(n489), .ZN(n723) );
  INV_X1 U596 ( .A(n723), .ZN(n565) );
  NOR2_X1 U597 ( .A1(G900), .A2(n561), .ZN(n491) );
  NAND2_X1 U598 ( .A1(n491), .A2(G902), .ZN(n492) );
  NAND2_X1 U599 ( .A1(n561), .A2(G952), .ZN(n563) );
  NAND2_X1 U600 ( .A1(n492), .A2(n563), .ZN(n493) );
  NAND2_X1 U601 ( .A1(n565), .A2(n493), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n495), .A2(n494), .ZN(n622) );
  XNOR2_X1 U603 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n500) );
  XNOR2_X1 U604 ( .A(KEYINPUT18), .B(KEYINPUT89), .ZN(n499) );
  XNOR2_X1 U605 ( .A(n500), .B(n499), .ZN(n503) );
  NAND2_X1 U606 ( .A1(n561), .A2(G224), .ZN(n501) );
  XNOR2_X1 U607 ( .A(n501), .B(KEYINPUT90), .ZN(n502) );
  XNOR2_X1 U608 ( .A(n503), .B(n502), .ZN(n507) );
  XNOR2_X1 U609 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U610 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U611 ( .A(n754), .B(n508), .ZN(n657) );
  INV_X1 U612 ( .A(n509), .ZN(n638) );
  NAND2_X1 U613 ( .A1(n510), .A2(G210), .ZN(n512) );
  INV_X1 U614 ( .A(KEYINPUT79), .ZN(n511) );
  XNOR2_X1 U615 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U616 ( .A(KEYINPUT38), .B(n559), .Z(n605) );
  XNOR2_X1 U617 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n514) );
  XNOR2_X1 U618 ( .A(n515), .B(n514), .ZN(n546) );
  XNOR2_X1 U619 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U620 ( .A(n521), .B(n520), .ZN(n526) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n524) );
  NAND2_X1 U622 ( .A1(G214), .A2(n522), .ZN(n523) );
  XNOR2_X1 U623 ( .A(n524), .B(n523), .ZN(n525) );
  NOR2_X1 U624 ( .A1(G902), .A2(n644), .ZN(n531) );
  XNOR2_X1 U625 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n529) );
  INV_X1 U626 ( .A(G475), .ZN(n643) );
  XNOR2_X1 U627 ( .A(n533), .B(n532), .ZN(n537) );
  XNOR2_X1 U628 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U629 ( .A(n537), .B(n536), .ZN(n539) );
  XNOR2_X1 U630 ( .A(n538), .B(n539), .ZN(n542) );
  NAND2_X1 U631 ( .A1(G217), .A2(n540), .ZN(n541) );
  XNOR2_X1 U632 ( .A(n542), .B(n541), .ZN(n743) );
  NAND2_X1 U633 ( .A1(n743), .A2(n543), .ZN(n544) );
  XNOR2_X1 U634 ( .A(n544), .B(G478), .ZN(n582) );
  INV_X1 U635 ( .A(n582), .ZN(n545) );
  OR2_X1 U636 ( .A1(n583), .A2(n545), .ZN(n690) );
  NOR2_X1 U637 ( .A1(n546), .A2(n690), .ZN(n635) );
  XOR2_X1 U638 ( .A(G134), .B(n635), .Z(G36) );
  NAND2_X1 U639 ( .A1(n583), .A2(n545), .ZN(n686) );
  NOR2_X1 U640 ( .A1(n546), .A2(n686), .ZN(n548) );
  XNOR2_X1 U641 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n547) );
  XNOR2_X1 U642 ( .A(n548), .B(n547), .ZN(n615) );
  XOR2_X1 U643 ( .A(n615), .B(G131), .Z(G33) );
  INV_X1 U644 ( .A(n559), .ZN(n557) );
  XOR2_X1 U645 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n555) );
  INV_X1 U646 ( .A(n558), .ZN(n695) );
  XNOR2_X1 U647 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n549) );
  INV_X1 U648 ( .A(n577), .ZN(n594) );
  NOR2_X1 U649 ( .A1(n686), .A2(n608), .ZN(n552) );
  NAND2_X1 U650 ( .A1(n552), .A2(n595), .ZN(n629) );
  NOR2_X1 U651 ( .A1(n594), .A2(n629), .ZN(n553) );
  NAND2_X1 U652 ( .A1(n695), .A2(n553), .ZN(n554) );
  XOR2_X1 U653 ( .A(n555), .B(n554), .Z(n556) );
  NOR2_X1 U654 ( .A1(n557), .A2(n556), .ZN(n634) );
  XOR2_X1 U655 ( .A(G140), .B(n634), .Z(G42) );
  XNOR2_X1 U656 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n560) );
  NOR2_X1 U657 ( .A1(G898), .A2(n561), .ZN(n562) );
  XOR2_X1 U658 ( .A(KEYINPUT91), .B(n562), .Z(n755) );
  NAND2_X1 U659 ( .A1(n755), .A2(G902), .ZN(n564) );
  NAND2_X1 U660 ( .A1(n564), .A2(n563), .ZN(n566) );
  AND2_X1 U661 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U662 ( .A(KEYINPUT69), .ZN(n568) );
  XNOR2_X1 U663 ( .A(n568), .B(KEYINPUT0), .ZN(n569) );
  INV_X1 U664 ( .A(n698), .ZN(n570) );
  NAND2_X1 U665 ( .A1(n570), .A2(n708), .ZN(n571) );
  INV_X1 U666 ( .A(KEYINPUT73), .ZN(n572) );
  AND2_X1 U667 ( .A1(n609), .A2(n577), .ZN(n574) );
  INV_X1 U668 ( .A(KEYINPUT103), .ZN(n576) );
  NOR2_X2 U669 ( .A1(n577), .A2(n706), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT104), .ZN(n578) );
  NAND2_X1 U671 ( .A1(n578), .A2(n595), .ZN(n580) );
  NAND2_X1 U672 ( .A1(n583), .A2(n582), .ZN(n624) );
  NAND2_X1 U673 ( .A1(n584), .A2(n391), .ZN(n585) );
  XNOR2_X1 U674 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n588) );
  INV_X1 U675 ( .A(KEYINPUT87), .ZN(n590) );
  XNOR2_X1 U676 ( .A(n591), .B(n590), .ZN(n593) );
  INV_X1 U677 ( .A(KEYINPUT44), .ZN(n592) );
  NAND2_X1 U678 ( .A1(n774), .A2(KEYINPUT44), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n596), .A2(n391), .ZN(n671) );
  NAND2_X1 U680 ( .A1(n686), .A2(n690), .ZN(n620) );
  INV_X1 U681 ( .A(n620), .ZN(n700) );
  XOR2_X1 U682 ( .A(n700), .B(KEYINPUT80), .Z(n621) );
  NOR2_X1 U683 ( .A1(n601), .A2(n597), .ZN(n598) );
  XOR2_X1 U684 ( .A(KEYINPUT95), .B(n598), .Z(n599) );
  NAND2_X1 U685 ( .A1(n599), .A2(n609), .ZN(n674) );
  INV_X1 U686 ( .A(n609), .ZN(n711) );
  NAND2_X1 U687 ( .A1(n600), .A2(n711), .ZN(n715) );
  NOR2_X1 U688 ( .A1(n601), .A2(n715), .ZN(n602) );
  XNOR2_X1 U689 ( .A(n602), .B(KEYINPUT31), .ZN(n689) );
  NAND2_X1 U690 ( .A1(n674), .A2(n689), .ZN(n603) );
  INV_X1 U691 ( .A(n605), .ZN(n696) );
  NAND2_X1 U692 ( .A1(n696), .A2(n695), .ZN(n699) );
  XOR2_X1 U693 ( .A(KEYINPUT41), .B(KEYINPUT109), .Z(n606) );
  XNOR2_X1 U694 ( .A(n607), .B(n606), .ZN(n729) );
  XNOR2_X1 U695 ( .A(n610), .B(KEYINPUT28), .ZN(n612) );
  INV_X1 U696 ( .A(n550), .ZN(n611) );
  NAND2_X1 U697 ( .A1(n612), .A2(n611), .ZN(n619) );
  XNOR2_X1 U698 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n613) );
  XNOR2_X1 U699 ( .A(n614), .B(n613), .ZN(n775) );
  BUF_X1 U700 ( .A(n616), .Z(n617) );
  INV_X1 U701 ( .A(n617), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n622), .A2(n559), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n623), .B(KEYINPUT107), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n681) );
  NOR2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n631) );
  XNOR2_X1 U706 ( .A(KEYINPUT111), .B(KEYINPUT36), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X1 U708 ( .A1(n632), .A2(n358), .ZN(n692) );
  XNOR2_X1 U709 ( .A(KEYINPUT83), .B(n692), .ZN(n633) );
  NOR2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n768) );
  NOR2_X2 U712 ( .A1(n748), .A2(n768), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n638), .A2(KEYINPUT2), .ZN(n639) );
  XOR2_X1 U714 ( .A(KEYINPUT67), .B(n639), .Z(n640) );
  NAND2_X1 U715 ( .A1(n694), .A2(KEYINPUT2), .ZN(n642) );
  XOR2_X1 U716 ( .A(n644), .B(KEYINPUT59), .Z(n645) );
  XNOR2_X1 U717 ( .A(n646), .B(n645), .ZN(n649) );
  INV_X1 U718 ( .A(G952), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n647), .A2(G953), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n649), .A2(n668), .ZN(n651) );
  INV_X1 U721 ( .A(KEYINPUT60), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(G60) );
  INV_X1 U723 ( .A(n734), .ZN(n742) );
  NAND2_X1 U724 ( .A1(n742), .A2(G217), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n652), .B(KEYINPUT119), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(n655) );
  INV_X1 U727 ( .A(n668), .ZN(n746) );
  NOR2_X1 U728 ( .A1(n655), .A2(n746), .ZN(G66) );
  INV_X1 U729 ( .A(G210), .ZN(n656) );
  XOR2_X1 U730 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n658) );
  XNOR2_X1 U731 ( .A(n355), .B(n658), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n661), .A2(n668), .ZN(n663) );
  INV_X1 U734 ( .A(KEYINPUT56), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G51) );
  XNOR2_X1 U736 ( .A(n665), .B(KEYINPUT62), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n667), .B(n666), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n670), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U740 ( .A(G101), .B(n671), .Z(G3) );
  NOR2_X1 U741 ( .A1(n674), .A2(n686), .ZN(n672) );
  XOR2_X1 U742 ( .A(KEYINPUT112), .B(n672), .Z(n673) );
  XNOR2_X1 U743 ( .A(G104), .B(n673), .ZN(G6) );
  NOR2_X1 U744 ( .A1(n674), .A2(n690), .ZN(n676) );
  XNOR2_X1 U745 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U747 ( .A(G107), .B(n677), .ZN(G9) );
  XOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .Z(n680) );
  INV_X1 U749 ( .A(n690), .ZN(n678) );
  NAND2_X1 U750 ( .A1(n683), .A2(n678), .ZN(n679) );
  XNOR2_X1 U751 ( .A(n680), .B(n679), .ZN(G30) );
  XOR2_X1 U752 ( .A(G143), .B(n681), .Z(G45) );
  XOR2_X1 U753 ( .A(G146), .B(KEYINPUT113), .Z(n685) );
  INV_X1 U754 ( .A(n686), .ZN(n682) );
  NAND2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n685), .B(n684), .ZN(G48) );
  NOR2_X1 U757 ( .A1(n686), .A2(n689), .ZN(n687) );
  XOR2_X1 U758 ( .A(KEYINPUT114), .B(n687), .Z(n688) );
  XNOR2_X1 U759 ( .A(G113), .B(n688), .ZN(G15) );
  NOR2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U761 ( .A(G116), .B(n691), .Z(G18) );
  XNOR2_X1 U762 ( .A(G125), .B(n692), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U764 ( .A(n694), .B(KEYINPUT2), .ZN(n728) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n705) );
  BUF_X1 U769 ( .A(n703), .Z(n704) );
  NOR2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n358), .A2(n706), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n707), .B(KEYINPUT50), .ZN(n714) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U774 ( .A(KEYINPUT49), .B(n710), .Z(n712) );
  NOR2_X1 U775 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U778 ( .A(KEYINPUT51), .B(n717), .ZN(n718) );
  NOR2_X1 U779 ( .A1(n729), .A2(n718), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U781 ( .A(n721), .B(KEYINPUT52), .ZN(n722) );
  NOR2_X1 U782 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U783 ( .A1(n724), .A2(G952), .ZN(n725) );
  XNOR2_X1 U784 ( .A(KEYINPUT115), .B(n725), .ZN(n726) );
  NOR2_X1 U785 ( .A1(G953), .A2(n726), .ZN(n727) );
  NAND2_X1 U786 ( .A1(n728), .A2(n727), .ZN(n731) );
  NOR2_X1 U787 ( .A1(n729), .A2(n704), .ZN(n730) );
  NOR2_X1 U788 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U789 ( .A(KEYINPUT53), .B(n732), .ZN(G75) );
  NOR2_X1 U790 ( .A1(n734), .A2(n733), .ZN(n740) );
  XOR2_X1 U791 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n736) );
  XNOR2_X1 U792 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n735) );
  XNOR2_X1 U793 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U794 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U795 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U796 ( .A1(n741), .A2(n746), .ZN(G54) );
  NAND2_X1 U797 ( .A1(n742), .A2(G478), .ZN(n745) );
  XOR2_X1 U798 ( .A(KEYINPUT118), .B(n743), .Z(n744) );
  XNOR2_X1 U799 ( .A(n745), .B(n744), .ZN(n747) );
  NOR2_X1 U800 ( .A1(n747), .A2(n746), .ZN(G63) );
  NOR2_X1 U801 ( .A1(n748), .A2(G953), .ZN(n749) );
  XOR2_X1 U802 ( .A(KEYINPUT120), .B(n749), .Z(n753) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n750) );
  XNOR2_X1 U804 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U805 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U806 ( .A1(n753), .A2(n752), .ZN(n760) );
  XNOR2_X1 U807 ( .A(n754), .B(KEYINPUT121), .ZN(n756) );
  NOR2_X1 U808 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U809 ( .A(n757), .B(KEYINPUT122), .Z(n758) );
  XNOR2_X1 U810 ( .A(KEYINPUT123), .B(n758), .ZN(n759) );
  XNOR2_X1 U811 ( .A(n760), .B(n759), .ZN(G69) );
  XNOR2_X1 U812 ( .A(n761), .B(KEYINPUT92), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(n769) );
  XNOR2_X1 U814 ( .A(n769), .B(KEYINPUT124), .ZN(n764) );
  XNOR2_X1 U815 ( .A(G227), .B(n764), .ZN(n765) );
  NAND2_X1 U816 ( .A1(G900), .A2(n765), .ZN(n766) );
  NAND2_X1 U817 ( .A1(G953), .A2(n766), .ZN(n767) );
  XNOR2_X1 U818 ( .A(n767), .B(KEYINPUT125), .ZN(n772) );
  XOR2_X1 U819 ( .A(n769), .B(n768), .Z(n770) );
  NOR2_X1 U820 ( .A1(n770), .A2(G953), .ZN(n771) );
  NOR2_X1 U821 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U822 ( .A(KEYINPUT126), .B(n773), .Z(G72) );
  XOR2_X1 U823 ( .A(n357), .B(G122), .Z(G24) );
  XOR2_X1 U824 ( .A(n775), .B(G137), .Z(G39) );
  XNOR2_X1 U825 ( .A(n776), .B(n353), .ZN(G21) );
endmodule

