

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U555 ( .A1(n815), .A2(n524), .ZN(n817) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n653) );
  AND2_X1 U557 ( .A1(n779), .A2(n522), .ZN(n521) );
  NOR2_X2 U558 ( .A1(G2104), .A2(n542), .ZN(n612) );
  OR2_X1 U559 ( .A1(n778), .A2(n777), .ZN(n522) );
  OR2_X1 U560 ( .A1(n777), .A2(n769), .ZN(n523) );
  AND2_X1 U561 ( .A1(n824), .A2(n526), .ZN(n524) );
  XOR2_X1 U562 ( .A(KEYINPUT78), .B(n585), .Z(n525) );
  OR2_X1 U563 ( .A1(n814), .A2(n813), .ZN(n526) );
  AND2_X1 U564 ( .A1(n696), .A2(n695), .ZN(n699) );
  AND2_X1 U565 ( .A1(n722), .A2(n721), .ZN(n724) );
  AND2_X1 U566 ( .A1(n732), .A2(G171), .ZN(n725) );
  BUF_X1 U567 ( .A(n728), .Z(n739) );
  XNOR2_X1 U568 ( .A(n747), .B(KEYINPUT32), .ZN(n755) );
  INV_X1 U569 ( .A(KEYINPUT106), .ZN(n765) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  NOR2_X2 U571 ( .A1(n633), .A2(n533), .ZN(n658) );
  INV_X1 U572 ( .A(KEYINPUT107), .ZN(n816) );
  NOR2_X1 U573 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U574 ( .A(n817), .B(n816), .ZN(n831) );
  XNOR2_X1 U575 ( .A(n589), .B(KEYINPUT15), .ZN(n1007) );
  NAND2_X1 U576 ( .A1(n581), .A2(n580), .ZN(n1008) );
  XNOR2_X1 U577 ( .A(n549), .B(n548), .ZN(n690) );
  BUF_X1 U578 ( .A(n690), .Z(G160) );
  XNOR2_X1 U579 ( .A(KEYINPUT9), .B(KEYINPUT71), .ZN(n530) );
  NAND2_X1 U580 ( .A1(G90), .A2(n653), .ZN(n528) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n633) );
  INV_X1 U582 ( .A(G651), .ZN(n533) );
  NAND2_X1 U583 ( .A1(G77), .A2(n658), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U585 ( .A(n530), .B(n529), .ZN(n538) );
  NOR2_X1 U586 ( .A1(G651), .A2(n633), .ZN(n531) );
  XOR2_X2 U587 ( .A(KEYINPUT65), .B(n531), .Z(n662) );
  NAND2_X1 U588 ( .A1(n662), .A2(G52), .ZN(n532) );
  XNOR2_X1 U589 ( .A(n532), .B(KEYINPUT70), .ZN(n536) );
  NOR2_X1 U590 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X2 U591 ( .A(KEYINPUT1), .B(n534), .Z(n654) );
  NAND2_X1 U592 ( .A1(G64), .A2(n654), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U594 ( .A1(n538), .A2(n537), .ZN(G171) );
  AND2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n874) );
  NAND2_X1 U596 ( .A1(n874), .A2(G113), .ZN(n547) );
  XOR2_X1 U597 ( .A(KEYINPUT17), .B(n539), .Z(n561) );
  NAND2_X1 U598 ( .A1(G137), .A2(n561), .ZN(n541) );
  INV_X2 U599 ( .A(G2105), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G125), .A2(n612), .ZN(n540) );
  NAND2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n545) );
  AND2_X4 U602 ( .A1(n542), .A2(G2104), .ZN(n878) );
  NAND2_X1 U603 ( .A1(G101), .A2(n878), .ZN(n543) );
  XNOR2_X1 U604 ( .A(KEYINPUT23), .B(n543), .ZN(n544) );
  NOR2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X1 U607 ( .A(KEYINPUT66), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n653), .A2(G89), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G76), .A2(n658), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U612 ( .A(KEYINPUT5), .B(n553), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n654), .A2(G63), .ZN(n554) );
  XOR2_X1 U614 ( .A(KEYINPUT79), .B(n554), .Z(n556) );
  NAND2_X1 U615 ( .A1(n662), .A2(G51), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(KEYINPUT7), .B(n560), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  NAND2_X1 U624 ( .A1(G102), .A2(n878), .ZN(n563) );
  BUF_X1 U625 ( .A(n561), .Z(n616) );
  NAND2_X1 U626 ( .A1(G138), .A2(n616), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G114), .A2(n874), .ZN(n565) );
  NAND2_X1 U629 ( .A1(G126), .A2(n612), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT89), .B(n566), .Z(n567) );
  NOR2_X1 U632 ( .A1(n568), .A2(n567), .ZN(G164) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U635 ( .A(G223), .ZN(n833) );
  NAND2_X1 U636 ( .A1(n833), .A2(G567), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  INV_X1 U638 ( .A(G860), .ZN(n603) );
  NAND2_X1 U639 ( .A1(n653), .A2(G81), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U641 ( .A1(G68), .A2(n658), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT76), .B(KEYINPUT13), .Z(n574) );
  XNOR2_X1 U644 ( .A(n575), .B(n574), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G56), .A2(n654), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT14), .ZN(n577) );
  XNOR2_X1 U647 ( .A(KEYINPUT75), .B(n577), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n662), .A2(G43), .ZN(n580) );
  NOR2_X1 U649 ( .A1(n603), .A2(n1008), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n582), .B(KEYINPUT77), .ZN(G153) );
  INV_X1 U651 ( .A(G171), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G54), .A2(n662), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G92), .A2(n653), .ZN(n584) );
  NAND2_X1 U655 ( .A1(G66), .A2(n654), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n658), .A2(G79), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n586), .A2(n525), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n589) );
  OR2_X1 U660 ( .A1(n1007), .A2(G868), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U662 ( .A1(G78), .A2(n658), .ZN(n592) );
  XOR2_X1 U663 ( .A(KEYINPUT72), .B(n592), .Z(n597) );
  NAND2_X1 U664 ( .A1(G65), .A2(n654), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G53), .A2(n662), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U667 ( .A(KEYINPUT73), .B(n595), .Z(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n653), .A2(G91), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(G299) );
  INV_X1 U671 ( .A(G868), .ZN(n600) );
  NOR2_X1 U672 ( .A1(G286), .A2(n600), .ZN(n602) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U674 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n604), .A2(n1007), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n1008), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G868), .A2(n1007), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G99), .A2(n878), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G111), .A2(n874), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U685 ( .A(KEYINPUT80), .B(n611), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n612), .A2(G123), .ZN(n613) );
  XOR2_X1 U687 ( .A(KEYINPUT18), .B(n613), .Z(n614) );
  NOR2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n616), .A2(G135), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n928) );
  XNOR2_X1 U691 ( .A(G2096), .B(n928), .ZN(n619) );
  NOR2_X1 U692 ( .A1(n619), .A2(G2100), .ZN(n620) );
  XNOR2_X1 U693 ( .A(n620), .B(KEYINPUT81), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G67), .A2(n654), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G55), .A2(n662), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G93), .A2(n653), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G80), .A2(n658), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n672) );
  NAND2_X1 U701 ( .A1(G559), .A2(n1007), .ZN(n627) );
  XOR2_X1 U702 ( .A(n1008), .B(n627), .Z(n670) );
  XOR2_X1 U703 ( .A(n670), .B(KEYINPUT82), .Z(n628) );
  NOR2_X1 U704 ( .A1(G860), .A2(n628), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n672), .B(n629), .ZN(G145) );
  NAND2_X1 U706 ( .A1(G49), .A2(n662), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n654), .A2(n632), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G87), .A2(n633), .ZN(n634) );
  XOR2_X1 U711 ( .A(KEYINPUT83), .B(n634), .Z(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G75), .A2(n658), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G62), .A2(n654), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G88), .A2(n653), .ZN(n639) );
  XNOR2_X1 U717 ( .A(KEYINPUT85), .B(n639), .ZN(n640) );
  NOR2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n662), .A2(G50), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n643), .A2(n642), .ZN(G303) );
  INV_X1 U721 ( .A(G303), .ZN(G166) );
  NAND2_X1 U722 ( .A1(n653), .A2(G85), .ZN(n644) );
  XOR2_X1 U723 ( .A(KEYINPUT67), .B(n644), .Z(n646) );
  NAND2_X1 U724 ( .A1(n658), .A2(G72), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U726 ( .A(KEYINPUT68), .B(n647), .ZN(n650) );
  NAND2_X1 U727 ( .A1(G60), .A2(n654), .ZN(n648) );
  XNOR2_X1 U728 ( .A(KEYINPUT69), .B(n648), .ZN(n649) );
  NOR2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n662), .A2(G47), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n652), .A2(n651), .ZN(G290) );
  NAND2_X1 U732 ( .A1(G86), .A2(n653), .ZN(n656) );
  NAND2_X1 U733 ( .A1(G61), .A2(n654), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U735 ( .A(KEYINPUT84), .B(n657), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n658), .A2(G73), .ZN(n659) );
  XOR2_X1 U737 ( .A(KEYINPUT2), .B(n659), .Z(n660) );
  NOR2_X1 U738 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U739 ( .A1(n662), .A2(G48), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n664), .A2(n663), .ZN(G305) );
  XNOR2_X1 U741 ( .A(KEYINPUT19), .B(G288), .ZN(n669) );
  XNOR2_X1 U742 ( .A(G166), .B(n672), .ZN(n667) );
  XNOR2_X1 U743 ( .A(G290), .B(G299), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n665), .B(G305), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n669), .B(n668), .ZN(n904) );
  XNOR2_X1 U747 ( .A(n670), .B(n904), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n671), .A2(G868), .ZN(n674) );
  OR2_X1 U749 ( .A1(G868), .A2(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n675) );
  XNOR2_X1 U753 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U756 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XOR2_X1 U757 ( .A(KEYINPUT74), .B(G132), .Z(G219) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G219), .A2(G220), .ZN(n680) );
  XNOR2_X1 U760 ( .A(KEYINPUT22), .B(n680), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n681), .A2(G96), .ZN(n682) );
  NOR2_X1 U762 ( .A1(n682), .A2(G218), .ZN(n683) );
  XNOR2_X1 U763 ( .A(n683), .B(KEYINPUT87), .ZN(n838) );
  NAND2_X1 U764 ( .A1(n838), .A2(G2106), .ZN(n688) );
  NAND2_X1 U765 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U766 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U767 ( .A1(G108), .A2(n685), .ZN(n837) );
  NAND2_X1 U768 ( .A1(G567), .A2(n837), .ZN(n686) );
  XNOR2_X1 U769 ( .A(KEYINPUT88), .B(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(n688), .A2(n687), .ZN(n839) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U772 ( .A1(n839), .A2(n689), .ZN(n836) );
  NAND2_X1 U773 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U774 ( .A1(n690), .A2(G40), .ZN(n692) );
  INV_X1 U775 ( .A(KEYINPUT90), .ZN(n691) );
  XNOR2_X2 U776 ( .A(n692), .B(n691), .ZN(n783) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n781) );
  NAND2_X1 U778 ( .A1(n783), .A2(n781), .ZN(n728) );
  INV_X1 U779 ( .A(n728), .ZN(n720) );
  NAND2_X1 U780 ( .A1(n720), .A2(G1996), .ZN(n693) );
  XNOR2_X1 U781 ( .A(n693), .B(KEYINPUT26), .ZN(n696) );
  AND2_X1 U782 ( .A1(n739), .A2(G1341), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n694), .A2(n1008), .ZN(n695) );
  INV_X1 U784 ( .A(n699), .ZN(n698) );
  INV_X1 U785 ( .A(n1007), .ZN(n697) );
  NAND2_X1 U786 ( .A1(n698), .A2(n697), .ZN(n706) );
  NAND2_X1 U787 ( .A1(n1007), .A2(n699), .ZN(n704) );
  AND2_X1 U788 ( .A1(n720), .A2(G2067), .ZN(n700) );
  XOR2_X1 U789 ( .A(n700), .B(KEYINPUT102), .Z(n702) );
  NAND2_X1 U790 ( .A1(n739), .A2(G1348), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U792 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U793 ( .A1(n706), .A2(n705), .ZN(n712) );
  INV_X1 U794 ( .A(G299), .ZN(n997) );
  NAND2_X1 U795 ( .A1(n720), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U796 ( .A(KEYINPUT27), .B(n707), .ZN(n710) );
  AND2_X1 U797 ( .A1(G1956), .A2(n728), .ZN(n708) );
  XNOR2_X1 U798 ( .A(KEYINPUT100), .B(n708), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U800 ( .A1(n997), .A2(n713), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U802 ( .A1(n713), .A2(n997), .ZN(n715) );
  XNOR2_X1 U803 ( .A(KEYINPUT101), .B(KEYINPUT28), .ZN(n714) );
  XNOR2_X1 U804 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U806 ( .A(n718), .B(KEYINPUT29), .ZN(n727) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n954) );
  NOR2_X1 U808 ( .A1(n954), .A2(n728), .ZN(n719) );
  XNOR2_X1 U809 ( .A(n719), .B(KEYINPUT97), .ZN(n722) );
  OR2_X1 U810 ( .A1(n720), .A2(G1961), .ZN(n721) );
  INV_X1 U811 ( .A(KEYINPUT98), .ZN(n723) );
  XNOR2_X1 U812 ( .A(n724), .B(n723), .ZN(n732) );
  XOR2_X1 U813 ( .A(KEYINPUT99), .B(n725), .Z(n726) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n737) );
  NAND2_X1 U815 ( .A1(G8), .A2(n728), .ZN(n777) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n777), .ZN(n751) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n739), .ZN(n748) );
  NOR2_X1 U818 ( .A1(n751), .A2(n748), .ZN(n729) );
  NAND2_X1 U819 ( .A1(G8), .A2(n729), .ZN(n730) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U821 ( .A1(G168), .A2(n731), .ZN(n734) );
  NOR2_X1 U822 ( .A1(G171), .A2(n732), .ZN(n733) );
  NOR2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n735), .B(KEYINPUT31), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U826 ( .A(n738), .B(KEYINPUT103), .ZN(n749) );
  NAND2_X1 U827 ( .A1(n749), .A2(G286), .ZN(n745) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n739), .ZN(n740) );
  XNOR2_X1 U829 ( .A(n740), .B(KEYINPUT104), .ZN(n742) );
  NOR2_X1 U830 ( .A1(n777), .A2(G1971), .ZN(n741) );
  NOR2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n743), .A2(G303), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n746), .A2(G8), .ZN(n747) );
  NAND2_X1 U835 ( .A1(G8), .A2(n748), .ZN(n753) );
  INV_X1 U836 ( .A(n749), .ZN(n750) );
  NOR2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n755), .A2(n754), .ZN(n771) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n756) );
  XNOR2_X1 U841 ( .A(KEYINPUT105), .B(n756), .ZN(n757) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n768) );
  INV_X1 U843 ( .A(n768), .ZN(n1006) );
  AND2_X1 U844 ( .A1(n757), .A2(n1006), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n771), .A2(n758), .ZN(n761) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n1005) );
  INV_X1 U847 ( .A(n777), .ZN(n759) );
  AND2_X1 U848 ( .A1(n1005), .A2(n759), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n763) );
  INV_X1 U850 ( .A(KEYINPUT64), .ZN(n762) );
  XNOR2_X1 U851 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X2 U852 ( .A1(n764), .A2(KEYINPUT33), .ZN(n766) );
  XNOR2_X1 U853 ( .A(n766), .B(n765), .ZN(n767) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n1002) );
  AND2_X1 U855 ( .A1(n767), .A2(n1002), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n768), .A2(KEYINPUT33), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n523), .ZN(n780) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n771), .A2(n773), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n774), .A2(n777), .ZN(n779) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U863 ( .A(n775), .B(KEYINPUT96), .Z(n776) );
  XNOR2_X1 U864 ( .A(KEYINPUT24), .B(n776), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n780), .A2(n521), .ZN(n815) );
  INV_X1 U866 ( .A(n781), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n813) );
  INV_X1 U868 ( .A(n813), .ZN(n828) );
  NAND2_X1 U869 ( .A1(n616), .A2(G140), .ZN(n784) );
  XOR2_X1 U870 ( .A(KEYINPUT91), .B(n784), .Z(n786) );
  NAND2_X1 U871 ( .A1(n878), .A2(G104), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U873 ( .A(KEYINPUT34), .B(n787), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G116), .A2(n874), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G128), .A2(n612), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U877 ( .A(n790), .B(KEYINPUT35), .Z(n791) );
  NOR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U879 ( .A(KEYINPUT36), .B(n793), .Z(n794) );
  XOR2_X1 U880 ( .A(KEYINPUT92), .B(n794), .Z(n899) );
  XNOR2_X1 U881 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U882 ( .A1(n899), .A2(n826), .ZN(n944) );
  NAND2_X1 U883 ( .A1(n828), .A2(n944), .ZN(n824) );
  NAND2_X1 U884 ( .A1(G117), .A2(n874), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G129), .A2(n612), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U887 ( .A1(n878), .A2(G105), .ZN(n797) );
  XOR2_X1 U888 ( .A(KEYINPUT38), .B(n797), .Z(n798) );
  NOR2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n616), .A2(G141), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n888) );
  NAND2_X1 U892 ( .A1(G1996), .A2(n888), .ZN(n812) );
  NAND2_X1 U893 ( .A1(G95), .A2(n878), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G131), .A2(n616), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n809) );
  NAND2_X1 U896 ( .A1(n874), .A2(G107), .ZN(n804) );
  XOR2_X1 U897 ( .A(KEYINPUT93), .B(n804), .Z(n806) );
  NAND2_X1 U898 ( .A1(n612), .A2(G119), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U900 ( .A(KEYINPUT94), .B(n807), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U902 ( .A(n810), .B(KEYINPUT95), .ZN(n896) );
  NAND2_X1 U903 ( .A1(G1991), .A2(n896), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n927) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n999) );
  NOR2_X1 U906 ( .A1(n927), .A2(n999), .ZN(n814) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n888), .ZN(n924) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n896), .ZN(n931) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n818) );
  XNOR2_X1 U910 ( .A(KEYINPUT108), .B(n818), .ZN(n819) );
  NOR2_X1 U911 ( .A1(n931), .A2(n819), .ZN(n820) );
  NOR2_X1 U912 ( .A1(n820), .A2(n927), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n924), .A2(n821), .ZN(n822) );
  XOR2_X1 U914 ( .A(n822), .B(KEYINPUT39), .Z(n823) );
  XNOR2_X1 U915 ( .A(KEYINPUT109), .B(n823), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n899), .A2(n826), .ZN(n932) );
  NAND2_X1 U918 ( .A1(n827), .A2(n932), .ZN(n829) );
  NAND2_X1 U919 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U920 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U921 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U924 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n839), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n841) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n843) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U940 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1981), .B(G1971), .Z(n849) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1956), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U946 ( .A(n850), .B(KEYINPUT41), .Z(n852) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U949 ( .A(G2474), .B(G1976), .Z(n854) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1961), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U953 ( .A1(G100), .A2(n878), .ZN(n858) );
  NAND2_X1 U954 ( .A1(G112), .A2(n874), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n859), .B(KEYINPUT111), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G136), .A2(n616), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U959 ( .A1(n612), .A2(G124), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT44), .B(n862), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U962 ( .A1(G103), .A2(n878), .ZN(n866) );
  NAND2_X1 U963 ( .A1(G139), .A2(n616), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U965 ( .A1(n874), .A2(G115), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n867), .B(KEYINPUT114), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G127), .A2(n612), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n870), .Z(n871) );
  NOR2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n934) );
  XOR2_X1 U971 ( .A(G164), .B(n934), .Z(n873) );
  XNOR2_X1 U972 ( .A(n928), .B(n873), .ZN(n895) );
  NAND2_X1 U973 ( .A1(n874), .A2(G118), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(KEYINPUT112), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G130), .A2(n612), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n884) );
  XNOR2_X1 U977 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G106), .A2(n878), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G142), .A2(n616), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n893) );
  XOR2_X1 U983 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n886) );
  XNOR2_X1 U984 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(KEYINPUT117), .B(n887), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n888), .B(KEYINPUT118), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U989 ( .A(G160), .B(n891), .Z(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n896), .B(G162), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U995 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n1008), .B(G286), .ZN(n903) );
  XNOR2_X1 U997 ( .A(G171), .B(n1007), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U1001 ( .A(G2451), .B(G2443), .Z(n908) );
  XNOR2_X1 U1002 ( .A(G2427), .B(G2454), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1004 ( .A(n909), .B(G2446), .Z(n911) );
  XNOR2_X1 U1005 ( .A(G1341), .B(G1348), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1007 ( .A(G2435), .B(KEYINPUT110), .Z(n913) );
  XNOR2_X1 U1008 ( .A(G2430), .B(G2438), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1010 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1011 ( .A1(G14), .A2(n916), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  INV_X1 U1020 ( .A(n922), .ZN(G401) );
  INV_X1 U1021 ( .A(KEYINPUT55), .ZN(n969) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n925), .B(KEYINPUT51), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n942) );
  XNOR2_X1 U1026 ( .A(G160), .B(G2084), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(G2072), .B(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(G164), .B(G2078), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1033 ( .A(KEYINPUT119), .B(n937), .Z(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT50), .B(n938), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n969), .A2(n946), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n1024) );
  XOR2_X1 U1041 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n962) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G2072), .B(G33), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1045 ( .A(KEYINPUT121), .B(n950), .Z(n953) );
  XOR2_X1 U1046 ( .A(KEYINPUT120), .B(G25), .Z(n951) );
  XNOR2_X1 U1047 ( .A(G1991), .B(n951), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(G1996), .B(G32), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n954), .B(G27), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1052 ( .A(KEYINPUT122), .B(n957), .Z(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n960), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n962), .B(n961), .ZN(n968) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(KEYINPUT124), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n963), .B(G34), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(G2084), .B(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(G2090), .B(G35), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n1025) );
  OR2_X1 U1062 ( .A1(n969), .A2(n1025), .ZN(n996) );
  XNOR2_X1 U1063 ( .A(KEYINPUT125), .B(G1961), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n970), .B(G5), .ZN(n989) );
  XNOR2_X1 U1065 ( .A(G1341), .B(G19), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G6), .B(G1981), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n978) );
  XOR2_X1 U1068 ( .A(G4), .B(KEYINPUT126), .Z(n974) );
  XNOR2_X1 U1069 ( .A(G1348), .B(KEYINPUT59), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(n974), .B(n973), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(G1956), .B(G20), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n979), .B(KEYINPUT60), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(G23), .B(G1976), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(G1986), .B(KEYINPUT127), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(n982), .B(G24), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(KEYINPUT58), .B(n985), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(G21), .B(G1966), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT61), .B(n992), .ZN(n994) );
  INV_X1 U1087 ( .A(G16), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n1022) );
  XOR2_X1 U1090 ( .A(KEYINPUT56), .B(G16), .Z(n1020) );
  XNOR2_X1 U1091 ( .A(n997), .B(G1956), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(G1961), .B(G301), .ZN(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1018) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G168), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1097 ( .A(n1004), .B(KEYINPUT57), .ZN(n1016) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1007), .B(G1348), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1008), .B(G1341), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(G303), .B(G1971), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1029) );
  NOR2_X1 U1110 ( .A1(KEYINPUT55), .A2(G29), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(G11), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1114 ( .A(n1030), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

