//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT66), .Z(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  AND3_X1   g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n209), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n208), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(G58), .A2(G68), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n222), .A2(G50), .A3(new_n223), .ZN(new_n224));
  OAI22_X1  g0024(.A1(new_n216), .A2(new_n217), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n209), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT64), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n225), .B(new_n231), .C1(new_n217), .C2(new_n216), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n236), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  INV_X1    g0046(.A(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT72), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(KEYINPUT10), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n208), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n255), .A2(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n260), .B1(G20), .B2(new_n204), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n262), .A2(new_n218), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n226), .A2(new_n208), .A3(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n201), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(G1), .B2(new_n208), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(new_n201), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n266), .B1(new_n201), .B2(new_n267), .C1(new_n261), .C2(new_n263), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT9), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G223), .A2(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n218), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n280), .B(new_n282), .C1(G77), .C2(new_n276), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT69), .B(G45), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n207), .B(G274), .C1(new_n284), .C2(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G226), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n207), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n283), .B(new_n285), .C1(new_n286), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G200), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n270), .A2(new_n273), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT71), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n254), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n253), .A2(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n297), .A2(new_n300), .A3(new_n253), .A4(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n271), .C1(G179), .C2(new_n295), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n255), .A2(new_n265), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n267), .B2(new_n255), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT77), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(KEYINPUT77), .B(new_n310), .C1(new_n267), .C2(new_n255), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT7), .B1(new_n318), .B2(new_n208), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  NOR4_X1   g0120(.A1(new_n316), .A2(new_n317), .A3(new_n320), .A4(G20), .ZN(new_n321));
  OAI21_X1  g0121(.A(G68), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n202), .A2(new_n203), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n323), .B2(new_n221), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n258), .A2(G159), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT16), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n263), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n322), .A2(KEYINPUT16), .A3(new_n327), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n315), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  INV_X1    g0133(.A(G33), .ZN(new_n334));
  INV_X1    g0134(.A(G87), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G223), .A2(G1698), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n286), .B2(G1698), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n336), .B1(new_n338), .B2(new_n276), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n285), .B1(new_n339), .B2(new_n293), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n240), .B(new_n282), .C1(new_n290), .C2(new_n289), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n333), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n286), .A2(G1698), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G223), .B2(G1698), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n344), .A2(new_n318), .B1(new_n334), .B2(new_n335), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n282), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G232), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n346), .A2(new_n348), .A3(new_n298), .A4(new_n285), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n342), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT78), .B1(new_n332), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n274), .A2(new_n208), .A3(new_n275), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n320), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n318), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n203), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n329), .B1(new_n355), .B2(new_n326), .ZN(new_n356));
  INV_X1    g0156(.A(new_n263), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n331), .A3(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n313), .A2(new_n314), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n350), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT78), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT17), .B1(new_n351), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G169), .B1(new_n340), .B2(new_n341), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n346), .A2(new_n348), .A3(G179), .A4(new_n285), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n358), .A2(new_n359), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT18), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n350), .A2(new_n358), .A3(new_n359), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(KEYINPUT17), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n363), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G238), .A2(G1698), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n276), .B(new_n372), .C1(new_n240), .C2(G1698), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n282), .C1(G107), .C2(new_n276), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n285), .ZN(new_n375));
  INV_X1    g0175(.A(G244), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n294), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G190), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G20), .A2(G77), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT15), .B(G87), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n380), .B1(new_n255), .B2(new_n259), .C1(new_n256), .C2(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n382), .A2(new_n357), .ZN(new_n383));
  INV_X1    g0183(.A(G77), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n265), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n267), .B2(new_n384), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n379), .B(new_n387), .C1(new_n333), .C2(new_n378), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n387), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n390), .B(new_n391), .C1(G169), .C2(new_n378), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n309), .A2(new_n371), .A3(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n265), .A2(KEYINPUT12), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n203), .A2(G20), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n226), .A2(G1), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT12), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n396), .B1(new_n256), .B2(new_n384), .C1(new_n259), .C2(new_n201), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n357), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT11), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n395), .B1(new_n396), .B2(new_n398), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT11), .B1(new_n399), .B2(new_n357), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n203), .B1(new_n267), .B2(KEYINPUT12), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n294), .A2(KEYINPUT73), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n347), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(G238), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n207), .A2(G274), .ZN(new_n412));
  AND2_X1   g0212(.A1(KEYINPUT69), .A2(G45), .ZN(new_n413));
  NOR2_X1   g0213(.A1(KEYINPUT69), .A2(G45), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G41), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n240), .A2(G1698), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G226), .B2(G1698), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n418), .B1(new_n420), .B2(new_n318), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n417), .B1(new_n421), .B2(new_n282), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n407), .B1(new_n411), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(G238), .B1(new_n347), .B2(new_n409), .ZN(new_n424));
  AOI211_X1 g0224(.A(KEYINPUT73), .B(new_n282), .C1(new_n290), .C2(new_n289), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n407), .B(new_n422), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(G169), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n426), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(KEYINPUT14), .A3(G169), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n426), .A2(G179), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n407), .B1(new_n431), .B2(KEYINPUT74), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT74), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n411), .A2(new_n438), .A3(new_n422), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n436), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT76), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  AOI211_X1 g0243(.A(new_n443), .B(new_n440), .C1(new_n430), .C2(new_n434), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n406), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n433), .A2(G200), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n405), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n437), .A2(new_n439), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n427), .A2(new_n298), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(KEYINPUT75), .A3(new_n449), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n394), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(G238), .A2(G1698), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n376), .A2(G1698), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n459), .C1(new_n316), .C2(new_n317), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G116), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n293), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G250), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n207), .B2(G45), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n293), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT81), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n293), .A3(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n293), .A2(G274), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n207), .A2(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n463), .A2(new_n470), .A3(G190), .A4(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n335), .A2(new_n478), .A3(new_n244), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n418), .A2(new_n208), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT19), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n208), .B(G68), .C1(new_n316), .C2(new_n317), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT19), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n256), .B2(new_n478), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(new_n357), .B1(new_n265), .B2(new_n381), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n397), .A2(G20), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n263), .B(new_n487), .C1(G1), .C2(new_n334), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n488), .A2(new_n335), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n463), .A2(new_n470), .A3(new_n474), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G200), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n462), .A2(new_n473), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(KEYINPUT82), .A3(G190), .A4(new_n470), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n477), .A2(new_n490), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n465), .A2(new_n293), .A3(KEYINPUT81), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT81), .B1(new_n465), .B2(new_n293), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n498), .A2(new_n462), .A3(new_n473), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n389), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n491), .A2(new_n305), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n486), .B1(new_n381), .B2(new_n488), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n276), .A2(G250), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n277), .B1(new_n505), .B2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G1698), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(G244), .C1(new_n317), .C2(new_n316), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n376), .B1(new_n274), .B2(new_n275), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n511), .C2(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n282), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT79), .ZN(new_n514));
  INV_X1    g0314(.A(G45), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G1), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G41), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n514), .B1(new_n471), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n472), .B1(new_n518), .B2(G41), .ZN(new_n522));
  INV_X1    g0322(.A(G274), .ZN(new_n523));
  INV_X1    g0323(.A(new_n218), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n292), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT79), .A4(new_n517), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n520), .A2(new_n293), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n521), .A2(new_n526), .B1(new_n527), .B2(G257), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT80), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n513), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n521), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(G257), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n531), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(G200), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n535), .A2(new_n478), .A3(G107), .ZN(new_n536));
  XNOR2_X1  g0336(.A(G97), .B(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n538), .A2(new_n208), .B1(new_n384), .B2(new_n259), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n244), .B1(new_n353), .B2(new_n354), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n357), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  MUX2_X1   g0341(.A(new_n487), .B(new_n488), .S(G97), .Z(new_n542));
  AND2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n513), .A2(new_n528), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n534), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n528), .A2(new_n529), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n528), .A2(new_n529), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(new_n389), .A4(new_n513), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n513), .A2(new_n528), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n305), .B1(new_n541), .B2(new_n542), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n504), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G250), .B(new_n277), .C1(new_n316), .C2(new_n317), .ZN(new_n554));
  OAI211_X1 g0354(.A(G257), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n555));
  INV_X1    g0355(.A(G294), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n554), .B(new_n555), .C1(new_n334), .C2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n282), .B1(new_n527), .B2(G264), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n389), .A3(new_n531), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n531), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n305), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n208), .B(G87), .C1(new_n316), .C2(new_n317), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT22), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n461), .A2(G20), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n208), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n244), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT24), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n563), .A2(new_n571), .A3(new_n568), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n263), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n488), .A2(new_n244), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT84), .B1(new_n487), .B2(G107), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT84), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n265), .A2(new_n576), .A3(new_n244), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT25), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT25), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n575), .A2(new_n580), .A3(new_n577), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n574), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n559), .B(new_n561), .C1(new_n573), .C2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n572), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n571), .B1(new_n563), .B2(new_n568), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n357), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n560), .A2(G190), .ZN(new_n588));
  AOI21_X1  g0388(.A(G200), .B1(new_n558), .B2(new_n531), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n587), .B(new_n582), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n265), .A2(new_n247), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n488), .B2(new_n247), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n262), .A2(new_n218), .B1(G20), .B2(new_n247), .ZN(new_n594));
  AOI21_X1  g0394(.A(G20), .B1(G33), .B2(G283), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n334), .A2(G97), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT83), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT83), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT20), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(KEYINPUT20), .B(new_n594), .C1(new_n597), .C2(new_n598), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n593), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n277), .A2(G257), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G264), .A2(G1698), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n606), .C1(new_n316), .C2(new_n317), .ZN(new_n607));
  INV_X1    g0407(.A(G303), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n274), .A2(new_n608), .A3(new_n275), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n282), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n520), .A2(G270), .A3(new_n293), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n305), .B1(new_n612), .B2(new_n531), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n604), .A2(KEYINPUT21), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n531), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n616), .B(new_n603), .C1(new_n298), .C2(new_n615), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(G169), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n603), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n615), .A2(new_n389), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n604), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n614), .A2(new_n617), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n553), .A2(new_n591), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n457), .A2(new_n624), .ZN(G372));
  NAND3_X1  g0425(.A1(new_n332), .A2(KEYINPUT78), .A3(new_n350), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n360), .A2(new_n361), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n369), .B1(new_n628), .B2(KEYINPUT17), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n454), .A2(new_n392), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n445), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n367), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n303), .B(new_n304), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n307), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n561), .A2(new_n559), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n587), .B2(new_n582), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n614), .A2(new_n620), .A3(new_n622), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n590), .B(new_n504), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n546), .A2(new_n552), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n504), .A2(new_n590), .ZN(new_n643));
  INV_X1    g0443(.A(new_n641), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n620), .A2(new_n622), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n645), .A2(new_n584), .A3(new_n614), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n643), .A2(new_n644), .A3(new_n646), .A4(KEYINPUT85), .ZN(new_n647));
  INV_X1    g0447(.A(new_n503), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n549), .A2(new_n551), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n504), .A3(KEYINPUT26), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n495), .A2(new_n503), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n552), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n648), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n642), .A2(new_n647), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n457), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n635), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(KEYINPUT86), .ZN(G369));
  NAND2_X1  g0458(.A1(new_n397), .A2(new_n208), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(new_n603), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n639), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n623), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n665), .B1(new_n587), .B2(new_n582), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n591), .A2(new_n671), .B1(new_n584), .B2(new_n665), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n639), .A2(new_n665), .ZN(new_n674));
  INV_X1    g0474(.A(new_n591), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(new_n638), .B2(new_n665), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(G399));
  NOR2_X1   g0477(.A1(new_n227), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n479), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n224), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT87), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n664), .A2(KEYINPUT31), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n560), .B1(new_n530), .B2(new_n533), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT88), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT88), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n688), .B(new_n560), .C1(new_n530), .C2(new_n533), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n615), .A2(new_n491), .A3(new_n389), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n610), .A2(new_n611), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n521), .B2(new_n526), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n499), .A3(G179), .A4(new_n558), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n696), .B2(new_n550), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n499), .A2(new_n558), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n544), .A3(new_n621), .A4(KEYINPUT30), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n685), .B1(new_n692), .B2(new_n700), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n624), .A2(new_n665), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n697), .A2(new_n699), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n690), .B1(new_n686), .B2(KEYINPUT88), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n689), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n704), .B1(new_n707), .B2(new_n665), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n701), .A2(KEYINPUT89), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n702), .A2(new_n703), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n641), .A2(KEYINPUT90), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT90), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n546), .B2(new_n552), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n713), .A2(new_n640), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n654), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT29), .B(new_n665), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n655), .A2(new_n665), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n712), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n684), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(new_n226), .A2(G20), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G45), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n679), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT91), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT91), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n670), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G330), .B2(new_n668), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n218), .B1(G20), .B2(new_n305), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n227), .A2(new_n276), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n251), .B2(G45), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n224), .B2(new_n284), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n227), .A2(new_n318), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n741), .A2(G355), .B1(new_n247), .B2(new_n227), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n735), .B(new_n736), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n333), .A2(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G20), .A3(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n608), .ZN(new_n746));
  NOR4_X1   g0546(.A1(new_n208), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n276), .B(new_n746), .C1(G329), .C2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G283), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n744), .A2(G20), .A3(new_n298), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT93), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(KEYINPUT93), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n298), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n208), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n748), .B1(new_n749), .B2(new_n753), .C1(new_n556), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(G20), .A2(G179), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT92), .Z(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n298), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n333), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G311), .A2(new_n760), .B1(new_n762), .B2(G326), .ZN(new_n763));
  INV_X1    g0563(.A(G322), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n761), .A2(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n759), .A2(new_n333), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT33), .B(G317), .Z(new_n769));
  OAI221_X1 g0569(.A(new_n763), .B1(new_n764), .B2(new_n766), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G58), .A2(new_n765), .B1(new_n760), .B2(G77), .ZN(new_n771));
  INV_X1    g0571(.A(new_n762), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n771), .B1(new_n201), .B2(new_n772), .C1(new_n203), .C2(new_n768), .ZN(new_n773));
  INV_X1    g0573(.A(new_n753), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G107), .ZN(new_n775));
  INV_X1    g0575(.A(new_n747), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n776), .A2(KEYINPUT32), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n755), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(G97), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT32), .B1(new_n776), .B2(new_n777), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n745), .A2(new_n335), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n318), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n775), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n756), .A2(new_n770), .B1(new_n773), .B2(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n743), .B(new_n729), .C1(new_n785), .C2(new_n736), .ZN(new_n786));
  INV_X1    g0586(.A(new_n735), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n668), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n732), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(G396));
  OR3_X1    g0590(.A1(new_n392), .A2(KEYINPUT96), .A3(new_n665), .ZN(new_n791));
  OAI21_X1  g0591(.A(KEYINPUT96), .B1(new_n392), .B2(new_n665), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n391), .A2(new_n664), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n791), .A2(new_n792), .B1(new_n393), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n719), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n791), .A2(new_n792), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n393), .A2(new_n793), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n655), .A2(new_n665), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n712), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n712), .A2(new_n795), .A3(new_n799), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT97), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n730), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n800), .B1(new_n804), .B2(KEYINPUT98), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(KEYINPUT98), .B2(new_n804), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n736), .A2(new_n733), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n729), .B1(new_n384), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G143), .A2(new_n765), .B1(new_n760), .B2(G159), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n810), .B2(new_n772), .C1(new_n257), .C2(new_n768), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT34), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n755), .A2(new_n202), .ZN(new_n813));
  INV_X1    g0613(.A(G132), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n276), .B1(new_n745), .B2(new_n201), .C1(new_n776), .C2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(new_n774), .C2(G68), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n318), .B1(new_n745), .B2(new_n244), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT95), .Z(new_n818));
  NAND2_X1  g0618(.A1(new_n774), .A2(G87), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n478), .B2(new_n755), .C1(new_n820), .C2(new_n776), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n818), .B(new_n821), .C1(G294), .C2(new_n765), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G116), .A2(new_n760), .B1(new_n762), .B2(G303), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n749), .B2(new_n768), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT94), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n812), .A2(new_n816), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n736), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n808), .B1(new_n826), .B2(new_n827), .C1(new_n798), .C2(new_n734), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n806), .A2(new_n828), .ZN(G384));
  NAND2_X1  g0629(.A1(new_n633), .A2(new_n662), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n392), .A2(new_n664), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n799), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n405), .A2(new_n665), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n445), .A2(new_n455), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT14), .B1(new_n433), .B2(G169), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n429), .B(new_n305), .C1(new_n432), .C2(new_n426), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n441), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n443), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n435), .A2(KEYINPUT76), .A3(new_n441), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n406), .B(new_n664), .C1(new_n842), .C2(new_n454), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n833), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  INV_X1    g0646(.A(new_n311), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n358), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n662), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n629), .B2(new_n367), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n364), .A2(new_n365), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n848), .B1(new_n852), .B2(new_n849), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n626), .A2(new_n627), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n366), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n358), .A2(new_n359), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n849), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n856), .A2(new_n627), .A3(new_n626), .A4(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n846), .B1(new_n851), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n855), .A2(new_n859), .ZN(new_n862));
  OAI211_X1 g0662(.A(KEYINPUT38), .B(new_n862), .C1(new_n371), .C2(new_n850), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n830), .B1(new_n845), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n445), .A2(new_n664), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n363), .A2(new_n367), .A3(new_n370), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n662), .B1(new_n358), .B2(new_n359), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT99), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n368), .A2(new_n366), .A3(new_n871), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n857), .A2(new_n852), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n858), .A3(new_n360), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(KEYINPUT99), .A3(KEYINPUT37), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n859), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT100), .B1(new_n881), .B2(new_n846), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT100), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n883), .B(KEYINPUT38), .C1(new_n872), .C2(new_n880), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n869), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n866), .B1(new_n867), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n457), .A2(new_n721), .A3(new_n718), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n635), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n888), .B(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT101), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n707), .B2(new_n665), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n692), .A2(new_n700), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(KEYINPUT101), .A3(new_n664), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n704), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n701), .B1(new_n624), .B2(new_n665), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n794), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n844), .A2(KEYINPUT40), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n863), .B1(new_n882), .B2(new_n884), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n844), .A2(new_n864), .A3(new_n898), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n899), .A2(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n896), .A2(new_n897), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n457), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(G330), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n891), .A2(new_n908), .B1(new_n207), .B2(new_n724), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n891), .B2(new_n908), .ZN(new_n910));
  INV_X1    g0710(.A(new_n538), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n247), .B(new_n220), .C1(new_n911), .C2(KEYINPUT35), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(KEYINPUT35), .B2(new_n911), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT36), .Z(new_n914));
  OR3_X1    g0714(.A1(new_n224), .A2(new_n384), .A3(new_n323), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n201), .A2(G68), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n207), .B(G13), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  OR3_X1    g0717(.A1(new_n910), .A2(new_n914), .A3(new_n917), .ZN(G367));
  NOR2_X1   g0718(.A1(new_n713), .A2(new_n715), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n543), .A2(new_n665), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n638), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n552), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n665), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT42), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n674), .A2(new_n584), .A3(new_n590), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n920), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n649), .A2(new_n664), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n923), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n924), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT43), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n490), .A2(new_n665), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT102), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n503), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT103), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(KEYINPUT103), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n504), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n923), .B(KEYINPUT104), .C1(new_n924), .C2(new_n928), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n933), .A2(new_n934), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n931), .A2(new_n943), .A3(new_n932), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n934), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n926), .A2(new_n927), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n949), .B1(new_n673), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT105), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n951), .A2(new_n673), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n944), .A2(new_n955), .A3(new_n948), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT106), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT106), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n944), .A2(new_n958), .A3(new_n955), .A4(new_n948), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n952), .A2(new_n957), .A3(new_n953), .A4(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n950), .A2(new_n676), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT45), .Z(new_n964));
  NOR2_X1   g0764(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n950), .A2(new_n676), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n965), .B1(new_n950), .B2(new_n676), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n670), .A2(KEYINPUT108), .A3(new_n672), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n669), .A2(KEYINPUT109), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n925), .B1(new_n672), .B2(new_n674), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n722), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n964), .A2(new_n969), .A3(new_n971), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n973), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n722), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n678), .B(KEYINPUT41), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n725), .A2(G1), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n961), .A2(new_n962), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n236), .A2(new_n738), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n735), .A2(new_n736), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n228), .B2(new_n381), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n730), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n762), .A2(G143), .ZN(new_n992));
  INV_X1    g0792(.A(new_n760), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n993), .B2(new_n201), .C1(new_n777), .C2(new_n768), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n318), .B1(new_n774), .B2(G77), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n996));
  INV_X1    g0796(.A(new_n745), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n997), .A2(G58), .B1(G137), .B2(new_n747), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n203), .B2(new_n755), .C1(new_n766), .C2(new_n257), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n1000));
  OR4_X1    g0800(.A1(new_n994), .A2(new_n996), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n749), .A2(new_n993), .B1(new_n768), .B2(new_n556), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G311), .B2(new_n762), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n745), .A2(new_n247), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT46), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT110), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n774), .A2(G97), .B1(KEYINPUT110), .B2(new_n1005), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n276), .B1(new_n747), .B2(G317), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n244), .B2(new_n755), .C1(new_n1004), .C2(KEYINPUT46), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G303), .B2(new_n765), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1003), .A2(new_n1006), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1001), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n991), .B1(new_n1014), .B2(new_n736), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n941), .B2(new_n787), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n987), .A2(new_n1016), .ZN(G387));
  NOR2_X1   g0817(.A1(new_n978), .A2(new_n679), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n722), .B2(new_n976), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n255), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G50), .A2(new_n765), .B1(new_n767), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G68), .A2(new_n760), .B1(new_n762), .B2(G159), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n774), .A2(G97), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n276), .B1(new_n745), .B2(new_n384), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n755), .A2(new_n381), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G150), .C2(new_n747), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n276), .B1(new_n747), .B2(G326), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n755), .A2(new_n749), .B1(new_n745), .B2(new_n556), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G303), .A2(new_n760), .B1(new_n765), .B2(G317), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n820), .B2(new_n768), .C1(new_n764), .C2(new_n772), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT49), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1028), .B1(new_n247), .B2(new_n753), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1027), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n827), .B1(new_n1038), .B2(KEYINPUT113), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(KEYINPUT113), .B2(new_n1038), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n738), .B1(new_n241), .B2(new_n284), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n680), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n741), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1020), .A2(new_n201), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT50), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n515), .B1(new_n203), .B2(new_n384), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1045), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1043), .A2(new_n1047), .B1(G107), .B2(new_n228), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n729), .B1(new_n1048), .B2(new_n989), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1040), .B(new_n1049), .C1(new_n672), .C2(new_n787), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n976), .A2(new_n984), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1019), .A2(new_n1052), .ZN(G393));
  XNOR2_X1  g0853(.A(new_n970), .B(new_n673), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n678), .B(new_n980), .C1(new_n1054), .C2(new_n978), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n951), .A2(new_n735), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n248), .A2(new_n737), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n989), .C1(new_n478), .C2(new_n228), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n997), .A2(G283), .B1(G322), .B2(new_n747), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT115), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1060), .A2(new_n318), .A3(new_n775), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n767), .A2(G303), .B1(G116), .B2(new_n779), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1061), .B1(KEYINPUT116), .B2(new_n1062), .C1(new_n556), .C2(new_n993), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT116), .B2(new_n1062), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G311), .A2(new_n765), .B1(new_n762), .B2(G317), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT52), .Z(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n762), .B1(new_n765), .B2(G159), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  AOI22_X1  g0868(.A1(G50), .A2(new_n767), .B1(new_n760), .B2(new_n1020), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n318), .B1(new_n779), .B2(G77), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n997), .A2(G68), .B1(G143), .B2(new_n747), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT114), .ZN(new_n1072));
  AND4_X1   g0872(.A1(new_n819), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1064), .A2(new_n1066), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1058), .B(new_n730), .C1(new_n1074), .C2(new_n827), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT117), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1054), .A2(new_n984), .B1(new_n1056), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1055), .A2(new_n1077), .ZN(G390));
  AND3_X1   g0878(.A1(new_n710), .A2(G330), .A3(new_n798), .ZN(new_n1079));
  OAI21_X1  g0879(.A(KEYINPUT118), .B1(new_n1079), .B2(new_n844), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n844), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT118), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(new_n711), .C2(new_n794), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n844), .A2(new_n898), .A3(G330), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n833), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n798), .B(new_n665), .C1(new_n716), .C2(new_n717), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n832), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1079), .B2(new_n844), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n898), .A2(G330), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n1081), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n457), .A2(G330), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n890), .B1(new_n905), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n867), .B1(new_n1088), .B2(new_n844), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n900), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1079), .A2(new_n844), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n867), .B1(new_n833), .B2(new_n844), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1099), .C1(new_n887), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n351), .A2(new_n362), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n366), .A2(new_n871), .A3(KEYINPUT37), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1102), .A2(new_n873), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1105), .A2(new_n879), .B1(new_n870), .B2(new_n871), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n883), .B1(new_n1106), .B2(KEYINPUT38), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n881), .A2(KEYINPUT100), .A3(new_n846), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(new_n869), .B1(KEYINPUT39), .B2(new_n864), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n867), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n845), .A2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1110), .A2(new_n1112), .B1(new_n900), .B2(new_n1097), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1101), .B1(new_n1113), .B2(new_n1084), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1096), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n679), .B1(new_n1096), .B2(new_n1114), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1114), .A2(new_n985), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n755), .A2(new_n777), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n318), .B(new_n1119), .C1(G125), .C2(new_n747), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n745), .A2(new_n257), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT53), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1120), .B(new_n1122), .C1(new_n201), .C2(new_n753), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G128), .A2(new_n762), .B1(new_n767), .B2(G137), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1124), .B1(new_n814), .B2(new_n766), .C1(new_n993), .C2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G97), .A2(new_n760), .B1(new_n767), .B2(G107), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n247), .B2(new_n766), .C1(new_n749), .C2(new_n772), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n276), .B(new_n782), .C1(G294), .C2(new_n747), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n203), .B2(new_n753), .C1(new_n384), .C2(new_n755), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1123), .A2(new_n1126), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n736), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n729), .B1(new_n255), .B2(new_n807), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n887), .C2(new_n734), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1117), .A2(new_n1118), .A3(new_n1134), .ZN(G378));
  OAI221_X1 g0935(.A(new_n830), .B1(new_n865), .B2(new_n845), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n899), .A2(new_n900), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n901), .A2(new_n902), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n308), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n308), .A2(new_n1139), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n269), .B2(new_n662), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n271), .A3(new_n849), .A4(new_n1141), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND4_X1   g0945(.A1(G330), .A2(new_n1137), .A3(new_n1138), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n903), .B2(G330), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1136), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1137), .A2(G330), .A3(new_n1138), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1145), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n903), .A2(G330), .A3(new_n1145), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n888), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1085), .A2(new_n833), .B1(new_n1091), .B2(new_n1089), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1095), .B1(new_n1114), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1156), .A3(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n678), .B(new_n1157), .C1(new_n1158), .C2(KEYINPUT119), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT119), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1160), .B(KEYINPUT57), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1145), .A2(new_n734), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n729), .B1(new_n201), .B2(new_n807), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n755), .A2(new_n257), .B1(new_n745), .B2(new_n1125), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G128), .A2(new_n765), .B1(new_n767), .B2(G132), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n810), .B2(new_n993), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(G125), .C2(new_n762), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT59), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n774), .A2(G159), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n478), .A2(new_n768), .B1(new_n766), .B2(new_n244), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n247), .A2(new_n772), .B1(new_n993), .B2(new_n381), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n753), .A2(new_n202), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n318), .A2(new_n416), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n997), .B2(G77), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n203), .B2(new_n755), .C1(new_n749), .C2(new_n776), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1178), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1184));
  AND4_X1   g0984(.A1(new_n1174), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1164), .B1(new_n1185), .B2(new_n827), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1163), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1154), .B2(new_n984), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1162), .A2(new_n1188), .ZN(G375));
  OR2_X1    g0989(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n982), .A3(new_n1096), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n814), .A2(new_n772), .B1(new_n768), .B2(new_n1125), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G137), .B2(new_n765), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT122), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n318), .B1(new_n747), .B2(G128), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n201), .B2(new_n755), .C1(new_n777), .C2(new_n745), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1196), .B(new_n1177), .C1(G150), .C2(new_n760), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n247), .A2(new_n768), .B1(new_n772), .B2(new_n556), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G107), .B2(new_n760), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n318), .B1(new_n753), .B2(new_n384), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT121), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT121), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n776), .A2(new_n608), .B1(new_n478), .B2(new_n745), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1025), .B(new_n1204), .C1(new_n765), .C2(G283), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1200), .A2(new_n1202), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n827), .B1(new_n1198), .B2(new_n1206), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n729), .B(new_n1207), .C1(new_n203), .C2(new_n807), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT123), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT120), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n844), .A2(new_n1210), .A3(new_n734), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT120), .B1(new_n1081), .B2(new_n733), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1093), .B2(new_n984), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1191), .A2(new_n1214), .ZN(G381));
  NAND3_X1  g1015(.A1(new_n1019), .A2(new_n789), .A3(new_n1052), .ZN(new_n1216));
  OR4_X1    g1016(.A1(G384), .A2(G378), .A3(G381), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(G390), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n987), .A2(new_n1016), .A3(new_n1218), .ZN(new_n1219));
  OR3_X1    g1019(.A1(new_n1217), .A2(G375), .A3(new_n1219), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n663), .A2(G213), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT124), .Z(new_n1222));
  OR2_X1    g1022(.A1(G378), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G375), .C2(new_n1223), .ZN(G409));
  NAND2_X1  g1024(.A1(G387), .A2(G390), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G393), .A2(G396), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT125), .B1(new_n1226), .B2(new_n1216), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1225), .A2(new_n1219), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(KEYINPUT125), .A3(new_n1216), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1225), .A2(new_n1219), .B1(new_n1230), .B2(new_n1228), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1221), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1188), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1118), .A2(new_n1134), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1188), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1154), .A2(new_n982), .A3(new_n1156), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1117), .B(new_n1235), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1233), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n678), .B(new_n1096), .C1(new_n1190), .C2(new_n1240), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1190), .A2(new_n1240), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1214), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n806), .A3(new_n828), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G384), .B(new_n1214), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT62), .B1(new_n1239), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1222), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT126), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1248), .A2(KEYINPUT126), .A3(new_n1222), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1246), .A2(KEYINPUT62), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1247), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1244), .A2(new_n1245), .A3(G2897), .A4(new_n1233), .ZN(new_n1256));
  INV_X1    g1056(.A(G2897), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1222), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1246), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1252), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1232), .B1(new_n1255), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1246), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1239), .A2(new_n1246), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(KEYINPUT63), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1239), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1259), .A2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1232), .A2(KEYINPUT61), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1264), .A2(new_n1266), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1263), .A2(new_n1270), .ZN(G405));
  OR2_X1    g1071(.A1(new_n1246), .A2(KEYINPUT127), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1246), .A2(KEYINPUT127), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1234), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G378), .B1(new_n1162), .B2(new_n1188), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1272), .B(new_n1273), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1274), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(KEYINPUT127), .A3(new_n1246), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1231), .B2(new_n1229), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1276), .A2(new_n1232), .A3(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(G402));
endmodule


