

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784;

  NOR2_X1 U374 ( .A1(n743), .A2(G902), .ZN(n487) );
  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n521) );
  AND2_X1 U376 ( .A1(n562), .A2(KEYINPUT46), .ZN(n352) );
  NAND2_X2 U377 ( .A1(n643), .A2(n700), .ZN(n645) );
  XNOR2_X2 U378 ( .A(n518), .B(n517), .ZN(n719) );
  INV_X1 U379 ( .A(n577), .ZN(n587) );
  XNOR2_X1 U380 ( .A(n354), .B(G478), .ZN(n568) );
  OR2_X1 U381 ( .A1(n642), .A2(n641), .ZN(n700) );
  AND2_X1 U382 ( .A1(n377), .A2(n357), .ZN(n373) );
  XNOR2_X1 U383 ( .A(n450), .B(KEYINPUT75), .ZN(n611) );
  NOR2_X2 U384 ( .A1(n568), .A2(n543), .ZN(n688) );
  XNOR2_X1 U385 ( .A(n494), .B(KEYINPUT24), .ZN(n495) );
  XNOR2_X2 U386 ( .A(n487), .B(G469), .ZN(n556) );
  XNOR2_X1 U387 ( .A(n458), .B(n408), .ZN(n512) );
  XNOR2_X1 U388 ( .A(n457), .B(G119), .ZN(n408) );
  INV_X1 U389 ( .A(KEYINPUT3), .ZN(n457) );
  INV_X1 U390 ( .A(G116), .ZN(n459) );
  XNOR2_X1 U391 ( .A(n516), .B(KEYINPUT68), .ZN(n517) );
  XNOR2_X1 U392 ( .A(n773), .B(G146), .ZN(n507) );
  NAND2_X1 U393 ( .A1(n635), .A2(n436), .ZN(n435) );
  NAND2_X1 U394 ( .A1(KEYINPUT2), .A2(n438), .ZN(n436) );
  INV_X1 U395 ( .A(KEYINPUT65), .ZN(n438) );
  NAND2_X1 U396 ( .A1(n373), .A2(n372), .ZN(n442) );
  INV_X1 U397 ( .A(G237), .ZN(n470) );
  INV_X1 U398 ( .A(G902), .ZN(n471) );
  XNOR2_X1 U399 ( .A(G131), .B(KEYINPUT4), .ZN(n480) );
  XOR2_X1 U400 ( .A(G137), .B(G140), .Z(n490) );
  XNOR2_X1 U401 ( .A(n464), .B(G128), .ZN(n479) );
  INV_X1 U402 ( .A(G143), .ZN(n464) );
  XNOR2_X1 U403 ( .A(n462), .B(n410), .ZN(n409) );
  INV_X1 U404 ( .A(KEYINPUT88), .ZN(n410) );
  XNOR2_X1 U405 ( .A(n697), .B(n415), .ZN(n584) );
  INV_X1 U406 ( .A(KEYINPUT80), .ZN(n415) );
  NAND2_X1 U407 ( .A1(n587), .A2(n586), .ZN(n604) );
  INV_X1 U408 ( .A(KEYINPUT30), .ZN(n400) );
  XNOR2_X1 U409 ( .A(n461), .B(n539), .ZN(n407) );
  XNOR2_X1 U410 ( .A(KEYINPUT16), .B(G110), .ZN(n460) );
  INV_X1 U411 ( .A(KEYINPUT7), .ZN(n535) );
  XNOR2_X1 U412 ( .A(n479), .B(G134), .ZN(n418) );
  XNOR2_X1 U413 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U414 ( .A(G101), .B(G104), .Z(n486) );
  NAND2_X1 U415 ( .A1(n355), .A2(n386), .ZN(n385) );
  XNOR2_X1 U416 ( .A(n719), .B(n542), .ZN(n384) );
  INV_X1 U417 ( .A(n602), .ZN(n440) );
  INV_X1 U418 ( .A(n782), .ZN(n390) );
  XOR2_X1 U419 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n509) );
  XNOR2_X1 U420 ( .A(G116), .B(G137), .ZN(n511) );
  AND2_X1 U421 ( .A1(n433), .A2(n434), .ZN(n432) );
  NAND2_X1 U422 ( .A1(n437), .A2(n435), .ZN(n434) );
  NAND2_X1 U423 ( .A1(n634), .A2(n438), .ZN(n437) );
  NAND2_X1 U424 ( .A1(n705), .A2(n706), .ZN(n702) );
  INV_X1 U425 ( .A(n426), .ZN(n421) );
  INV_X1 U426 ( .A(n604), .ZN(n405) );
  INV_X2 U427 ( .A(G953), .ZN(n765) );
  XOR2_X1 U428 ( .A(KEYINPUT95), .B(KEYINPUT98), .Z(n526) );
  XNOR2_X1 U429 ( .A(G143), .B(G140), .ZN(n525) );
  XNOR2_X1 U430 ( .A(G113), .B(G131), .ZN(n414) );
  XNOR2_X1 U431 ( .A(KEYINPUT96), .B(KEYINPUT12), .ZN(n527) );
  XOR2_X1 U432 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n528) );
  XNOR2_X1 U433 ( .A(n409), .B(n463), .ZN(n468) );
  XNOR2_X1 U434 ( .A(n446), .B(n445), .ZN(n639) );
  INV_X1 U435 ( .A(KEYINPUT48), .ZN(n445) );
  NOR2_X1 U436 ( .A1(n448), .A2(n576), .ZN(n447) );
  NAND2_X1 U437 ( .A1(n427), .A2(n359), .ZN(n736) );
  XNOR2_X1 U438 ( .A(n394), .B(n392), .ZN(n735) );
  XNOR2_X1 U439 ( .A(n393), .B(KEYINPUT41), .ZN(n392) );
  NOR2_X1 U440 ( .A1(n702), .A2(n595), .ZN(n394) );
  INV_X1 U441 ( .A(KEYINPUT108), .ZN(n393) );
  INV_X1 U442 ( .A(n552), .ZN(n417) );
  XNOR2_X1 U443 ( .A(n519), .B(n400), .ZN(n399) );
  XNOR2_X1 U444 ( .A(n553), .B(KEYINPUT106), .ZN(n554) );
  OR2_X1 U445 ( .A1(n716), .A2(KEYINPUT103), .ZN(n376) );
  BUF_X1 U446 ( .A(n719), .Z(n401) );
  NAND2_X1 U447 ( .A1(G953), .A2(G900), .ZN(n775) );
  XNOR2_X1 U448 ( .A(n541), .B(n397), .ZN(n749) );
  XNOR2_X1 U449 ( .A(n538), .B(n537), .ZN(n541) );
  XNOR2_X1 U450 ( .A(n482), .B(n429), .ZN(n428) );
  XNOR2_X1 U451 ( .A(n485), .B(n486), .ZN(n429) );
  XNOR2_X1 U452 ( .A(n454), .B(n452), .ZN(n782) );
  XNOR2_X1 U453 ( .A(n558), .B(n453), .ZN(n452) );
  NAND2_X1 U454 ( .A1(n735), .A2(n563), .ZN(n454) );
  INV_X1 U455 ( .A(KEYINPUT109), .ZN(n453) );
  XNOR2_X1 U456 ( .A(n561), .B(n560), .ZN(n784) );
  XNOR2_X1 U457 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n560) );
  AND2_X1 U458 ( .A1(n416), .A2(n587), .ZN(n697) );
  XNOR2_X1 U459 ( .A(n580), .B(KEYINPUT36), .ZN(n416) );
  NOR2_X1 U460 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U461 ( .A(n592), .ZN(n403) );
  NOR2_X1 U462 ( .A1(n353), .A2(n382), .ZN(n381) );
  INV_X1 U463 ( .A(n384), .ZN(n382) );
  INV_X1 U464 ( .A(n688), .ZN(n692) );
  OR2_X1 U465 ( .A1(n716), .A2(n614), .ZN(n353) );
  OR2_X1 U466 ( .A1(G902), .A2(n749), .ZN(n354) );
  AND2_X1 U467 ( .A1(n423), .A2(n420), .ZN(n355) );
  OR2_X1 U468 ( .A1(n556), .A2(n715), .ZN(n356) );
  AND2_X1 U469 ( .A1(n376), .A2(n599), .ZN(n357) );
  AND2_X1 U470 ( .A1(n589), .A2(n588), .ZN(n358) );
  INV_X1 U471 ( .A(n450), .ZN(n703) );
  AND2_X1 U472 ( .A1(n419), .A2(n426), .ZN(n359) );
  AND2_X1 U473 ( .A1(n534), .A2(G221), .ZN(n360) );
  AND2_X1 U474 ( .A1(G214), .A2(n521), .ZN(n361) );
  BUF_X1 U475 ( .A(n577), .Z(n716) );
  NAND2_X1 U476 ( .A1(n716), .A2(n614), .ZN(n362) );
  AND2_X1 U477 ( .A1(n422), .A2(n405), .ZN(n363) );
  XOR2_X1 U478 ( .A(KEYINPUT85), .B(KEYINPUT33), .Z(n364) );
  XOR2_X1 U479 ( .A(n598), .B(KEYINPUT22), .Z(n365) );
  XOR2_X1 U480 ( .A(n591), .B(n590), .Z(n366) );
  XNOR2_X1 U481 ( .A(G902), .B(KEYINPUT15), .ZN(n634) );
  XNOR2_X1 U482 ( .A(n507), .B(n428), .ZN(n743) );
  INV_X1 U483 ( .A(KEYINPUT46), .ZN(n449) );
  XNOR2_X1 U484 ( .A(n407), .B(n512), .ZN(n764) );
  AND2_X1 U485 ( .A1(n635), .A2(n438), .ZN(n367) );
  AND2_X1 U486 ( .A1(n633), .A2(KEYINPUT65), .ZN(n368) );
  NOR2_X2 U487 ( .A1(G902), .A2(n647), .ZN(n533) );
  OR2_X1 U488 ( .A1(n569), .A2(n568), .ZN(n595) );
  XNOR2_X1 U489 ( .A(n694), .B(KEYINPUT101), .ZN(n565) );
  OR2_X2 U490 ( .A1(n565), .A2(n688), .ZN(n450) );
  AND2_X1 U491 ( .A1(n373), .A2(n372), .ZN(n369) );
  NAND2_X1 U492 ( .A1(n375), .A2(n374), .ZN(n372) );
  XNOR2_X1 U493 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U494 ( .A1(n543), .A2(n568), .ZN(n694) );
  XNOR2_X1 U495 ( .A(n540), .B(n418), .ZN(n397) );
  XNOR2_X1 U496 ( .A(n418), .B(n480), .ZN(n773) );
  XNOR2_X1 U497 ( .A(n495), .B(n360), .ZN(n411) );
  BUF_X1 U498 ( .A(n413), .Z(n370) );
  XNOR2_X1 U499 ( .A(n481), .B(G107), .ZN(n482) );
  XNOR2_X1 U500 ( .A(n556), .B(KEYINPUT1), .ZN(n577) );
  NOR2_X1 U501 ( .A1(n715), .A2(n556), .ZN(n608) );
  XNOR2_X1 U502 ( .A(n411), .B(n771), .ZN(n753) );
  AND2_X1 U503 ( .A1(n639), .A2(n456), .ZN(n640) );
  XNOR2_X1 U504 ( .A(n502), .B(n501), .ZN(n712) );
  BUF_X1 U505 ( .A(n742), .Z(n751) );
  NAND2_X1 U506 ( .A1(n600), .A2(n384), .ZN(n383) );
  AND2_X2 U507 ( .A1(n442), .A2(n371), .ZN(n624) );
  XNOR2_X1 U508 ( .A(n371), .B(G119), .ZN(G21) );
  XNOR2_X2 U509 ( .A(n601), .B(KEYINPUT32), .ZN(n371) );
  INV_X1 U510 ( .A(KEYINPUT103), .ZN(n374) );
  INV_X1 U511 ( .A(n600), .ZN(n375) );
  NAND2_X1 U512 ( .A1(n600), .A2(n378), .ZN(n377) );
  AND2_X1 U513 ( .A1(n716), .A2(KEYINPUT103), .ZN(n378) );
  XNOR2_X2 U514 ( .A(n379), .B(KEYINPUT19), .ZN(n413) );
  NAND2_X2 U515 ( .A1(n564), .A2(n706), .ZN(n379) );
  XNOR2_X2 U516 ( .A(n380), .B(n473), .ZN(n564) );
  NAND2_X1 U517 ( .A1(n667), .A2(n634), .ZN(n380) );
  NAND2_X1 U518 ( .A1(n381), .A2(n600), .ZN(n601) );
  NOR2_X1 U519 ( .A1(n383), .A2(n362), .ZN(n674) );
  OR2_X1 U520 ( .A1(n384), .A2(n364), .ZN(n425) );
  NAND2_X1 U521 ( .A1(n384), .A2(n364), .ZN(n426) );
  NOR2_X1 U522 ( .A1(n546), .A2(n384), .ZN(n547) );
  XNOR2_X1 U523 ( .A(n507), .B(n515), .ZN(n656) );
  XNOR2_X1 U524 ( .A(n385), .B(n366), .ZN(n404) );
  NAND2_X1 U525 ( .A1(n363), .A2(n609), .ZN(n386) );
  NAND2_X1 U526 ( .A1(n387), .A2(n449), .ZN(n389) );
  NAND2_X1 U527 ( .A1(n390), .A2(n562), .ZN(n387) );
  NAND2_X1 U528 ( .A1(n389), .A2(n388), .ZN(n391) );
  NAND2_X1 U529 ( .A1(n352), .A2(n390), .ZN(n388) );
  NAND2_X1 U530 ( .A1(n447), .A2(n391), .ZN(n446) );
  XNOR2_X1 U531 ( .A(n395), .B(n489), .ZN(n451) );
  XNOR2_X1 U532 ( .A(n524), .B(n361), .ZN(n395) );
  NAND2_X1 U533 ( .A1(n639), .A2(n585), .ZN(n776) );
  NAND2_X1 U534 ( .A1(n396), .A2(n689), .ZN(n583) );
  NAND2_X1 U535 ( .A1(n582), .A2(KEYINPUT74), .ZN(n396) );
  NOR2_X2 U536 ( .A1(n611), .A2(KEYINPUT47), .ZN(n581) );
  XNOR2_X2 U537 ( .A(n533), .B(n532), .ZN(n569) );
  NAND2_X1 U538 ( .A1(n624), .A2(KEYINPUT44), .ZN(n441) );
  XNOR2_X1 U539 ( .A(n469), .B(n764), .ZN(n667) );
  INV_X2 U540 ( .A(G125), .ZN(n444) );
  NAND2_X1 U541 ( .A1(n630), .A2(n398), .ZN(n631) );
  NAND2_X1 U542 ( .A1(n629), .A2(n783), .ZN(n398) );
  NAND2_X1 U543 ( .A1(n608), .A2(n399), .ZN(n520) );
  XNOR2_X2 U544 ( .A(n402), .B(KEYINPUT39), .ZN(n559) );
  NAND2_X1 U545 ( .A1(n571), .A2(n705), .ZN(n402) );
  NOR2_X2 U546 ( .A1(n605), .A2(n597), .ZN(n406) );
  NAND2_X1 U547 ( .A1(n404), .A2(n403), .ZN(n593) );
  XNOR2_X2 U548 ( .A(n406), .B(n365), .ZN(n600) );
  NAND2_X1 U549 ( .A1(n441), .A2(n440), .ZN(n618) );
  INV_X1 U550 ( .A(n425), .ZN(n422) );
  XNOR2_X1 U551 ( .A(n412), .B(n492), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n491), .B(KEYINPUT91), .ZN(n412) );
  INV_X1 U553 ( .A(n682), .ZN(n689) );
  NAND2_X1 U554 ( .A1(n682), .A2(KEYINPUT74), .ZN(n566) );
  NAND2_X1 U555 ( .A1(n563), .A2(n370), .ZN(n682) );
  XNOR2_X1 U556 ( .A(n555), .B(n554), .ZN(n557) );
  XNOR2_X1 U557 ( .A(n523), .B(n414), .ZN(n524) );
  XNOR2_X2 U558 ( .A(G122), .B(G104), .ZN(n523) );
  NAND2_X1 U559 ( .A1(n417), .A2(n688), .ZN(n546) );
  XNOR2_X2 U560 ( .A(n569), .B(KEYINPUT99), .ZN(n543) );
  OR2_X1 U561 ( .A1(n604), .A2(n425), .ZN(n419) );
  NAND2_X1 U562 ( .A1(n609), .A2(n421), .ZN(n420) );
  NAND2_X1 U563 ( .A1(n424), .A2(n609), .ZN(n423) );
  INV_X1 U564 ( .A(n427), .ZN(n424) );
  NAND2_X1 U565 ( .A1(n604), .A2(n364), .ZN(n427) );
  NAND2_X1 U566 ( .A1(n583), .A2(n584), .ZN(n448) );
  NOR2_X2 U567 ( .A1(n712), .A2(n713), .ZN(n586) );
  NAND2_X1 U568 ( .A1(n432), .A2(n430), .ZN(n643) );
  NAND2_X1 U569 ( .A1(n431), .A2(n367), .ZN(n430) );
  INV_X1 U570 ( .A(n439), .ZN(n431) );
  NAND2_X1 U571 ( .A1(n439), .A2(n368), .ZN(n433) );
  NAND2_X1 U572 ( .A1(n439), .A2(n633), .ZN(n701) );
  NAND2_X1 U573 ( .A1(n632), .A2(n758), .ZN(n439) );
  XNOR2_X2 U574 ( .A(n443), .B(KEYINPUT0), .ZN(n605) );
  NAND2_X1 U575 ( .A1(n413), .A2(n358), .ZN(n443) );
  XNOR2_X2 U576 ( .A(n444), .B(G146), .ZN(n488) );
  INV_X1 U577 ( .A(n489), .ZN(n522) );
  XNOR2_X1 U578 ( .A(n531), .B(n451), .ZN(n647) );
  XNOR2_X1 U579 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U580 ( .A(n488), .B(KEYINPUT10), .ZN(n489) );
  XOR2_X1 U581 ( .A(KEYINPUT78), .B(KEYINPUT35), .Z(n455) );
  NOR2_X1 U582 ( .A1(n638), .A2(n637), .ZN(n456) );
  INV_X1 U583 ( .A(n784), .ZN(n562) );
  INV_X1 U584 ( .A(KEYINPUT90), .ZN(n483) );
  INV_X1 U585 ( .A(KEYINPUT28), .ZN(n553) );
  XNOR2_X1 U586 ( .A(n536), .B(n535), .ZN(n537) );
  INV_X1 U587 ( .A(KEYINPUT67), .ZN(n590) );
  INV_X1 U588 ( .A(G472), .ZN(n516) );
  INV_X1 U589 ( .A(n757), .ZN(n660) );
  XNOR2_X1 U590 ( .A(n743), .B(n744), .ZN(n745) );
  XNOR2_X1 U591 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U592 ( .A(G113), .B(G101), .ZN(n458) );
  XNOR2_X1 U593 ( .A(n459), .B(G107), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n523), .B(n460), .ZN(n461) );
  XOR2_X1 U595 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n463) );
  XNOR2_X1 U596 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n462) );
  NAND2_X1 U597 ( .A1(G224), .A2(n765), .ZN(n465) );
  XNOR2_X1 U598 ( .A(n488), .B(n465), .ZN(n466) );
  XNOR2_X1 U599 ( .A(n466), .B(n479), .ZN(n467) );
  XNOR2_X1 U600 ( .A(n467), .B(n468), .ZN(n469) );
  NAND2_X1 U601 ( .A1(n471), .A2(n470), .ZN(n506) );
  NAND2_X1 U602 ( .A1(n506), .A2(G210), .ZN(n472) );
  XNOR2_X1 U603 ( .A(n472), .B(KEYINPUT89), .ZN(n473) );
  XOR2_X1 U604 ( .A(KEYINPUT70), .B(KEYINPUT38), .Z(n474) );
  XNOR2_X1 U605 ( .A(n564), .B(n474), .ZN(n705) );
  NAND2_X1 U606 ( .A1(G234), .A2(G237), .ZN(n475) );
  XNOR2_X1 U607 ( .A(n475), .B(KEYINPUT14), .ZN(n731) );
  NOR2_X1 U608 ( .A1(G953), .A2(G952), .ZN(n477) );
  NOR2_X1 U609 ( .A1(G902), .A2(n765), .ZN(n476) );
  NOR2_X1 U610 ( .A1(n477), .A2(n476), .ZN(n478) );
  AND2_X1 U611 ( .A1(n731), .A2(n478), .ZN(n589) );
  NAND2_X1 U612 ( .A1(n589), .A2(n775), .ZN(n544) );
  XOR2_X1 U613 ( .A(n490), .B(G110), .Z(n481) );
  NAND2_X1 U614 ( .A1(G227), .A2(n765), .ZN(n484) );
  XOR2_X1 U615 ( .A(n490), .B(n522), .Z(n771) );
  XOR2_X1 U616 ( .A(KEYINPUT23), .B(G110), .Z(n492) );
  XNOR2_X1 U617 ( .A(G119), .B(G128), .ZN(n491) );
  INV_X1 U618 ( .A(n493), .ZN(n494) );
  NAND2_X1 U619 ( .A1(n765), .A2(G234), .ZN(n496) );
  XOR2_X1 U620 ( .A(KEYINPUT8), .B(n496), .Z(n534) );
  NOR2_X1 U621 ( .A1(n753), .A2(G902), .ZN(n502) );
  XOR2_X1 U622 ( .A(KEYINPUT25), .B(KEYINPUT72), .Z(n499) );
  NAND2_X1 U623 ( .A1(G234), .A2(n634), .ZN(n497) );
  XNOR2_X1 U624 ( .A(KEYINPUT20), .B(n497), .ZN(n503) );
  NAND2_X1 U625 ( .A1(G217), .A2(n503), .ZN(n498) );
  XNOR2_X1 U626 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U627 ( .A(n500), .B(KEYINPUT92), .ZN(n501) );
  AND2_X1 U628 ( .A1(n503), .A2(G221), .ZN(n505) );
  INV_X1 U629 ( .A(KEYINPUT21), .ZN(n504) );
  XNOR2_X1 U630 ( .A(n505), .B(n504), .ZN(n713) );
  INV_X1 U631 ( .A(n586), .ZN(n715) );
  NAND2_X1 U632 ( .A1(n506), .A2(G214), .ZN(n706) );
  NAND2_X1 U633 ( .A1(n521), .A2(G210), .ZN(n508) );
  XNOR2_X1 U634 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U635 ( .A(n510), .B(KEYINPUT71), .Z(n514) );
  XNOR2_X1 U636 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U637 ( .A(n514), .B(n513), .ZN(n515) );
  NOR2_X1 U638 ( .A1(n656), .A2(G902), .ZN(n518) );
  NAND2_X1 U639 ( .A1(n706), .A2(n719), .ZN(n519) );
  NOR2_X2 U640 ( .A1(n544), .A2(n520), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n526), .B(n525), .ZN(n530) );
  XNOR2_X1 U642 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U643 ( .A(n530), .B(n529), .Z(n531) );
  XNOR2_X1 U644 ( .A(KEYINPUT13), .B(G475), .ZN(n532) );
  NAND2_X1 U645 ( .A1(G217), .A2(n534), .ZN(n538) );
  XOR2_X1 U646 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n536) );
  XNOR2_X1 U647 ( .A(n539), .B(G122), .ZN(n540) );
  NAND2_X1 U648 ( .A1(n559), .A2(n565), .ZN(n699) );
  XNOR2_X1 U649 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n542) );
  NOR2_X1 U650 ( .A1(n713), .A2(n544), .ZN(n545) );
  NAND2_X1 U651 ( .A1(n712), .A2(n545), .ZN(n552) );
  NAND2_X1 U652 ( .A1(n547), .A2(n706), .ZN(n579) );
  XNOR2_X1 U653 ( .A(n579), .B(KEYINPUT104), .ZN(n548) );
  NOR2_X1 U654 ( .A1(n548), .A2(n587), .ZN(n549) );
  XNOR2_X1 U655 ( .A(KEYINPUT43), .B(n549), .ZN(n550) );
  XNOR2_X1 U656 ( .A(n550), .B(KEYINPUT105), .ZN(n551) );
  INV_X1 U657 ( .A(n564), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n551), .A2(n578), .ZN(n673) );
  AND2_X1 U659 ( .A1(n699), .A2(n673), .ZN(n585) );
  XOR2_X1 U660 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n558) );
  INV_X1 U661 ( .A(n401), .ZN(n603) );
  NOR2_X1 U662 ( .A1(n603), .A2(n552), .ZN(n555) );
  NOR2_X1 U663 ( .A1(n557), .A2(n556), .ZN(n563) );
  NAND2_X1 U664 ( .A1(n559), .A2(n688), .ZN(n561) );
  NAND2_X1 U665 ( .A1(n566), .A2(n450), .ZN(n567) );
  NAND2_X1 U666 ( .A1(n567), .A2(KEYINPUT47), .ZN(n575) );
  NAND2_X1 U667 ( .A1(n569), .A2(n568), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n592), .A2(n578), .ZN(n570) );
  AND2_X1 U669 ( .A1(n571), .A2(n570), .ZN(n686) );
  XNOR2_X1 U670 ( .A(n686), .B(KEYINPUT76), .ZN(n573) );
  NOR2_X1 U671 ( .A1(KEYINPUT74), .A2(KEYINPUT47), .ZN(n572) );
  NOR2_X1 U672 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U673 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U674 ( .A(KEYINPUT69), .B(n581), .ZN(n582) );
  INV_X1 U675 ( .A(n776), .ZN(n632) );
  NAND2_X1 U676 ( .A1(G953), .A2(G898), .ZN(n588) );
  INV_X1 U677 ( .A(n605), .ZN(n609) );
  INV_X1 U678 ( .A(KEYINPUT34), .ZN(n591) );
  XNOR2_X2 U679 ( .A(n593), .B(n455), .ZN(n783) );
  INV_X1 U680 ( .A(KEYINPUT81), .ZN(n627) );
  INV_X1 U681 ( .A(KEYINPUT44), .ZN(n621) );
  AND2_X1 U682 ( .A1(n627), .A2(n621), .ZN(n602) );
  OR2_X1 U683 ( .A1(KEYINPUT81), .A2(n602), .ZN(n594) );
  NOR2_X1 U684 ( .A1(n783), .A2(n594), .ZN(n620) );
  INV_X1 U685 ( .A(n595), .ZN(n708) );
  INV_X1 U686 ( .A(n713), .ZN(n596) );
  NAND2_X1 U687 ( .A1(n708), .A2(n596), .ZN(n597) );
  INV_X1 U688 ( .A(KEYINPUT66), .ZN(n598) );
  INV_X1 U689 ( .A(n712), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n401), .A2(n614), .ZN(n599) );
  OR2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n724) );
  NOR2_X1 U692 ( .A1(n724), .A2(n605), .ZN(n607) );
  XNOR2_X1 U693 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n606) );
  XNOR2_X1 U694 ( .A(n607), .B(n606), .ZN(n695) );
  NOR2_X1 U695 ( .A1(n356), .A2(n401), .ZN(n610) );
  NAND2_X1 U696 ( .A1(n610), .A2(n609), .ZN(n679) );
  NAND2_X1 U697 ( .A1(n695), .A2(n679), .ZN(n613) );
  INV_X1 U698 ( .A(n611), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n613), .A2(n612), .ZN(n616) );
  INV_X1 U700 ( .A(n674), .ZN(n615) );
  AND2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n624), .A2(n621), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n622), .A2(KEYINPUT82), .ZN(n626) );
  INV_X1 U706 ( .A(KEYINPUT82), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X2 U710 ( .A(n631), .B(KEYINPUT45), .ZN(n758) );
  INV_X1 U711 ( .A(KEYINPUT2), .ZN(n633) );
  INV_X1 U712 ( .A(n634), .ZN(n635) );
  INV_X1 U713 ( .A(n758), .ZN(n642) );
  INV_X1 U714 ( .A(n673), .ZN(n638) );
  NAND2_X1 U715 ( .A1(KEYINPUT2), .A2(n699), .ZN(n636) );
  XOR2_X1 U716 ( .A(KEYINPUT73), .B(n636), .Z(n637) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT77), .ZN(n641) );
  INV_X1 U718 ( .A(KEYINPUT64), .ZN(n644) );
  XNOR2_X2 U719 ( .A(n645), .B(n644), .ZN(n742) );
  NAND2_X1 U720 ( .A1(n742), .A2(G475), .ZN(n649) );
  XOR2_X1 U721 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n646) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(n651) );
  INV_X1 U723 ( .A(G952), .ZN(n650) );
  AND2_X1 U724 ( .A1(n650), .A2(G953), .ZN(n757) );
  NOR2_X2 U725 ( .A1(n651), .A2(n757), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n652), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U727 ( .A1(n742), .A2(G472), .ZN(n658) );
  XOR2_X1 U728 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n654) );
  XNOR2_X1 U729 ( .A(KEYINPUT62), .B(KEYINPUT86), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  INV_X1 U733 ( .A(n659), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n662), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U736 ( .A1(n742), .A2(G210), .ZN(n669) );
  XNOR2_X1 U737 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n663), .B(KEYINPUT55), .ZN(n664) );
  XOR2_X1 U739 ( .A(n664), .B(KEYINPUT54), .Z(n665) );
  XOR2_X1 U740 ( .A(n665), .B(KEYINPUT121), .Z(n666) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X2 U743 ( .A1(n670), .A2(n757), .ZN(n672) );
  XOR2_X1 U744 ( .A(KEYINPUT56), .B(KEYINPUT79), .Z(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(n671), .ZN(G51) );
  XNOR2_X1 U746 ( .A(n673), .B(G140), .ZN(G42) );
  XNOR2_X1 U747 ( .A(G101), .B(n674), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n675), .B(KEYINPUT113), .ZN(G3) );
  NOR2_X1 U749 ( .A1(n692), .A2(n679), .ZN(n676) );
  XOR2_X1 U750 ( .A(G104), .B(n676), .Z(G6) );
  XOR2_X1 U751 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n678) );
  XNOR2_X1 U752 ( .A(G107), .B(KEYINPUT27), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n678), .B(n677), .ZN(n681) );
  NOR2_X1 U754 ( .A1(n694), .A2(n679), .ZN(n680) );
  XOR2_X1 U755 ( .A(n681), .B(n680), .Z(G9) );
  XOR2_X1 U756 ( .A(n369), .B(G110), .Z(G12) );
  NOR2_X1 U757 ( .A1(n682), .A2(n694), .ZN(n684) );
  XNOR2_X1 U758 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n683) );
  XNOR2_X1 U759 ( .A(n684), .B(n683), .ZN(n685) );
  XOR2_X1 U760 ( .A(G128), .B(n685), .Z(G30) );
  XOR2_X1 U761 ( .A(G143), .B(n686), .Z(n687) );
  XNOR2_X1 U762 ( .A(KEYINPUT116), .B(n687), .ZN(G45) );
  XOR2_X1 U763 ( .A(G146), .B(KEYINPUT117), .Z(n691) );
  NAND2_X1 U764 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U765 ( .A(n691), .B(n690), .ZN(G48) );
  NOR2_X1 U766 ( .A1(n695), .A2(n692), .ZN(n693) );
  XOR2_X1 U767 ( .A(G113), .B(n693), .Z(G15) );
  NOR2_X1 U768 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U769 ( .A(G116), .B(n696), .Z(G18) );
  XNOR2_X1 U770 ( .A(G125), .B(n697), .ZN(n698) );
  XNOR2_X1 U771 ( .A(n698), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U772 ( .A(G134), .B(n699), .ZN(G36) );
  AND2_X1 U773 ( .A1(n701), .A2(n700), .ZN(n740) );
  NOR2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U775 ( .A(n704), .B(KEYINPUT119), .ZN(n710) );
  OR2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U777 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U778 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n711), .A2(n736), .ZN(n728) );
  AND2_X1 U780 ( .A1(n712), .A2(n713), .ZN(n714) );
  XNOR2_X1 U781 ( .A(KEYINPUT49), .B(n714), .ZN(n722) );
  XOR2_X1 U782 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n718) );
  NAND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U784 ( .A(n718), .B(n717), .ZN(n720) );
  NOR2_X1 U785 ( .A1(n720), .A2(n401), .ZN(n721) );
  NAND2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U788 ( .A(KEYINPUT51), .B(n725), .Z(n726) );
  NAND2_X1 U789 ( .A1(n726), .A2(n735), .ZN(n727) );
  NAND2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U791 ( .A(n729), .B(KEYINPUT120), .ZN(n730) );
  XOR2_X1 U792 ( .A(KEYINPUT52), .B(n730), .Z(n733) );
  NAND2_X1 U793 ( .A1(G952), .A2(n731), .ZN(n732) );
  NOR2_X1 U794 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U795 ( .A1(G953), .A2(n734), .ZN(n738) );
  NAND2_X1 U796 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U797 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U798 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U799 ( .A(KEYINPUT53), .B(n741), .ZN(G75) );
  NAND2_X1 U800 ( .A1(n751), .A2(G469), .ZN(n746) );
  XOR2_X1 U801 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n744) );
  NOR2_X1 U802 ( .A1(n757), .A2(n747), .ZN(G54) );
  NAND2_X1 U803 ( .A1(n751), .A2(G478), .ZN(n748) );
  XNOR2_X1 U804 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U805 ( .A1(n757), .A2(n750), .ZN(G63) );
  NAND2_X1 U806 ( .A1(n751), .A2(G217), .ZN(n755) );
  INV_X1 U807 ( .A(KEYINPUT123), .ZN(n752) );
  XNOR2_X1 U808 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U809 ( .A1(n757), .A2(n756), .ZN(G66) );
  NAND2_X1 U810 ( .A1(n758), .A2(n765), .ZN(n763) );
  NAND2_X1 U811 ( .A1(G224), .A2(G953), .ZN(n759) );
  XNOR2_X1 U812 ( .A(n759), .B(KEYINPUT61), .ZN(n760) );
  XNOR2_X1 U813 ( .A(KEYINPUT124), .B(n760), .ZN(n761) );
  NAND2_X1 U814 ( .A1(n761), .A2(G898), .ZN(n762) );
  NAND2_X1 U815 ( .A1(n763), .A2(n762), .ZN(n770) );
  INV_X1 U816 ( .A(n764), .ZN(n767) );
  OR2_X1 U817 ( .A1(G898), .A2(n765), .ZN(n766) );
  NAND2_X1 U818 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n768), .B(KEYINPUT125), .ZN(n769) );
  XNOR2_X1 U820 ( .A(n770), .B(n769), .ZN(G69) );
  XOR2_X1 U821 ( .A(n771), .B(KEYINPUT90), .Z(n772) );
  XNOR2_X1 U822 ( .A(n773), .B(n772), .ZN(n777) );
  XNOR2_X1 U823 ( .A(n777), .B(G227), .ZN(n774) );
  NOR2_X1 U824 ( .A1(n775), .A2(n774), .ZN(n780) );
  XOR2_X1 U825 ( .A(n777), .B(n776), .Z(n778) );
  NOR2_X1 U826 ( .A1(G953), .A2(n778), .ZN(n779) );
  NOR2_X1 U827 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U828 ( .A(n781), .B(KEYINPUT126), .ZN(G72) );
  XOR2_X1 U829 ( .A(G137), .B(n782), .Z(G39) );
  XNOR2_X1 U830 ( .A(n783), .B(G122), .ZN(G24) );
  XOR2_X1 U831 ( .A(n784), .B(G131), .Z(G33) );
endmodule

