//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n187));
  INV_X1    g001(.A(G478), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT15), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT9), .B(G234), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(G217), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G116), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(G122), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n202), .A2(G122), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G107), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n210), .A3(new_n207), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n201), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT13), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n195), .B2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT13), .A3(G128), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n198), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G134), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(KEYINPUT82), .A3(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n208), .A2(KEYINPUT14), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g039(.A(G107), .B1(new_n206), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n198), .ZN(new_n228));
  OAI21_X1  g042(.A(G134), .B1(new_n228), .B2(new_n196), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n200), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n230), .A2(new_n211), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n223), .A2(KEYINPUT83), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT83), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n212), .A2(new_n222), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n194), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n221), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT82), .B1(new_n217), .B2(G134), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n211), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n210), .B1(new_n206), .B2(new_n207), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n200), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT83), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n227), .A2(new_n231), .ZN(new_n243));
  AND4_X1   g057(.A1(new_n234), .A2(new_n242), .A3(new_n243), .A4(new_n194), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n235), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n189), .B1(new_n245), .B2(G902), .ZN(new_n246));
  NAND2_X1  g060(.A1(G234), .A2(G237), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(G952), .A3(new_n192), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT21), .B(G898), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT84), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(G902), .A3(G953), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n234), .A3(new_n243), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n193), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n232), .A2(new_n234), .A3(new_n194), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G902), .ZN(new_n257));
  INV_X1    g071(.A(new_n189), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n246), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G140), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G125), .ZN(new_n262));
  INV_X1    g076(.A(G125), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G140), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  XNOR2_X1  g080(.A(G125), .B(G140), .ZN(new_n267));
  INV_X1    g081(.A(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT18), .A2(G131), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G237), .A2(G953), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n273), .A2(G143), .A3(G214), .ZN(new_n274));
  AOI21_X1  g088(.A(G143), .B1(new_n273), .B2(G214), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(G214), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n215), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(G143), .A3(G214), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(new_n271), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT79), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n270), .A2(new_n276), .A3(new_n280), .A4(KEYINPUT79), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G113), .B(G122), .ZN(new_n286));
  INV_X1    g100(.A(G104), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n286), .B(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G131), .B1(new_n274), .B2(new_n275), .ZN(new_n289));
  INV_X1    g103(.A(G131), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n278), .A2(new_n290), .A3(new_n279), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT17), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT17), .B(G131), .C1(new_n274), .C2(new_n275), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT16), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n261), .A3(G125), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n265), .B2(new_n295), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n268), .ZN(new_n298));
  OAI211_X1 g112(.A(G146), .B(new_n296), .C1(new_n265), .C2(new_n295), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n293), .A2(new_n294), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n285), .A2(new_n288), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(new_n289), .B2(new_n291), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT19), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n262), .B(new_n264), .C1(KEYINPUT81), .C2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n305), .B(new_n268), .C1(new_n267), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n299), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n289), .A2(new_n291), .A3(new_n302), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n309), .A2(new_n310), .B1(new_n283), .B2(new_n284), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n301), .B1(new_n311), .B2(new_n288), .ZN(new_n312));
  NOR2_X1   g126(.A1(G475), .A2(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT20), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(new_n316), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n301), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n288), .B1(new_n285), .B2(new_n300), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n257), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G475), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n187), .B1(new_n260), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n258), .B1(new_n256), .B2(new_n257), .ZN(new_n325));
  AOI211_X1 g139(.A(G902), .B(new_n189), .C1(new_n254), .C2(new_n255), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n315), .A2(new_n317), .B1(G475), .B2(new_n321), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT85), .A4(new_n252), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n203), .A2(new_n205), .A3(G119), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n202), .A2(G119), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(KEYINPUT5), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G113), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n287), .A2(G107), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n210), .A2(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(G101), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(new_n287), .B2(G107), .ZN(new_n344));
  AOI21_X1  g158(.A(G101), .B1(new_n287), .B2(G107), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n210), .A3(G104), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n337), .A2(KEYINPUT2), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G113), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n333), .A2(new_n335), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n340), .A2(new_n349), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n287), .A2(G107), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n344), .A2(new_n347), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G101), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n333), .A2(new_n335), .A3(new_n353), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n353), .B1(new_n333), .B2(new_n335), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(G101), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n355), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT76), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n355), .B(new_n367), .C1(new_n362), .C2(new_n364), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G122), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n355), .B(new_n369), .C1(new_n362), .C2(new_n364), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n372), .A2(KEYINPUT6), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT77), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n371), .A2(KEYINPUT6), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n377), .A3(new_n373), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n268), .A2(G143), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n215), .A2(G146), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n215), .C2(G146), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G128), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT66), .B1(new_n379), .B2(KEYINPUT1), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT65), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n215), .B2(G146), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n268), .A2(KEYINPUT65), .A3(G143), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .A4(new_n380), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n263), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G143), .B(G146), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT0), .B(G128), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT64), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(KEYINPUT0), .A2(G128), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n387), .A2(new_n388), .A3(new_n380), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(KEYINPUT0), .A2(G128), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT64), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n381), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n394), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n391), .B1(new_n401), .B2(new_n263), .ZN(new_n402));
  INV_X1    g216(.A(G224), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n375), .A2(new_n376), .A3(new_n378), .A4(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT78), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n402), .B1(new_n407), .B2(KEYINPUT7), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(new_n403), .B2(G953), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n372), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n340), .A2(new_n354), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n343), .A2(new_n348), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n355), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n369), .B(KEYINPUT8), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(G902), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n406), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n406), .A2(new_n418), .A3(new_n420), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n332), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n401), .A2(new_n426), .A3(new_n359), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n387), .A2(new_n388), .A3(new_n380), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n195), .B1(new_n379), .B2(KEYINPUT1), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n390), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n349), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT10), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT11), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n199), .B2(G137), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n199), .A2(G137), .ZN(new_n436));
  INV_X1    g250(.A(G137), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT11), .A3(G134), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G131), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n435), .A2(new_n438), .A3(new_n290), .A4(new_n436), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n385), .A2(new_n390), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT10), .A3(new_n349), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n427), .A2(new_n433), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G140), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n192), .A2(G227), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n385), .A2(new_n390), .A3(new_n413), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n385), .A2(new_n413), .A3(KEYINPUT75), .A4(new_n390), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n431), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n442), .A2(KEYINPUT74), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n460), .A3(new_n456), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n450), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n427), .A2(new_n433), .A3(new_n444), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n440), .A2(new_n441), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n449), .B1(new_n467), .B2(new_n445), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n425), .B(new_n257), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n445), .A2(new_n449), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n467), .ZN(new_n471));
  INV_X1    g285(.A(new_n445), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n462), .B2(new_n463), .ZN(new_n473));
  OAI211_X1 g287(.A(G469), .B(new_n471), .C1(new_n473), .C2(new_n449), .ZN(new_n474));
  NAND2_X1  g288(.A1(G469), .A2(G902), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G221), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n191), .B2(new_n257), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n330), .A2(new_n424), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT23), .B1(new_n195), .B2(G119), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT72), .B1(new_n195), .B2(G119), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G119), .B(G128), .ZN(new_n486));
  XOR2_X1   g300(.A(KEYINPUT24), .B(G110), .Z(new_n487));
  OAI22_X1  g301(.A1(new_n485), .A2(G110), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n299), .A3(new_n269), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n298), .A2(new_n299), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n486), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n485), .A2(G110), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT22), .B(G137), .ZN(new_n495));
  INV_X1    g309(.A(G234), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n477), .A2(new_n496), .A3(G953), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n495), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n498), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n489), .A2(new_n493), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G217), .B1(new_n496), .B2(G902), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT71), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n502), .A2(G902), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT25), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n499), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n506), .A2(new_n507), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n504), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n505), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n360), .A2(new_n361), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n394), .A2(new_n396), .A3(new_n400), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n442), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n437), .A2(G134), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n199), .A2(G137), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n441), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n385), .B2(new_n390), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n517), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT69), .ZN(new_n526));
  INV_X1    g340(.A(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n443), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n466), .A2(new_n396), .A3(new_n400), .A4(new_n394), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n516), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT69), .B(new_n517), .C1(new_n519), .C2(new_n524), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(KEYINPUT28), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n273), .A2(G210), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT27), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT26), .B(G101), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n401), .A2(new_n466), .B1(new_n443), .B2(new_n527), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT28), .B1(new_n538), .B2(new_n516), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n533), .A2(KEYINPUT29), .A3(new_n537), .A4(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT29), .ZN(new_n542));
  INV_X1    g356(.A(new_n530), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT30), .B1(new_n519), .B2(new_n524), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT30), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n528), .A2(new_n529), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n543), .B1(new_n547), .B2(new_n517), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(new_n548), .B2(new_n537), .ZN(new_n549));
  INV_X1    g363(.A(new_n537), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n516), .B1(new_n528), .B2(new_n529), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(KEYINPUT68), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n525), .A2(new_n554), .A3(new_n530), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n550), .B(new_n539), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n257), .B(new_n541), .C1(new_n549), .C2(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n557), .A2(KEYINPUT70), .A3(G472), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT70), .B1(new_n557), .B2(G472), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n519), .A2(KEYINPUT30), .A3(new_n524), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n545), .B1(new_n528), .B2(new_n529), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n517), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n537), .A3(new_n530), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT31), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n548), .A2(new_n566), .A3(new_n537), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n539), .B1(new_n553), .B2(new_n555), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n565), .B(new_n567), .C1(new_n537), .C2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(G472), .A2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT32), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT32), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n515), .B1(new_n560), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n482), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  NAND3_X1  g392(.A1(new_n476), .A2(new_n514), .A3(new_n479), .ZN(new_n579));
  INV_X1    g393(.A(new_n571), .ZN(new_n580));
  INV_X1    g394(.A(G472), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n569), .B2(new_n257), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n583), .B(KEYINPUT86), .Z(new_n584));
  AND3_X1   g398(.A1(new_n406), .A2(new_n418), .A3(new_n420), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n420), .B1(new_n406), .B2(new_n418), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n331), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n252), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT87), .B1(new_n232), .B2(new_n234), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  OAI22_X1  g404(.A1(new_n244), .A2(new_n235), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT87), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n253), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n255), .A3(new_n254), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n591), .A2(new_n594), .A3(G478), .A4(new_n257), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT88), .B(G478), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n245), .B2(G902), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n323), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n587), .A2(new_n588), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n584), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT34), .B(G104), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  INV_X1    g417(.A(new_n327), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n328), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n587), .A2(new_n588), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n584), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT89), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT35), .B(G107), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  NOR2_X1   g424(.A1(new_n587), .A2(new_n480), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n569), .A2(new_n257), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n612), .A2(G472), .B1(new_n569), .B2(new_n570), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n511), .A2(new_n513), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n498), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n494), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n257), .A3(new_n512), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n324), .B2(new_n329), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n611), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT37), .B(G110), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT90), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT91), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n621), .B(new_n624), .ZN(G12));
  NAND2_X1  g439(.A1(new_n557), .A2(G472), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT70), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n557), .A2(KEYINPUT70), .A3(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n573), .B1(new_n569), .B2(new_n570), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n569), .A2(new_n573), .A3(new_n570), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n248), .B(KEYINPUT92), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(G900), .B2(new_n251), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT93), .Z(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n604), .A2(new_n328), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n476), .A2(new_n618), .A3(new_n479), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n632), .A2(new_n424), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  XOR2_X1   g455(.A(new_n635), .B(KEYINPUT39), .Z(new_n642));
  AND2_X1   g456(.A1(new_n481), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT40), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n422), .A2(new_n423), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT38), .Z(new_n646));
  NAND2_X1  g460(.A1(new_n531), .A2(new_n532), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n550), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n516), .B1(new_n544), .B2(new_n546), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n537), .B1(new_n649), .B2(new_n543), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n257), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(G472), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT94), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT94), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n651), .A2(new_n654), .A3(G472), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n631), .B2(new_n630), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n327), .A2(new_n328), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n331), .A3(new_n619), .A4(new_n658), .ZN(new_n659));
  OR3_X1    g473(.A1(new_n644), .A2(new_n646), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT95), .B(G143), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G45));
  NAND3_X1  g476(.A1(new_n598), .A2(new_n323), .A3(new_n636), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n638), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n632), .A2(new_n424), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT96), .B(G146), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G48));
  OAI21_X1  g481(.A(new_n257), .B1(new_n464), .B2(new_n468), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G469), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n479), .A3(new_n469), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT97), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT97), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n669), .A2(new_n672), .A3(new_n479), .A4(new_n469), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n576), .A2(new_n600), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND3_X1  g491(.A1(new_n576), .A2(new_n606), .A3(new_n674), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  NAND4_X1  g493(.A1(new_n674), .A2(new_n632), .A3(new_n424), .A4(new_n620), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  OAI211_X1 g495(.A(new_n658), .B(new_n331), .C1(new_n585), .C2(new_n586), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT100), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n645), .A2(new_n684), .A3(new_n331), .A4(new_n658), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n671), .A2(new_n252), .A3(new_n673), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n533), .A2(new_n540), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT99), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n533), .A2(new_n540), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n550), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n565), .A2(new_n567), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n570), .B(KEYINPUT98), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n612), .A2(G472), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n514), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n687), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n686), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n686), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND3_X1  g520(.A1(new_n424), .A2(new_n673), .A3(new_n671), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n598), .A2(new_n323), .A3(new_n636), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n698), .A3(new_n618), .A4(new_n697), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n263), .ZN(G27));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n422), .A2(new_n331), .A3(new_n423), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n470), .A2(KEYINPUT102), .A3(new_n467), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n465), .A2(new_n466), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n715), .B1(new_n716), .B2(new_n450), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n714), .B(new_n717), .C1(new_n473), .C2(new_n449), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n469), .B(new_n475), .C1(new_n718), .C2(new_n425), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT103), .B1(new_n719), .B2(new_n479), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(KEYINPUT103), .A3(new_n479), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n632), .A3(new_n514), .A4(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n712), .B1(new_n723), .B2(new_n663), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n479), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n585), .A2(new_n586), .A3(new_n332), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n722), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n576), .A3(KEYINPUT42), .A4(new_n708), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  OAI21_X1  g546(.A(KEYINPUT104), .B1(new_n723), .B2(new_n637), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  INV_X1    g548(.A(new_n637), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n729), .A2(new_n576), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT105), .B(G134), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G36));
  NAND2_X1  g553(.A1(new_n598), .A2(new_n328), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT43), .ZN(new_n741));
  OR3_X1    g555(.A1(new_n741), .A2(new_n613), .A3(new_n619), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT106), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n473), .A2(new_n449), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n471), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n749), .B(G469), .C1(new_n748), .C2(new_n718), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n475), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n475), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n469), .A3(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n479), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(new_n642), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n713), .B1(new_n742), .B2(new_n743), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n745), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  XNOR2_X1  g574(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n632), .A2(new_n514), .A3(new_n663), .A4(new_n713), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT47), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n763), .B(new_n764), .C1(new_n756), .C2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  NAND2_X1  g584(.A1(new_n674), .A2(new_n728), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n771), .A2(new_n515), .A3(new_n248), .A4(new_n657), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT118), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n773), .A2(new_n323), .A3(new_n598), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n741), .A2(new_n633), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(new_n771), .ZN(new_n776));
  INV_X1    g590(.A(new_n696), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n692), .B2(new_n694), .ZN(new_n778));
  OR4_X1    g592(.A1(new_n582), .A2(new_n776), .A3(new_n619), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n674), .A2(new_n332), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT116), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n775), .A2(new_n699), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n646), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT50), .Z(new_n786));
  NAND3_X1  g600(.A1(new_n669), .A2(new_n478), .A3(new_n469), .ZN(new_n787));
  INV_X1    g601(.A(new_n763), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n756), .A2(new_n766), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n775), .A2(new_n699), .A3(new_n713), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n786), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n576), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n776), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT48), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n773), .A2(new_n599), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n192), .A2(G952), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n775), .A2(new_n707), .A3(new_n699), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n787), .B(KEYINPUT115), .Z(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n788), .B2(new_n789), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n791), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n781), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n786), .B(KEYINPUT117), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n793), .B(new_n800), .C1(new_n806), .C2(KEYINPUT51), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n325), .B2(new_n326), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n246), .A2(KEYINPUT110), .A3(new_n259), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n638), .A2(new_n811), .A3(new_n323), .A4(new_n635), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n632), .A2(new_n812), .A3(new_n728), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n663), .A2(new_n778), .A3(new_n582), .A4(new_n619), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n729), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n727), .A2(new_n728), .A3(new_n722), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n709), .A3(KEYINPUT111), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n813), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n640), .B1(new_n707), .B2(new_n709), .ZN(new_n820));
  INV_X1    g634(.A(new_n725), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n618), .A2(new_n635), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n657), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n685), .B2(new_n683), .ZN(new_n824));
  INV_X1    g638(.A(new_n665), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n820), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n819), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n330), .A2(new_n613), .A3(new_n618), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n576), .A2(new_n482), .B1(new_n829), .B2(new_n611), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n576), .B(new_n674), .C1(new_n600), .C2(new_n606), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n811), .A2(new_n328), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n599), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n583), .A2(new_n833), .A3(new_n252), .A4(new_n424), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n830), .A2(new_n831), .A3(new_n680), .A4(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n686), .A2(new_n703), .A3(new_n700), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n703), .B1(new_n686), .B2(new_n700), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n724), .A2(new_n730), .B1(new_n733), .B2(new_n736), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n686), .A2(new_n657), .A3(new_n821), .A4(new_n822), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n665), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT52), .B1(new_n842), .B2(new_n820), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n828), .A2(new_n839), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  OR3_X1    g659(.A1(new_n844), .A2(KEYINPUT113), .A3(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n577), .A2(new_n621), .A3(new_n680), .A4(new_n834), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n705), .A2(new_n847), .A3(new_n831), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n731), .A2(new_n737), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n850), .A2(new_n828), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n632), .A2(new_n424), .A3(new_n639), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT112), .B1(new_n852), .B2(new_n710), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n815), .A2(new_n424), .A3(new_n674), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n855), .A3(new_n640), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n665), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT52), .B1(new_n857), .B2(new_n824), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT113), .B1(new_n844), .B2(new_n845), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n846), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n844), .A2(new_n845), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n828), .A4(new_n858), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n861), .A2(new_n862), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n807), .A2(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n669), .A2(new_n469), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(KEYINPUT49), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT109), .Z(new_n872));
  INV_X1    g686(.A(new_n657), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n514), .A2(new_n331), .A3(new_n479), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n874), .B(new_n740), .C1(KEYINPUT49), .C2(new_n870), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n646), .A2(new_n872), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n876), .ZN(G75));
  NOR2_X1   g691(.A1(new_n192), .A2(G952), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n257), .B1(new_n865), .B2(new_n866), .ZN(new_n880));
  AOI211_X1 g694(.A(KEYINPUT119), .B(KEYINPUT56), .C1(new_n880), .C2(G210), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n405), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT55), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n879), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n884), .B2(new_n881), .ZN(G51));
  XNOR2_X1  g700(.A(new_n867), .B(new_n864), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n475), .B(KEYINPUT57), .Z(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n464), .B2(new_n468), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n750), .B(KEYINPUT120), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n878), .B1(new_n890), .B2(new_n892), .ZN(G54));
  NAND3_X1  g707(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  INV_X1    g708(.A(new_n312), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n878), .ZN(G60));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT59), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n887), .A2(new_n591), .A3(new_n594), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n879), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n868), .A2(new_n900), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n591), .A2(new_n594), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n867), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT122), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n867), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n502), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n867), .B2(new_n908), .ZN(new_n914));
  AOI211_X1 g728(.A(KEYINPUT122), .B(new_n907), .C1(new_n865), .C2(new_n866), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n616), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n916), .A3(new_n879), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n917), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT61), .B1(new_n917), .B2(KEYINPUT121), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(G66));
  INV_X1    g734(.A(new_n250), .ZN(new_n921));
  OAI21_X1  g735(.A(G953), .B1(new_n921), .B2(new_n403), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n839), .B2(G953), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT123), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n882), .B1(G898), .B2(new_n192), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(G69));
  AOI21_X1  g740(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n305), .B1(new_n267), .B2(new_n306), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT124), .Z(new_n931));
  XNOR2_X1  g745(.A(new_n547), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n857), .B(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n660), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n576), .A2(new_n643), .A3(new_n728), .A4(new_n833), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n759), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n769), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n932), .B1(new_n939), .B2(new_n192), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n757), .A2(new_n576), .A3(new_n686), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n759), .A2(new_n840), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n769), .A3(new_n933), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(G953), .ZN(new_n944));
  INV_X1    g758(.A(G900), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n932), .B1(new_n945), .B2(new_n192), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n929), .B1(new_n940), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n927), .A2(new_n928), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT127), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n929), .B(new_n950), .C1(new_n940), .C2(new_n947), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G72));
  OR2_X1    g768(.A1(new_n939), .A2(new_n848), .ZN(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  AOI21_X1  g771(.A(new_n650), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n943), .B2(new_n848), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n649), .A2(new_n537), .A3(new_n543), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n878), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n548), .A2(new_n537), .ZN(new_n962));
  INV_X1    g776(.A(new_n564), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n861), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n958), .A2(new_n965), .ZN(G57));
endmodule


