

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(G651), .A2(n567), .ZN(n791) );
  NAND2_X2 U552 ( .A1(n702), .A2(n595), .ZN(n650) );
  OR2_X1 U553 ( .A1(n634), .A2(n928), .ZN(n633) );
  XNOR2_X1 U554 ( .A(n521), .B(n520), .ZN(n586) );
  XNOR2_X1 U555 ( .A(n519), .B(KEYINPUT17), .ZN(n520) );
  INV_X1 U556 ( .A(KEYINPUT66), .ZN(n519) );
  INV_X1 U557 ( .A(KEYINPUT26), .ZN(n600) );
  INV_X1 U558 ( .A(KEYINPUT13), .ZN(n608) );
  XNOR2_X1 U559 ( .A(n608), .B(KEYINPUT75), .ZN(n609) );
  XNOR2_X1 U560 ( .A(n610), .B(n609), .ZN(n614) );
  NAND2_X1 U561 ( .A1(n749), .A2(n594), .ZN(n701) );
  XNOR2_X1 U562 ( .A(G651), .B(KEYINPUT69), .ZN(n534) );
  INV_X1 U563 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U564 ( .A1(n525), .A2(G2104), .ZN(n517) );
  XNOR2_X1 U565 ( .A(n517), .B(KEYINPUT65), .ZN(n592) );
  INV_X1 U566 ( .A(n592), .ZN(n518) );
  INV_X1 U567 ( .A(n518), .ZN(n886) );
  NAND2_X1 U568 ( .A1(n886), .A2(G102), .ZN(n524) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  INV_X1 U570 ( .A(n586), .ZN(n522) );
  INV_X1 U571 ( .A(n522), .ZN(n884) );
  NAND2_X1 U572 ( .A1(G138), .A2(n884), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n524), .A2(n523), .ZN(n529) );
  NOR2_X2 U574 ( .A1(G2104), .A2(n525), .ZN(n878) );
  NAND2_X1 U575 ( .A1(G126), .A2(n878), .ZN(n527) );
  AND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U577 ( .A1(G114), .A2(n879), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U579 ( .A1(n529), .A2(n528), .ZN(G164) );
  XOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .Z(n567) );
  NAND2_X1 U581 ( .A1(G52), .A2(n791), .ZN(n533) );
  NOR2_X1 U582 ( .A1(G543), .A2(n534), .ZN(n531) );
  XOR2_X1 U583 ( .A(KEYINPUT70), .B(KEYINPUT1), .Z(n530) );
  XNOR2_X2 U584 ( .A(n531), .B(n530), .ZN(n795) );
  NAND2_X1 U585 ( .A1(G64), .A2(n795), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n541) );
  XNOR2_X1 U587 ( .A(KEYINPUT9), .B(KEYINPUT72), .ZN(n539) );
  NOR2_X2 U588 ( .A1(n567), .A2(n534), .ZN(n792) );
  NAND2_X1 U589 ( .A1(G77), .A2(n792), .ZN(n537) );
  NOR2_X1 U590 ( .A1(G543), .A2(G651), .ZN(n796) );
  NAND2_X1 U591 ( .A1(n796), .A2(G90), .ZN(n535) );
  XOR2_X1 U592 ( .A(KEYINPUT71), .B(n535), .Z(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U594 ( .A(n539), .B(n538), .Z(n540) );
  NOR2_X1 U595 ( .A1(n541), .A2(n540), .ZN(G171) );
  INV_X1 U596 ( .A(G171), .ZN(G301) );
  NAND2_X1 U597 ( .A1(G51), .A2(n791), .ZN(n543) );
  NAND2_X1 U598 ( .A1(G63), .A2(n795), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U600 ( .A(KEYINPUT6), .B(n544), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n796), .A2(G89), .ZN(n545) );
  XNOR2_X1 U602 ( .A(n545), .B(KEYINPUT4), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G76), .A2(n792), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT5), .B(n548), .Z(n549) );
  XNOR2_X1 U606 ( .A(KEYINPUT80), .B(n549), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U608 ( .A(KEYINPUT7), .B(n552), .Z(G168) );
  XOR2_X1 U609 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U610 ( .A1(n796), .A2(G88), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G75), .A2(n792), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G50), .A2(n791), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G62), .A2(n795), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(G166) );
  INV_X1 U617 ( .A(G166), .ZN(G303) );
  XOR2_X1 U618 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n560) );
  NAND2_X1 U619 ( .A1(G73), .A2(n792), .ZN(n559) );
  XNOR2_X1 U620 ( .A(n560), .B(n559), .ZN(n564) );
  NAND2_X1 U621 ( .A1(G48), .A2(n791), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G86), .A2(n796), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n795), .A2(G61), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(G305) );
  NAND2_X1 U627 ( .A1(G87), .A2(n567), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G74), .A2(G651), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U630 ( .A1(n795), .A2(n570), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n791), .A2(G49), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U633 ( .A1(n791), .A2(G47), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G72), .A2(n792), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n796), .A2(G85), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT68), .B(n575), .Z(n576) );
  NOR2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n795), .A2(G60), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G290) );
  NAND2_X1 U641 ( .A1(G53), .A2(n791), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G65), .A2(n795), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n796), .A2(G91), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G78), .A2(n792), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n804) );
  NOR2_X1 U648 ( .A1(G164), .A2(G1384), .ZN(n702) );
  NAND2_X1 U649 ( .A1(G137), .A2(n586), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n879), .A2(G113), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U652 ( .A(n589), .B(KEYINPUT67), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G125), .A2(n878), .ZN(n590) );
  AND2_X1 U654 ( .A1(n591), .A2(n590), .ZN(n749) );
  NAND2_X1 U655 ( .A1(G101), .A2(n592), .ZN(n593) );
  XOR2_X1 U656 ( .A(KEYINPUT23), .B(n593), .Z(n750) );
  AND2_X1 U657 ( .A1(G40), .A2(n750), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT90), .B(n701), .Z(n595) );
  INV_X1 U659 ( .A(n650), .ZN(n645) );
  NAND2_X1 U660 ( .A1(n645), .A2(G2072), .ZN(n596) );
  XNOR2_X1 U661 ( .A(n596), .B(KEYINPUT27), .ZN(n598) );
  INV_X1 U662 ( .A(G1956), .ZN(n939) );
  NOR2_X1 U663 ( .A1(n939), .A2(n645), .ZN(n597) );
  NOR2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n637) );
  OR2_X1 U665 ( .A1(n804), .A2(n637), .ZN(n599) );
  XNOR2_X1 U666 ( .A(KEYINPUT28), .B(n599), .ZN(n642) );
  XOR2_X1 U667 ( .A(G1996), .B(KEYINPUT94), .Z(n1003) );
  NOR2_X1 U668 ( .A1(n650), .A2(n1003), .ZN(n601) );
  XNOR2_X1 U669 ( .A(n601), .B(n600), .ZN(n603) );
  NAND2_X1 U670 ( .A1(n650), .A2(G1341), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n618) );
  NAND2_X1 U672 ( .A1(G43), .A2(n791), .ZN(n616) );
  NAND2_X1 U673 ( .A1(n796), .A2(G81), .ZN(n604) );
  XOR2_X1 U674 ( .A(KEYINPUT12), .B(n604), .Z(n607) );
  NAND2_X1 U675 ( .A1(G68), .A2(n792), .ZN(n605) );
  XOR2_X1 U676 ( .A(n605), .B(KEYINPUT74), .Z(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G56), .A2(n795), .ZN(n611) );
  XNOR2_X1 U679 ( .A(n611), .B(KEYINPUT14), .ZN(n612) );
  XNOR2_X1 U680 ( .A(KEYINPUT73), .B(n612), .ZN(n613) );
  NOR2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U682 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X2 U683 ( .A(n617), .B(KEYINPUT76), .ZN(n929) );
  NOR2_X1 U684 ( .A1(n618), .A2(n929), .ZN(n620) );
  INV_X1 U685 ( .A(KEYINPUT64), .ZN(n619) );
  XNOR2_X1 U686 ( .A(n620), .B(n619), .ZN(n634) );
  NAND2_X1 U687 ( .A1(n791), .A2(G54), .ZN(n622) );
  NAND2_X1 U688 ( .A1(G79), .A2(n792), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U690 ( .A1(G66), .A2(n795), .ZN(n624) );
  NAND2_X1 U691 ( .A1(G92), .A2(n796), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U693 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U694 ( .A(KEYINPUT15), .B(n627), .Z(n628) );
  XNOR2_X1 U695 ( .A(KEYINPUT78), .B(n628), .ZN(n789) );
  AND2_X1 U696 ( .A1(n650), .A2(G1348), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n629), .B(KEYINPUT95), .ZN(n631) );
  NAND2_X1 U698 ( .A1(n645), .A2(G2067), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n636) );
  INV_X1 U701 ( .A(n789), .ZN(n928) );
  NAND2_X1 U702 ( .A1(n928), .A2(n634), .ZN(n635) );
  NAND2_X1 U703 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U704 ( .A1(n804), .A2(n637), .ZN(n638) );
  NAND2_X1 U705 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U706 ( .A(KEYINPUT96), .B(n640), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U708 ( .A(KEYINPUT29), .B(n643), .ZN(n649) );
  NAND2_X1 U709 ( .A1(G1961), .A2(n650), .ZN(n647) );
  XNOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n644), .B(KEYINPUT93), .ZN(n1002) );
  NAND2_X1 U712 ( .A1(n645), .A2(n1002), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n654) );
  NOR2_X1 U714 ( .A1(G301), .A2(n654), .ZN(n648) );
  NOR2_X1 U715 ( .A1(n649), .A2(n648), .ZN(n659) );
  NAND2_X1 U716 ( .A1(G8), .A2(n650), .ZN(n694) );
  NOR2_X1 U717 ( .A1(G1966), .A2(n694), .ZN(n670) );
  NOR2_X1 U718 ( .A1(G2084), .A2(n650), .ZN(n671) );
  NOR2_X1 U719 ( .A1(n670), .A2(n671), .ZN(n651) );
  NAND2_X1 U720 ( .A1(G8), .A2(n651), .ZN(n652) );
  XNOR2_X1 U721 ( .A(KEYINPUT30), .B(n652), .ZN(n653) );
  NOR2_X1 U722 ( .A1(G168), .A2(n653), .ZN(n656) );
  AND2_X1 U723 ( .A1(G301), .A2(n654), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(KEYINPUT31), .ZN(n658) );
  NOR2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n669) );
  INV_X1 U727 ( .A(n669), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n660), .A2(G286), .ZN(n666) );
  NOR2_X1 U729 ( .A1(G1971), .A2(n694), .ZN(n662) );
  NOR2_X1 U730 ( .A1(G2090), .A2(n650), .ZN(n661) );
  NOR2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n663), .A2(G303), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(KEYINPUT98), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U735 ( .A1(n667), .A2(G8), .ZN(n668) );
  XNOR2_X1 U736 ( .A(KEYINPUT32), .B(n668), .ZN(n676) );
  NOR2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n673) );
  NAND2_X1 U738 ( .A1(G8), .A2(n671), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U740 ( .A(n674), .B(KEYINPUT97), .Z(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n689) );
  NAND2_X1 U742 ( .A1(G166), .A2(G8), .ZN(n677) );
  OR2_X1 U743 ( .A1(G2090), .A2(n677), .ZN(n678) );
  AND2_X1 U744 ( .A1(n689), .A2(n678), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n679), .B(KEYINPUT99), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n680), .A2(n694), .ZN(n686) );
  NOR2_X1 U747 ( .A1(G1981), .A2(G305), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(KEYINPUT91), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT24), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n683), .A2(n694), .ZN(n684) );
  XOR2_X1 U751 ( .A(n684), .B(KEYINPUT92), .Z(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n700) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n917) );
  NOR2_X1 U755 ( .A1(n687), .A2(n917), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n918) );
  INV_X1 U758 ( .A(n918), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n690), .A2(n694), .ZN(n691) );
  AND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U761 ( .A1(KEYINPUT33), .A2(n693), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n917), .A2(KEYINPUT33), .ZN(n695) );
  OR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U764 ( .A(G1981), .B(G305), .Z(n914) );
  NAND2_X1 U765 ( .A1(n696), .A2(n914), .ZN(n697) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n730) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n744) );
  NAND2_X1 U769 ( .A1(G105), .A2(n886), .ZN(n703) );
  XNOR2_X1 U770 ( .A(n703), .B(KEYINPUT38), .ZN(n711) );
  NAND2_X1 U771 ( .A1(n878), .A2(G129), .ZN(n704) );
  XNOR2_X1 U772 ( .A(n704), .B(KEYINPUT88), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G117), .A2(n879), .ZN(n705) );
  NAND2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U775 ( .A1(G141), .A2(n884), .ZN(n707) );
  XNOR2_X1 U776 ( .A(KEYINPUT89), .B(n707), .ZN(n708) );
  NOR2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n873) );
  NAND2_X1 U779 ( .A1(G1996), .A2(n873), .ZN(n719) );
  NAND2_X1 U780 ( .A1(n878), .A2(G119), .ZN(n713) );
  NAND2_X1 U781 ( .A1(G131), .A2(n884), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U783 ( .A1(G95), .A2(n886), .ZN(n715) );
  NAND2_X1 U784 ( .A1(G107), .A2(n879), .ZN(n714) );
  NAND2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n716) );
  OR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n894) );
  NAND2_X1 U787 ( .A1(G1991), .A2(n894), .ZN(n718) );
  NAND2_X1 U788 ( .A1(n719), .A2(n718), .ZN(n977) );
  NAND2_X1 U789 ( .A1(n744), .A2(n977), .ZN(n737) );
  XNOR2_X1 U790 ( .A(KEYINPUT37), .B(G2067), .ZN(n733) );
  NAND2_X1 U791 ( .A1(n886), .A2(G104), .ZN(n721) );
  NAND2_X1 U792 ( .A1(G140), .A2(n884), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U794 ( .A(KEYINPUT34), .B(n722), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G128), .A2(n878), .ZN(n724) );
  NAND2_X1 U796 ( .A1(G116), .A2(n879), .ZN(n723) );
  NAND2_X1 U797 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U798 ( .A(KEYINPUT35), .B(n725), .Z(n726) );
  NOR2_X1 U799 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U800 ( .A(KEYINPUT36), .B(n728), .ZN(n896) );
  NOR2_X1 U801 ( .A1(n733), .A2(n896), .ZN(n968) );
  NAND2_X1 U802 ( .A1(n744), .A2(n968), .ZN(n741) );
  NAND2_X1 U803 ( .A1(n737), .A2(n741), .ZN(n729) );
  NOR2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n923) );
  NAND2_X1 U806 ( .A1(n923), .A2(n744), .ZN(n731) );
  NAND2_X1 U807 ( .A1(n732), .A2(n731), .ZN(n747) );
  NAND2_X1 U808 ( .A1(n733), .A2(n896), .ZN(n970) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n734) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n894), .ZN(n979) );
  NOR2_X1 U811 ( .A1(n734), .A2(n979), .ZN(n735) );
  XOR2_X1 U812 ( .A(KEYINPUT100), .B(n735), .Z(n736) );
  NAND2_X1 U813 ( .A1(n737), .A2(n736), .ZN(n738) );
  OR2_X1 U814 ( .A1(n873), .A2(G1996), .ZN(n985) );
  NAND2_X1 U815 ( .A1(n738), .A2(n985), .ZN(n740) );
  XNOR2_X1 U816 ( .A(KEYINPUT101), .B(KEYINPUT39), .ZN(n739) );
  XNOR2_X1 U817 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U818 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U819 ( .A1(n970), .A2(n743), .ZN(n745) );
  NAND2_X1 U820 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U822 ( .A(n748), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U823 ( .A1(n749), .A2(n750), .ZN(G160) );
  XNOR2_X1 U824 ( .A(G2451), .B(G2446), .ZN(n760) );
  XOR2_X1 U825 ( .A(G2430), .B(KEYINPUT103), .Z(n752) );
  XNOR2_X1 U826 ( .A(G2454), .B(G2435), .ZN(n751) );
  XNOR2_X1 U827 ( .A(n752), .B(n751), .ZN(n756) );
  XOR2_X1 U828 ( .A(G2438), .B(KEYINPUT102), .Z(n754) );
  XNOR2_X1 U829 ( .A(G1348), .B(G1341), .ZN(n753) );
  XNOR2_X1 U830 ( .A(n754), .B(n753), .ZN(n755) );
  XOR2_X1 U831 ( .A(n756), .B(n755), .Z(n758) );
  XNOR2_X1 U832 ( .A(G2443), .B(G2427), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U834 ( .A(n760), .B(n759), .ZN(n761) );
  AND2_X1 U835 ( .A1(n761), .A2(G14), .ZN(G401) );
  AND2_X1 U836 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U837 ( .A(G57), .ZN(G237) );
  INV_X1 U838 ( .A(G132), .ZN(G219) );
  INV_X1 U839 ( .A(G82), .ZN(G220) );
  NAND2_X1 U840 ( .A1(G7), .A2(G661), .ZN(n762) );
  XNOR2_X1 U841 ( .A(n762), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U842 ( .A(G223), .ZN(n829) );
  NAND2_X1 U843 ( .A1(n829), .A2(G567), .ZN(n763) );
  XOR2_X1 U844 ( .A(KEYINPUT11), .B(n763), .Z(G234) );
  XOR2_X1 U845 ( .A(G860), .B(KEYINPUT77), .Z(n771) );
  INV_X1 U846 ( .A(n929), .ZN(n764) );
  NAND2_X1 U847 ( .A1(n771), .A2(n764), .ZN(G153) );
  NOR2_X1 U848 ( .A1(G868), .A2(n789), .ZN(n765) );
  XNOR2_X1 U849 ( .A(n765), .B(KEYINPUT79), .ZN(n767) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n767), .A2(n766), .ZN(G284) );
  INV_X1 U852 ( .A(n804), .ZN(G299) );
  INV_X1 U853 ( .A(G868), .ZN(n811) );
  NOR2_X1 U854 ( .A1(G286), .A2(n811), .ZN(n769) );
  NOR2_X1 U855 ( .A1(G868), .A2(G299), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(G297) );
  INV_X1 U857 ( .A(G559), .ZN(n770) );
  NOR2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT81), .B(n772), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n773), .A2(n789), .ZN(n774) );
  XNOR2_X1 U861 ( .A(n774), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U862 ( .A1(n929), .A2(G868), .ZN(n775) );
  XNOR2_X1 U863 ( .A(KEYINPUT82), .B(n775), .ZN(n778) );
  NAND2_X1 U864 ( .A1(G868), .A2(n789), .ZN(n776) );
  NOR2_X1 U865 ( .A1(G559), .A2(n776), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(G282) );
  NAND2_X1 U867 ( .A1(G123), .A2(n878), .ZN(n779) );
  XOR2_X1 U868 ( .A(KEYINPUT83), .B(n779), .Z(n780) );
  XNOR2_X1 U869 ( .A(n780), .B(KEYINPUT18), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G111), .A2(n879), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n886), .A2(G99), .ZN(n784) );
  NAND2_X1 U873 ( .A1(G135), .A2(n884), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n978) );
  XNOR2_X1 U876 ( .A(n978), .B(G2096), .ZN(n788) );
  INV_X1 U877 ( .A(G2100), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(G156) );
  NAND2_X1 U879 ( .A1(n789), .A2(G559), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n790), .B(n929), .ZN(n809) );
  NOR2_X1 U881 ( .A1(G860), .A2(n809), .ZN(n801) );
  NAND2_X1 U882 ( .A1(n791), .A2(G55), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n800) );
  NAND2_X1 U885 ( .A1(G67), .A2(n795), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G93), .A2(n796), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n812) );
  XOR2_X1 U889 ( .A(n801), .B(n812), .Z(G145) );
  XOR2_X1 U890 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n802) );
  XNOR2_X1 U891 ( .A(G288), .B(n802), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n804), .B(n803), .ZN(n806) );
  XNOR2_X1 U893 ( .A(G290), .B(G166), .ZN(n805) );
  XNOR2_X1 U894 ( .A(n806), .B(n805), .ZN(n807) );
  XNOR2_X1 U895 ( .A(n812), .B(n807), .ZN(n808) );
  XNOR2_X1 U896 ( .A(G305), .B(n808), .ZN(n900) );
  XOR2_X1 U897 ( .A(n900), .B(n809), .Z(n810) );
  NOR2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n814) );
  NOR2_X1 U899 ( .A1(G868), .A2(n812), .ZN(n813) );
  NOR2_X1 U900 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U907 ( .A1(G220), .A2(G219), .ZN(n819) );
  XOR2_X1 U908 ( .A(KEYINPUT22), .B(n819), .Z(n820) );
  NOR2_X1 U909 ( .A1(G218), .A2(n820), .ZN(n821) );
  XNOR2_X1 U910 ( .A(KEYINPUT86), .B(n821), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n822), .A2(G96), .ZN(n833) );
  NAND2_X1 U912 ( .A1(n833), .A2(G2106), .ZN(n826) );
  NAND2_X1 U913 ( .A1(G69), .A2(G120), .ZN(n823) );
  NOR2_X1 U914 ( .A1(G237), .A2(n823), .ZN(n824) );
  NAND2_X1 U915 ( .A1(G108), .A2(n824), .ZN(n834) );
  NAND2_X1 U916 ( .A1(n834), .A2(G567), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n835) );
  NAND2_X1 U918 ( .A1(G483), .A2(G661), .ZN(n827) );
  NOR2_X1 U919 ( .A1(n835), .A2(n827), .ZN(n832) );
  NAND2_X1 U920 ( .A1(n832), .A2(G36), .ZN(n828) );
  XOR2_X1 U921 ( .A(KEYINPUT87), .B(n828), .Z(G176) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n835), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT43), .B(G2678), .Z(n837) );
  XNOR2_X1 U935 ( .A(KEYINPUT105), .B(KEYINPUT104), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT42), .B(G2090), .Z(n839) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2096), .B(G2100), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U943 ( .A(G2078), .B(G2084), .Z(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1956), .B(G1971), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1976), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n848), .B(G2474), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1981), .B(G1966), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1961), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U955 ( .A1(G124), .A2(n878), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n855), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n884), .A2(G136), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n856), .B(KEYINPUT106), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U960 ( .A1(G100), .A2(n886), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G112), .A2(n879), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U963 ( .A1(n862), .A2(n861), .ZN(G162) );
  NAND2_X1 U964 ( .A1(n886), .A2(G106), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G142), .A2(n884), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n865), .B(KEYINPUT45), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n879), .A2(G118), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT107), .B(n866), .Z(n868) );
  NAND2_X1 U970 ( .A1(n878), .A2(G130), .ZN(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U972 ( .A(KEYINPUT108), .B(n869), .Z(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n872), .B(G162), .ZN(n877) );
  XOR2_X1 U975 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n875) );
  XOR2_X1 U976 ( .A(n873), .B(KEYINPUT48), .Z(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U978 ( .A(n877), .B(n876), .Z(n892) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G127), .A2(n878), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G115), .A2(n879), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G139), .A2(n884), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n885), .B(KEYINPUT110), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n972) );
  XNOR2_X1 U989 ( .A(G164), .B(n972), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n898) );
  XOR2_X1 U991 ( .A(G160), .B(n978), .Z(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U995 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U996 ( .A(n900), .B(G286), .Z(n902) );
  XNOR2_X1 U997 ( .A(G171), .B(n928), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n903), .B(n929), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n904), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(KEYINPUT112), .B(n905), .ZN(G397) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n908), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n909), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT114), .B(n910), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(G16), .ZN(n964) );
  XNOR2_X1 U1013 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(n964), .B(n913), .ZN(n938) );
  XNOR2_X1 U1015 ( .A(G1966), .B(G168), .ZN(n915) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(KEYINPUT57), .B(n916), .ZN(n936) );
  XOR2_X1 U1018 ( .A(n917), .B(KEYINPUT122), .Z(n919) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n921) );
  XOR2_X1 U1020 ( .A(G1971), .B(G166), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G1956), .B(G299), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(G1961), .B(G301), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(G1348), .B(n928), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n929), .B(G1341), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(KEYINPUT123), .B(n934), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n966) );
  XOR2_X1 U1034 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n962) );
  XOR2_X1 U1035 ( .A(G1966), .B(G21), .Z(n949) );
  XNOR2_X1 U1036 ( .A(G20), .B(n939), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G1981), .B(G6), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(G1341), .B(G19), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1041 ( .A(KEYINPUT59), .B(G1348), .Z(n944) );
  XNOR2_X1 U1042 ( .A(G4), .B(n944), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT60), .B(n947), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT124), .B(G1961), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G5), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(G1986), .B(G24), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(G1971), .B(KEYINPUT125), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n955), .B(G22), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1055 ( .A(KEYINPUT58), .B(n958), .Z(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n962), .B(n961), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n967), .B(KEYINPUT127), .ZN(n998) );
  INV_X1 U1061 ( .A(n968), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n992) );
  XNOR2_X1 U1063 ( .A(G164), .B(G2078), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n971), .B(KEYINPUT117), .ZN(n974) );
  XOR2_X1 U1065 ( .A(G2072), .B(n972), .Z(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(KEYINPUT50), .B(n975), .ZN(n990) );
  XOR2_X1 U1068 ( .A(G160), .B(G2084), .Z(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n982) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1071 ( .A(KEYINPUT115), .B(n980), .Z(n981) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G2090), .B(G162), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n983), .B(KEYINPUT116), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n986), .Z(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1080 ( .A(KEYINPUT52), .B(n993), .Z(n994) );
  NOR2_X1 U1081 ( .A1(KEYINPUT55), .A2(n994), .ZN(n995) );
  XOR2_X1 U1082 ( .A(KEYINPUT118), .B(n995), .Z(n996) );
  NAND2_X1 U1083 ( .A1(n996), .A2(G29), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1022) );
  XNOR2_X1 U1085 ( .A(G1991), .B(G25), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G33), .B(G2072), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1009) );
  XOR2_X1 U1088 ( .A(G2067), .B(G26), .Z(n1001) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(G28), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(n1002), .B(G27), .Z(n1005) );
  XNOR2_X1 U1091 ( .A(n1003), .B(G32), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(n1010), .B(KEYINPUT53), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(G2084), .B(G34), .Z(n1011) );
  XNOR2_X1 U1097 ( .A(KEYINPUT54), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(G35), .B(G2090), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(n1016), .B(KEYINPUT55), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(G29), .B(KEYINPUT119), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(G11), .A2(n1019), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT120), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .ZN(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

