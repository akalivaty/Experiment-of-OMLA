//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(KEYINPUT67), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  INV_X1    g046(.A(new_n463), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(G160));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n479), .A2(new_n461), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(new_n487), .B2(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n461), .B2(G114), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G102), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n461), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n492), .A2(new_n494), .A3(G2104), .A4(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n479), .A2(new_n502), .A3(G138), .A4(new_n461), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT71), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT71), .A2(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT6), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n507), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n507), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT71), .B(G651), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n513), .A2(G88), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n510), .B2(new_n512), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  XNOR2_X1  g098(.A(KEYINPUT72), .B(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(G51), .ZN(new_n526));
  INV_X1    g101(.A(new_n507), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n527), .A2(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G168));
  XOR2_X1   g109(.A(KEYINPUT73), .B(G90), .Z(new_n535));
  NAND2_X1  g110(.A1(new_n513), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n520), .A2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n507), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(new_n517), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n536), .A2(new_n537), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n507), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n520), .A2(G43), .B1(new_n546), .B2(new_n517), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n513), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n507), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n513), .A2(G91), .B1(new_n558), .B2(G651), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n511), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n561), .A2(G53), .A3(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT74), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n510), .A2(new_n512), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  INV_X1    g140(.A(new_n562), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n561), .B1(new_n520), .B2(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n559), .B1(new_n568), .B2(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n533), .A2(KEYINPUT75), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n533), .A2(KEYINPUT75), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(G286));
  NAND2_X1  g149(.A1(new_n520), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n564), .A2(G87), .A3(new_n527), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G48), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT76), .B1(new_n564), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  AOI211_X1 g157(.A(new_n582), .B(new_n579), .C1(new_n510), .C2(new_n512), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n513), .A2(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n507), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(new_n517), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n513), .A2(G85), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n520), .A2(G47), .ZN(new_n594));
  INV_X1    g169(.A(new_n517), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n507), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n520), .A2(G54), .B1(new_n601), .B2(G651), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n513), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT10), .B1(new_n513), .B2(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g183(.A(KEYINPUT77), .B(new_n602), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G321));
  NOR2_X1   g187(.A1(G299), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G286), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  AOI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n617), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  OR3_X1    g196(.A1(new_n620), .A2(KEYINPUT78), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(KEYINPUT78), .B1(new_n620), .B2(new_n621), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n622), .B(new_n623), .C1(G868), .C2(new_n550), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n487), .A2(G135), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT79), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n481), .A2(G123), .ZN(new_n628));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT81), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n642), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT83), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n671), .A2(new_n672), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n670), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n670), .B2(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT84), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n687), .A2(new_n690), .A3(new_n688), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G6), .A2(G16), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n591), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n695), .A2(G23), .ZN(new_n704));
  NAND2_X1  g279(.A1(G288), .A2(KEYINPUT86), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT86), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n575), .A2(new_n576), .A3(new_n706), .A4(new_n577), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n704), .B1(new_n708), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT33), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT87), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n711), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n699), .A2(new_n703), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n481), .A2(G119), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(G107), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G2105), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n487), .B2(G131), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(new_n717), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT85), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  MUX2_X1   g305(.A(G24), .B(G290), .S(G16), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n716), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n734), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n695), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n695), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT95), .B(G1966), .Z(new_n742));
  XOR2_X1   g317(.A(new_n741), .B(new_n742), .Z(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  OR2_X1    g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n744), .A2(new_n717), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  NOR2_X1   g323(.A1(G5), .A2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT96), .Z(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G301), .B2(new_n695), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n747), .B1(new_n748), .B2(new_n751), .C1(new_n631), .C2(new_n717), .ZN(new_n752));
  OR3_X1    g327(.A1(new_n743), .A2(KEYINPUT97), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT97), .B1(new_n743), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n610), .A2(new_n695), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G4), .B2(new_n695), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT90), .B(G1348), .Z(new_n757));
  OAI211_X1 g332(.A(new_n753), .B(new_n754), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2090), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n717), .A2(G35), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n717), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(KEYINPUT29), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n762), .A2(new_n759), .A3(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n695), .A2(G19), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT91), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n549), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1341), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n764), .B(new_n770), .C1(new_n756), .C2(new_n757), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n717), .A2(G26), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT28), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n481), .A2(G128), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n775));
  INV_X1    g350(.A(G116), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G2105), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n487), .B2(G140), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT92), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G139), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n486), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n479), .A2(G127), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n461), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(G29), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G33), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(G29), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G2072), .Z(new_n795));
  INV_X1    g370(.A(G2078), .ZN(new_n796));
  NAND2_X1  g371(.A1(G164), .A2(G29), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G27), .B2(G29), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n796), .B2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n717), .A2(G32), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n481), .A2(G129), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n803));
  NAND3_X1  g378(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT26), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n803), .B(new_n805), .C1(new_n487), .C2(G141), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n801), .B1(new_n808), .B2(new_n717), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT94), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n751), .A2(new_n748), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n783), .A2(new_n800), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(G160), .A2(G29), .ZN(new_n815));
  INV_X1    g390(.A(G34), .ZN(new_n816));
  AOI21_X1  g391(.A(G29), .B1(new_n816), .B2(KEYINPUT24), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(KEYINPUT24), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G2084), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT93), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n695), .A2(G20), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT23), .Z(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G299), .B2(G16), .ZN(new_n825));
  INV_X1    g400(.A(G1956), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n820), .B2(new_n819), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n771), .A2(new_n814), .A3(new_n822), .A4(new_n828), .ZN(new_n829));
  NOR4_X1   g404(.A1(new_n737), .A2(new_n739), .A3(new_n758), .A4(new_n829), .ZN(G311));
  NOR3_X1   g405(.A1(new_n739), .A2(new_n758), .A3(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(new_n736), .ZN(G150));
  NAND2_X1  g407(.A1(new_n513), .A2(G93), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n520), .A2(G55), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n833), .B(new_n834), .C1(new_n595), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT99), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n610), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n549), .B(new_n836), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT98), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n843), .B2(new_n844), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n839), .B1(new_n846), .B2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(G160), .B(new_n489), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n631), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n481), .A2(G130), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n487), .A2(G142), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n461), .A2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n635), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n725), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT101), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n788), .A2(KEYINPUT100), .A3(new_n791), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G164), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n779), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(new_n807), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n807), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n858), .A2(KEYINPUT101), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n859), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n851), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n857), .B(new_n724), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT102), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n851), .B1(new_n873), .B2(new_n865), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n863), .A3(new_n864), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  OR2_X1    g454(.A1(G290), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(G290), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(new_n591), .ZN(new_n883));
  AOI21_X1  g458(.A(G305), .B1(new_n880), .B2(new_n881), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n708), .A2(G166), .ZN(new_n886));
  AOI21_X1  g461(.A(G303), .B1(new_n705), .B2(new_n707), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  OAI22_X1  g464(.A1(new_n883), .A2(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT42), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n889), .A2(KEYINPUT106), .A3(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n891), .B1(new_n896), .B2(KEYINPUT42), .ZN(new_n897));
  INV_X1    g472(.A(new_n606), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(KEYINPUT103), .A3(G299), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n513), .A2(G91), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n558), .A2(G651), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n904));
  AOI211_X1 g479(.A(KEYINPUT74), .B(new_n562), .C1(new_n510), .C2(new_n512), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n520), .A2(G53), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT9), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n900), .B1(new_n909), .B2(new_n606), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n899), .A2(new_n910), .B1(new_n909), .B2(new_n606), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n899), .A2(new_n910), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n899), .A2(KEYINPUT104), .A3(new_n910), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n909), .A2(new_n606), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n912), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n619), .B(new_n842), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n918), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n924), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n897), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n897), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(G868), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n836), .A2(new_n621), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(G295));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n932), .ZN(G331));
  XOR2_X1   g509(.A(new_n549), .B(new_n836), .Z(new_n935));
  OAI21_X1  g510(.A(G171), .B1(new_n572), .B2(new_n573), .ZN(new_n936));
  NOR2_X1   g511(.A1(G168), .A2(G171), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT75), .ZN(new_n942));
  NAND2_X1  g517(.A1(G168), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G301), .B1(new_n943), .B2(new_n571), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(new_n937), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(KEYINPUT109), .A3(new_n935), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n842), .B(new_n947), .C1(new_n944), .C2(new_n937), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n936), .A2(new_n938), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n947), .B1(new_n950), .B2(new_n842), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n941), .B(new_n946), .C1(new_n949), .C2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n842), .B1(new_n944), .B2(new_n937), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n939), .A2(new_n953), .A3(KEYINPUT110), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n945), .A2(new_n955), .A3(new_n935), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n920), .A2(new_n952), .B1(new_n918), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n889), .A2(KEYINPUT106), .A3(new_n890), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT106), .B1(new_n889), .B2(new_n890), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n918), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n954), .B(new_n956), .C1(new_n919), .C2(new_n911), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n952), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n919), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n896), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n962), .A2(new_n967), .A3(KEYINPUT43), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n920), .A2(new_n952), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n957), .A2(new_n918), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n896), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT43), .B1(new_n962), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n962), .A2(new_n967), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n962), .B2(new_n971), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(G397));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n464), .A2(KEYINPUT67), .A3(new_n465), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT67), .B1(new_n464), .B2(new_n465), .ZN(new_n983));
  OAI211_X1 g558(.A(G40), .B(new_n476), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n779), .B(new_n782), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n989), .A2(new_n808), .ZN(new_n990));
  INV_X1    g565(.A(new_n985), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT126), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(KEYINPUT47), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n807), .B(new_n986), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n989), .A2(new_n996), .A3(new_n728), .A4(new_n725), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n774), .A2(new_n782), .A3(new_n778), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n991), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n989), .A2(new_n996), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n724), .B(new_n728), .Z(new_n1001));
  OR2_X1    g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n1003));
  OR3_X1    g578(.A1(new_n991), .A2(G1986), .A3(G290), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n1002), .A2(new_n985), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1004), .A2(new_n1003), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n999), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n994), .A2(new_n995), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT63), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT112), .B(G8), .Z(new_n1010));
  INV_X1    g585(.A(new_n984), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n501), .A2(new_n503), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n497), .A2(new_n498), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1384), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n981), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n698), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n984), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1014), .A2(new_n1021), .A3(new_n1015), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n759), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1010), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1025));
  AND3_X1   g600(.A1(G303), .A2(G8), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT113), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n584), .A2(new_n590), .A3(G1981), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n582), .B1(new_n560), .B2(new_n579), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n564), .A2(KEYINPUT76), .A3(new_n580), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n513), .A2(G86), .B1(new_n588), .B2(new_n517), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1034), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1032), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1010), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n1019), .B2(new_n984), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(G1981), .B1(new_n584), .B2(new_n590), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1037), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n705), .A2(G1976), .A3(new_n707), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT52), .B1(new_n1048), .B2(new_n1042), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n705), .A2(G1976), .A3(new_n707), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1043), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1047), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(new_n1026), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1058), .A2(new_n1022), .A3(new_n1011), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1059), .A2(new_n759), .B1(new_n1017), .B2(new_n698), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1055), .B(new_n1057), .C1(new_n1060), .C2(new_n1010), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1030), .A2(new_n1062), .A3(G8), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1031), .A2(new_n1054), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1017), .A2(new_n1065), .A3(new_n742), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1020), .A2(new_n820), .A3(new_n1022), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1017), .B2(new_n742), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n614), .B(new_n1041), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1009), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1062), .A2(G8), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1009), .B1(new_n1072), .B2(new_n1057), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(new_n1063), .A3(new_n1054), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1047), .ZN(new_n1076));
  OR2_X1    g651(.A1(G288), .A2(G1976), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1045), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1063), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1078), .A2(new_n1043), .B1(new_n1079), .B2(new_n1054), .ZN(new_n1080));
  OAI21_X1  g655(.A(G8), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n533), .A2(new_n1041), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1082), .B(KEYINPUT121), .Z(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n533), .B(new_n1041), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(KEYINPUT51), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1041), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n1082), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(KEYINPUT62), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n981), .A2(new_n1011), .A3(new_n1016), .A4(new_n796), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1058), .A2(new_n1022), .A3(new_n1011), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n748), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1092), .A2(G2078), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1017), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(G171), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1064), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1090), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT62), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1075), .B(new_n1080), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n981), .A2(new_n1011), .A3(new_n1016), .A4(new_n986), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT118), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n984), .A2(G1996), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1107), .A2(new_n981), .A3(new_n1108), .A4(new_n1016), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT58), .B(G1341), .Z(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1019), .B2(new_n984), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1106), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n550), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT59), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1115), .A3(new_n550), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n909), .B2(KEYINPUT57), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n1119));
  NAND3_X1  g694(.A1(G299), .A2(KEYINPUT115), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT57), .B(new_n559), .C1(new_n568), .C2(new_n569), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n906), .A2(new_n908), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n559), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1017), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1129), .A2(new_n1130), .B1(new_n1094), .B2(new_n826), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1118), .A2(new_n1120), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n981), .A2(new_n1011), .A3(new_n1016), .A4(new_n1130), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1059), .B2(G1956), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1114), .A2(new_n1116), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n610), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1019), .A2(new_n984), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1094), .A2(new_n757), .B1(new_n782), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n610), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(KEYINPUT119), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(KEYINPUT119), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n1142), .A4(new_n1140), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1142), .A2(KEYINPUT60), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1128), .A2(new_n1150), .A3(new_n1131), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT117), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1151), .A2(new_n1152), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1138), .B(new_n1149), .C1(KEYINPUT61), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1128), .A2(new_n1131), .B1(new_n1144), .B2(new_n1142), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT120), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1092), .A2(new_n1091), .B1(new_n1094), .B2(new_n748), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1159), .B(G301), .C1(new_n1017), .C2(new_n1098), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n981), .A2(new_n1016), .A3(new_n1097), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n984), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n470), .A2(KEYINPUT122), .A3(G40), .A4(new_n476), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n981), .A2(new_n1016), .A3(new_n1097), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(KEYINPUT123), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1096), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(KEYINPUT54), .B(new_n1160), .C1(new_n1171), .C2(G301), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT125), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT54), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1170), .A2(new_n1167), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1159), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1174), .B1(new_n1176), .B2(G171), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1178), .A3(new_n1160), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1175), .A2(new_n1182), .A3(G301), .A4(new_n1159), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1183), .A2(new_n1174), .ZN(new_n1184));
  OAI211_X1 g759(.A(KEYINPUT124), .B(new_n1100), .C1(new_n1176), .C2(G171), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1064), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1180), .A2(new_n1181), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1158), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1154), .A2(KEYINPUT120), .A3(new_n1157), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1104), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1002), .ZN(new_n1191));
  XOR2_X1   g766(.A(G290), .B(G1986), .Z(new_n1192));
  AOI21_X1  g767(.A(new_n991), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1008), .B1(new_n1190), .B2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g769(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n692), .B2(new_n693), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n877), .B(new_n1197), .C1(new_n976), .C2(new_n977), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


