

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U324 ( .A(n375), .B(n332), .ZN(n333) );
  XNOR2_X1 U325 ( .A(n396), .B(n333), .ZN(n334) );
  XNOR2_X1 U326 ( .A(n340), .B(n339), .ZN(n341) );
  NOR2_X1 U327 ( .A1(n430), .A2(n519), .ZN(n456) );
  XNOR2_X1 U328 ( .A(n342), .B(n341), .ZN(n345) );
  NOR2_X1 U329 ( .A1(n533), .A2(n450), .ZN(n572) );
  XNOR2_X1 U330 ( .A(n451), .B(G190GAT), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(G120GAT), .B(G71GAT), .Z(n343) );
  XOR2_X1 U333 ( .A(G15GAT), .B(G127GAT), .Z(n361) );
  XNOR2_X1 U334 ( .A(n343), .B(n361), .ZN(n294) );
  XOR2_X1 U335 ( .A(KEYINPUT0), .B(KEYINPUT85), .Z(n293) );
  XNOR2_X1 U336 ( .A(G113GAT), .B(G134GAT), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n427) );
  XNOR2_X1 U338 ( .A(n294), .B(n427), .ZN(n300) );
  XOR2_X1 U339 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n296) );
  XNOR2_X1 U340 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n405) );
  XOR2_X1 U342 ( .A(G176GAT), .B(n405), .Z(n298) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U345 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(G99GAT), .Z(n302) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U349 ( .A(G183GAT), .B(KEYINPUT86), .Z(n304) );
  XNOR2_X1 U350 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n533) );
  INV_X1 U354 ( .A(KEYINPUT54), .ZN(n409) );
  XOR2_X1 U355 ( .A(G197GAT), .B(G22GAT), .Z(n310) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(G141GAT), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U358 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n312) );
  XNOR2_X1 U359 ( .A(G8GAT), .B(KEYINPUT70), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U361 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT68), .B(KEYINPUT74), .Z(n316) );
  NAND2_X1 U363 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U365 ( .A(KEYINPUT30), .B(n317), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U367 ( .A(G36GAT), .B(G50GAT), .Z(n322) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(KEYINPUT72), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n320), .B(KEYINPUT73), .ZN(n357) );
  XNOR2_X1 U370 ( .A(G15GAT), .B(n357), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U372 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U373 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n326) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(G29GAT), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U376 ( .A(KEYINPUT71), .B(n327), .Z(n374) );
  XNOR2_X1 U377 ( .A(G169GAT), .B(n374), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n575) );
  XOR2_X1 U379 ( .A(G64GAT), .B(G92GAT), .Z(n331) );
  XNOR2_X1 U380 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n396) );
  XOR2_X1 U382 ( .A(G99GAT), .B(G85GAT), .Z(n375) );
  AND2_X1 U383 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XOR2_X1 U384 ( .A(n334), .B(KEYINPUT31), .Z(n342) );
  XOR2_X1 U385 ( .A(G78GAT), .B(G148GAT), .Z(n336) );
  XNOR2_X1 U386 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n431) );
  XNOR2_X1 U388 ( .A(n431), .B(KEYINPUT32), .ZN(n340) );
  XOR2_X1 U389 ( .A(KEYINPUT78), .B(KEYINPUT76), .Z(n338) );
  XNOR2_X1 U390 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n337) );
  XOR2_X1 U391 ( .A(n338), .B(n337), .Z(n339) );
  XOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT13), .Z(n360) );
  XNOR2_X1 U393 ( .A(n343), .B(n360), .ZN(n344) );
  XNOR2_X1 U394 ( .A(n345), .B(n344), .ZN(n389) );
  XNOR2_X1 U395 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n346) );
  XOR2_X1 U396 ( .A(n389), .B(n346), .Z(n556) );
  INV_X1 U397 ( .A(n556), .ZN(n567) );
  NAND2_X1 U398 ( .A1(n575), .A2(n567), .ZN(n348) );
  INV_X1 U399 ( .A(KEYINPUT46), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n370) );
  XOR2_X1 U401 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n350) );
  XNOR2_X1 U402 ( .A(KEYINPUT80), .B(KEYINPUT82), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n369) );
  XOR2_X1 U404 ( .A(G64GAT), .B(G78GAT), .Z(n352) );
  XNOR2_X1 U405 ( .A(G71GAT), .B(G211GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U407 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n354) );
  XNOR2_X1 U408 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U410 ( .A(n356), .B(n355), .Z(n367) );
  XOR2_X1 U411 ( .A(n357), .B(KEYINPUT84), .Z(n359) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n365) );
  XOR2_X1 U414 ( .A(G8GAT), .B(G183GAT), .Z(n400) );
  XOR2_X1 U415 ( .A(n360), .B(n400), .Z(n363) );
  XOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .Z(n438) );
  XNOR2_X1 U417 ( .A(n361), .B(n438), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U421 ( .A(n369), .B(n368), .Z(n579) );
  NOR2_X1 U422 ( .A1(n370), .A2(n579), .ZN(n386) );
  XOR2_X1 U423 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n372) );
  XNOR2_X1 U424 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n385) );
  XOR2_X1 U427 ( .A(G36GAT), .B(G190GAT), .Z(n397) );
  XOR2_X1 U428 ( .A(n375), .B(n397), .Z(n377) );
  XNOR2_X1 U429 ( .A(G218GAT), .B(G92GAT), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U431 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n379) );
  NAND2_X1 U432 ( .A1(G232GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U434 ( .A(n381), .B(n380), .Z(n383) );
  XOR2_X1 U435 ( .A(G50GAT), .B(G162GAT), .Z(n432) );
  XNOR2_X1 U436 ( .A(n432), .B(G106GAT), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n563) );
  NAND2_X1 U439 ( .A1(n386), .A2(n563), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n387), .B(KEYINPUT47), .ZN(n394) );
  XNOR2_X1 U441 ( .A(n563), .B(KEYINPUT36), .ZN(n582) );
  INV_X1 U442 ( .A(n579), .ZN(n559) );
  NOR2_X1 U443 ( .A1(n582), .A2(n559), .ZN(n388) );
  XNOR2_X1 U444 ( .A(KEYINPUT45), .B(n388), .ZN(n390) );
  NAND2_X1 U445 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U446 ( .A(KEYINPUT116), .B(n391), .ZN(n392) );
  NOR2_X1 U447 ( .A1(n392), .A2(n575), .ZN(n393) );
  NOR2_X1 U448 ( .A1(n394), .A2(n393), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n395), .B(KEYINPUT48), .ZN(n549) );
  XOR2_X1 U450 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U451 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U453 ( .A(n401), .B(n400), .Z(n407) );
  XOR2_X1 U454 ( .A(KEYINPUT91), .B(G218GAT), .Z(n403) );
  XNOR2_X1 U455 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n402) );
  XNOR2_X1 U456 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U457 ( .A(G197GAT), .B(n404), .ZN(n447) );
  XOR2_X1 U458 ( .A(n405), .B(n447), .Z(n406) );
  XNOR2_X1 U459 ( .A(n407), .B(n406), .ZN(n465) );
  NOR2_X1 U460 ( .A1(n549), .A2(n465), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n409), .B(n408), .ZN(n430) );
  XOR2_X1 U462 ( .A(G85GAT), .B(G162GAT), .Z(n411) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(G120GAT), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U465 ( .A(G155GAT), .B(G148GAT), .Z(n413) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(G127GAT), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U468 ( .A(n415), .B(n414), .Z(n420) );
  XOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n417) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U472 ( .A(KEYINPUT6), .B(n418), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U474 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n422) );
  XNOR2_X1 U475 ( .A(KEYINPUT96), .B(G57GAT), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U477 ( .A(n424), .B(n423), .Z(n429) );
  XOR2_X1 U478 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n426) );
  XNOR2_X1 U479 ( .A(G141GAT), .B(KEYINPUT92), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n442) );
  XNOR2_X1 U481 ( .A(n427), .B(n442), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n519) );
  XOR2_X1 U483 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n446) );
  XOR2_X1 U486 ( .A(G204GAT), .B(KEYINPUT90), .Z(n436) );
  XNOR2_X1 U487 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U489 ( .A(n437), .B(KEYINPUT94), .Z(n440) );
  XNOR2_X1 U490 ( .A(n438), .B(KEYINPUT89), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U492 ( .A(n441), .B(KEYINPUT22), .Z(n444) );
  XNOR2_X1 U493 ( .A(n442), .B(KEYINPUT93), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U495 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U496 ( .A(n448), .B(n447), .ZN(n467) );
  NAND2_X1 U497 ( .A1(n456), .A2(n467), .ZN(n449) );
  XOR2_X1 U498 ( .A(KEYINPUT55), .B(n449), .Z(n450) );
  INV_X1 U499 ( .A(n563), .ZN(n543) );
  NAND2_X1 U500 ( .A1(n572), .A2(n543), .ZN(n453) );
  XOR2_X1 U501 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n451) );
  INV_X1 U502 ( .A(G204GAT), .ZN(n461) );
  XOR2_X1 U503 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n459) );
  INV_X1 U504 ( .A(n533), .ZN(n526) );
  NOR2_X1 U505 ( .A1(n526), .A2(n467), .ZN(n455) );
  XNOR2_X1 U506 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n551) );
  NAND2_X1 U508 ( .A1(n456), .A2(n551), .ZN(n457) );
  XOR2_X1 U509 ( .A(KEYINPUT126), .B(n457), .Z(n580) );
  INV_X1 U510 ( .A(n580), .ZN(n583) );
  OR2_X1 U511 ( .A1(n583), .A2(n389), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n461), .B(n460), .ZN(G1353GAT) );
  NAND2_X1 U514 ( .A1(n575), .A2(n389), .ZN(n492) );
  NOR2_X1 U515 ( .A1(n543), .A2(n559), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n462), .B(KEYINPUT16), .ZN(n476) );
  XOR2_X1 U517 ( .A(n465), .B(KEYINPUT27), .Z(n469) );
  NAND2_X1 U518 ( .A1(n519), .A2(n469), .ZN(n548) );
  XNOR2_X1 U519 ( .A(KEYINPUT67), .B(KEYINPUT28), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(n467), .ZN(n528) );
  NOR2_X1 U521 ( .A1(n548), .A2(n528), .ZN(n535) );
  NAND2_X1 U522 ( .A1(n533), .A2(n535), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT97), .B(n464), .Z(n475) );
  INV_X1 U524 ( .A(n519), .ZN(n473) );
  INV_X1 U525 ( .A(n465), .ZN(n523) );
  NAND2_X1 U526 ( .A1(n526), .A2(n523), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(n468), .Z(n471) );
  NAND2_X1 U529 ( .A1(n551), .A2(n469), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n488) );
  NAND2_X1 U533 ( .A1(n476), .A2(n488), .ZN(n505) );
  NOR2_X1 U534 ( .A1(n492), .A2(n505), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT99), .B(n477), .Z(n485) );
  NAND2_X1 U536 ( .A1(n485), .A2(n519), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n523), .A2(n485), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT100), .ZN(n481) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(n481), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U543 ( .A1(n485), .A2(n526), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U545 ( .A(G15GAT), .B(n484), .Z(G1326GAT) );
  NAND2_X1 U546 ( .A1(n528), .A2(n485), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U548 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n487), .B(KEYINPUT38), .ZN(n494) );
  NAND2_X1 U550 ( .A1(n559), .A2(n488), .ZN(n489) );
  NOR2_X1 U551 ( .A1(n582), .A2(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n517) );
  NOR2_X1 U554 ( .A1(n492), .A2(n517), .ZN(n493) );
  XOR2_X1 U555 ( .A(n494), .B(n493), .Z(n502) );
  NAND2_X1 U556 ( .A1(n519), .A2(n502), .ZN(n496) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT105), .Z(n498) );
  NAND2_X1 U560 ( .A1(n502), .A2(n523), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n500) );
  NAND2_X1 U563 ( .A1(n502), .A2(n526), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U565 ( .A(G43GAT), .B(n501), .Z(G1330GAT) );
  XOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT107), .Z(n504) );
  NAND2_X1 U567 ( .A1(n502), .A2(n528), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  INV_X1 U570 ( .A(n575), .ZN(n552) );
  NAND2_X1 U571 ( .A1(n567), .A2(n552), .ZN(n516) );
  NOR2_X1 U572 ( .A1(n505), .A2(n516), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n506), .B(KEYINPUT108), .ZN(n512) );
  NAND2_X1 U574 ( .A1(n519), .A2(n512), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  XOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT109), .Z(n510) );
  NAND2_X1 U577 ( .A1(n512), .A2(n523), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n512), .A2(n526), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U582 ( .A1(n512), .A2(n528), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n521) );
  NOR2_X1 U586 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U587 ( .A(KEYINPUT111), .B(n518), .Z(n529) );
  NAND2_X1 U588 ( .A1(n529), .A2(n519), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n523), .A2(n529), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n524), .B(KEYINPUT114), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n525), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n526), .A2(n529), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT44), .Z(n531) );
  NAND2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U600 ( .A1(n549), .A2(n533), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT117), .B(n536), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n575), .A2(n544), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n539) );
  NAND2_X1 U606 ( .A1(n544), .A2(n567), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n544), .A2(n579), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n562) );
  NOR2_X1 U618 ( .A1(n552), .A2(n562), .ZN(n553) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n556), .A2(n562), .ZN(n557) );
  XOR2_X1 U624 ( .A(n558), .B(n557), .Z(G1345GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n562), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n575), .A2(n572), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n569) );
  NAND2_X1 U634 ( .A1(n572), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT56), .Z(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n579), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(n574), .ZN(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  NAND2_X1 U642 ( .A1(n575), .A2(n580), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

