//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n558, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT69), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(KEYINPUT3), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n465), .A2(new_n470), .A3(G137), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n463), .A2(G2104), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT67), .Z(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n472), .A2(new_n485), .A3(new_n474), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n476), .A2(new_n484), .A3(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n465), .A2(new_n470), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n488), .A2(new_n471), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  AND2_X1   g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n465), .A2(new_n470), .A3(new_n471), .A4(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n465), .A2(new_n470), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n477), .A2(new_n478), .A3(G138), .A4(new_n471), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n498), .A2(new_n500), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT71), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  INV_X1    g090(.A(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n517), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT72), .A3(G543), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(new_n520), .B1(KEYINPUT5), .B2(new_n512), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n514), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n508), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n523), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  XOR2_X1   g103(.A(KEYINPUT73), .B(G51), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n513), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n521), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n511), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n521), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n530), .A2(new_n533), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n513), .A2(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n542), .B2(new_n522), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n525), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n543), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  AOI22_X1  g122(.A1(G43), .A2(new_n513), .B1(new_n532), .B2(G81), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n525), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT74), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(KEYINPUT74), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT75), .Z(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT76), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n513), .A2(G53), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(KEYINPUT77), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n562), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n531), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n532), .A2(G91), .B1(G651), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n532), .A2(G87), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT78), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT79), .Z(new_n574));
  NAND2_X1  g149(.A1(new_n513), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(G288));
  OAI211_X1 g151(.A(G86), .B(new_n521), .C1(new_n509), .C2(new_n510), .ZN(new_n577));
  OAI211_X1 g152(.A(G48), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n521), .A2(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT80), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n577), .B(new_n578), .C1(new_n582), .C2(new_n525), .ZN(G305));
  AOI22_X1  g158(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n525), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n522), .A2(new_n586), .ZN(new_n587));
  AOI211_X1 g162(.A(new_n585), .B(new_n587), .C1(G47), .C2(new_n513), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT81), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n532), .A2(G92), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT10), .Z(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n531), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n513), .A2(G54), .B1(G651), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n590), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n590), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G299), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  NOR2_X1   g181(.A1(new_n597), .A2(G559), .ZN(new_n607));
  OR3_X1    g182(.A1(new_n607), .A2(KEYINPUT82), .A3(new_n601), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT82), .B1(new_n607), .B2(new_n601), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n608), .B(new_n609), .C1(G868), .C2(new_n554), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n468), .A2(new_n469), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n479), .A2(new_n612), .A3(new_n471), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n489), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n491), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n471), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n616), .A2(new_n623), .ZN(G156));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n628), .B(new_n634), .Z(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n638), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(G401));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2096), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n645), .B2(KEYINPUT18), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT86), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(G227));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT87), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n656), .A2(new_n658), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n661), .A3(new_n659), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n666), .C1(new_n661), .C2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G288), .ZN(new_n674));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n675), .B2(G23), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT33), .B(G1976), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(G22), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n675), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(G1971), .Z(new_n683));
  MUX2_X1   g258(.A(G6), .B(G305), .S(G16), .Z(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n679), .A2(new_n680), .A3(new_n683), .A4(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(KEYINPUT34), .ZN(new_n688));
  NAND2_X1  g263(.A1(G290), .A2(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n675), .A2(G24), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT88), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(KEYINPUT88), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G1986), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n489), .A2(G131), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n491), .A2(G119), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n696), .B1(new_n702), .B2(new_n695), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  AND2_X1   g280(.A1(new_n693), .A2(G1986), .ZN(new_n706));
  NOR4_X1   g281(.A1(new_n688), .A2(new_n694), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n687), .A2(KEYINPUT34), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT89), .B(KEYINPUT36), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n712));
  OAI211_X1 g287(.A(KEYINPUT90), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n710), .A2(KEYINPUT90), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n675), .A2(G21), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G168), .B2(new_n675), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT95), .Z(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(G1966), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(G1966), .ZN(new_n719));
  NAND2_X1  g294(.A1(G301), .A2(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n675), .A2(G5), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT30), .B(G28), .ZN(new_n725));
  OR2_X1    g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n725), .A2(new_n695), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n621), .B2(new_n695), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT96), .ZN(new_n730));
  NOR4_X1   g305(.A1(new_n718), .A2(new_n719), .A3(new_n724), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT97), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G160), .B2(new_n695), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT91), .Z(new_n738));
  INV_X1    g313(.A(G2084), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n489), .A2(G141), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n491), .A2(G129), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT26), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI22_X1  g321(.A1(G105), .A2(new_n473), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n741), .A2(new_n742), .A3(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G32), .B(new_n748), .S(G29), .Z(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2072), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n695), .A2(G33), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n489), .A2(G139), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT25), .Z(new_n757));
  AOI22_X1  g332(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n757), .C1(new_n471), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n754), .B1(new_n759), .B2(G29), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n722), .A2(new_n723), .B1(new_n753), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n695), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n695), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n760), .A2(new_n753), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT92), .ZN(new_n767));
  AND4_X1   g342(.A1(new_n752), .A2(new_n761), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n738), .A2(new_n739), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n749), .A2(new_n751), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT94), .Z(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n732), .A2(new_n740), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G4), .A2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n598), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1348), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n695), .A2(G26), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT28), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n489), .A2(G140), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n491), .A2(G128), .ZN(new_n782));
  OR2_X1    g357(.A1(G104), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(new_n695), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n778), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n554), .A2(new_n675), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n675), .B2(G19), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G1341), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n695), .A2(G35), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G162), .B2(new_n695), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT29), .Z(new_n796));
  INV_X1    g371(.A(G2090), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n792), .B2(G1341), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n675), .A2(G20), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT23), .Z(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n797), .B2(new_n796), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n789), .A2(new_n793), .A3(new_n799), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n773), .B2(new_n774), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n713), .A2(new_n714), .A3(new_n775), .A4(new_n807), .ZN(G150));
  INV_X1    g383(.A(G150), .ZN(G311));
  NAND2_X1  g384(.A1(new_n521), .A2(G67), .ZN(new_n810));
  NAND2_X1  g385(.A1(G80), .A2(G543), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n525), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n513), .A2(G55), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n532), .A2(G93), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n554), .B2(KEYINPUT100), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n554), .A2(KEYINPUT100), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT38), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n598), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n824), .A2(new_n825), .A3(G860), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n817), .A2(G860), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  NAND2_X1  g404(.A1(new_n491), .A2(G130), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n471), .A2(G118), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G142), .B2(new_n489), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(new_n614), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n759), .B(new_n748), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n500), .A2(new_n502), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n498), .A2(new_n505), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n500), .A2(KEYINPUT101), .A3(new_n502), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n785), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n702), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n837), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G160), .B(new_n621), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n495), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT102), .Z(new_n850));
  AOI21_X1  g425(.A(G37), .B1(new_n846), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(G395));
  NAND2_X1  g429(.A1(new_n817), .A2(new_n601), .ZN(new_n855));
  XNOR2_X1  g430(.A(G290), .B(G303), .ZN(new_n856));
  XNOR2_X1  g431(.A(G288), .B(G305), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n856), .B(new_n857), .Z(new_n858));
  XOR2_X1   g433(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n820), .B(new_n607), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n597), .B(G299), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT41), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n862), .B2(new_n861), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n860), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n855), .B1(new_n866), .B2(new_n601), .ZN(G295));
  OAI21_X1  g442(.A(new_n855), .B1(new_n866), .B2(new_n601), .ZN(G331));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n869));
  XNOR2_X1  g444(.A(G301), .B(G286), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n820), .B(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n862), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n871), .A2(new_n863), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(KEYINPUT105), .ZN(new_n874));
  INV_X1    g449(.A(new_n858), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n874), .B(new_n875), .C1(KEYINPUT105), .C2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n858), .B1(new_n873), .B2(new_n872), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT43), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(KEYINPUT105), .ZN(new_n882));
  INV_X1    g457(.A(new_n872), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n873), .A2(KEYINPUT105), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n858), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n876), .A4(new_n878), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n869), .B1(new_n881), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n878), .A3(new_n876), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n876), .A2(new_n887), .ZN(new_n891));
  AOI22_X1  g466(.A1(KEYINPUT43), .A2(new_n890), .B1(new_n891), .B2(new_n879), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n869), .B2(new_n892), .ZN(G397));
  INV_X1    g468(.A(G1384), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n843), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(KEYINPUT45), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n476), .A2(G40), .A3(new_n484), .A4(new_n486), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT106), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n898), .A2(KEYINPUT107), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT107), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n903), .A2(G1986), .A3(G290), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT48), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(new_n903), .ZN(new_n908));
  INV_X1    g483(.A(G2067), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n785), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G1996), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n748), .B(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n702), .A2(new_n704), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n702), .A2(new_n704), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n910), .A2(new_n912), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  AOI211_X1 g490(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n910), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n908), .B1(new_n748), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(new_n908), .B2(new_n911), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n903), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT47), .Z(new_n923));
  NAND2_X1  g498(.A1(new_n910), .A2(new_n912), .ZN(new_n924));
  OAI22_X1  g499(.A1(new_n924), .A2(new_n914), .B1(G2067), .B2(new_n785), .ZN(new_n925));
  AOI211_X1 g500(.A(new_n916), .B(new_n923), .C1(new_n908), .C2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G290), .B(G1986), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n908), .B1(new_n927), .B2(new_n915), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT108), .Z(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n500), .A2(KEYINPUT101), .A3(new_n502), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT101), .B1(new_n500), .B2(new_n502), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n498), .A2(new_n505), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n930), .B1(new_n934), .B2(G1384), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n843), .A2(KEYINPUT109), .A3(new_n894), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  NOR2_X1   g514(.A1(G164), .A2(G1384), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(new_n936), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(G160), .A2(KEYINPUT106), .A3(G40), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n899), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n935), .A2(new_n939), .A3(new_n936), .A4(new_n937), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT120), .ZN(new_n949));
  INV_X1    g524(.A(G1348), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT120), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n942), .A2(new_n951), .A3(new_n946), .A4(new_n947), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n935), .A2(new_n937), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n900), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n909), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(KEYINPUT60), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT122), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT122), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n953), .A2(new_n959), .A3(KEYINPUT60), .A4(new_n956), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n953), .A2(new_n956), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT60), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n598), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  MUX2_X1   g541(.A(new_n940), .B(new_n895), .S(KEYINPUT45), .Z(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT56), .B(G2072), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n967), .A2(new_n946), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n943), .A2(new_n945), .B1(new_n936), .B2(new_n940), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n803), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n974), .A3(KEYINPUT121), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT121), .ZN(new_n976));
  AOI21_X1  g551(.A(G1956), .B1(new_n971), .B2(new_n972), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(new_n969), .ZN(new_n978));
  NAND2_X1  g553(.A1(G299), .A2(KEYINPUT57), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n565), .A2(new_n980), .A3(new_n569), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n975), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n982), .A2(new_n977), .A3(new_n969), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(KEYINPUT61), .A3(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT58), .B(G1341), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n955), .A2(new_n987), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n967), .A2(new_n911), .A3(new_n946), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n554), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT59), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT61), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n970), .A2(new_n974), .B1(new_n979), .B2(new_n981), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(new_n984), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n986), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n958), .A2(new_n964), .A3(new_n598), .A4(new_n960), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n966), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n962), .A2(new_n598), .A3(new_n985), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n998), .A2(new_n983), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT124), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT123), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n940), .A2(KEYINPUT45), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT117), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n954), .A2(new_n1005), .B1(new_n943), .B2(new_n945), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n935), .B2(new_n937), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT116), .B1(new_n1009), .B2(new_n900), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1966), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n948), .A2(G2084), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1002), .B(G8), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G168), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(KEYINPUT51), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n843), .A2(KEYINPUT109), .A3(new_n894), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT109), .B1(new_n843), .B2(new_n894), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1005), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(new_n1007), .A3(new_n946), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1003), .B(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1010), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1966), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n942), .A2(new_n946), .A3(new_n947), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n739), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1002), .B1(new_n1029), .B2(G8), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1001), .B1(new_n1017), .B2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1025), .A2(new_n1024), .B1(new_n1027), .B2(new_n739), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT123), .B1(new_n1032), .B2(new_n1014), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1033), .A2(new_n1013), .A3(KEYINPUT124), .A4(new_n1016), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1015), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT51), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1031), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n949), .A2(new_n723), .A3(new_n952), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n967), .A2(new_n946), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n764), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(G301), .B(KEYINPUT54), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n764), .A2(KEYINPUT53), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n896), .B2(KEYINPUT45), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n471), .B1(new_n483), .B2(KEYINPUT125), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(KEYINPUT125), .B2(new_n483), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1053), .A2(G40), .A3(new_n476), .A4(new_n486), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1054), .A2(KEYINPUT126), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(KEYINPUT126), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n897), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1049), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1024), .A2(new_n1050), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1048), .A2(new_n1058), .B1(new_n1060), .B2(new_n1049), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G305), .A2(G1981), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT49), .B1(new_n1062), .B2(KEYINPUT112), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1064), .B(new_n1065), .C1(G305), .C2(G1981), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(G1981), .A3(G305), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G305), .A2(G1981), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n899), .A2(new_n944), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n899), .A2(new_n944), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n935), .B(new_n937), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1073), .A2(KEYINPUT111), .A3(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT111), .B1(new_n1073), .B2(G8), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1068), .B(new_n1070), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n674), .A2(G1976), .ZN(new_n1077));
  INV_X1    g652(.A(G1976), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT52), .B1(G288), .B2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1077), .B(new_n1079), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n955), .B2(new_n1014), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1073), .A2(KEYINPUT111), .A3(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1086), .B2(new_n1077), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT115), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1077), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT52), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(new_n1080), .A4(new_n1076), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n948), .A2(G2090), .B1(new_n1044), .B2(G1971), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G303), .A2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1097), .A3(G8), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n971), .A2(new_n972), .A3(new_n797), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1971), .B1(new_n967), .B2(new_n946), .ZN(new_n1100));
  OAI21_X1  g675(.A(G8), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1095), .B(KEYINPUT55), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1061), .A2(new_n1093), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1000), .A2(new_n1042), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1029), .A2(G8), .A3(G168), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1104), .B(new_n1110), .C1(new_n1088), .C2(new_n1092), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1109), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1093), .A2(new_n1105), .ZN(new_n1115));
  OAI211_X1 g690(.A(KEYINPUT119), .B(new_n1112), .C1(new_n1115), .C2(new_n1110), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1090), .A2(new_n1080), .A3(new_n1076), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n1110), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1094), .A2(G8), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1102), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1118), .A2(KEYINPUT63), .A3(new_n1098), .A4(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1114), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G288), .A2(G1976), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT114), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1062), .B1(new_n1124), .B2(new_n1076), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1086), .B(KEYINPUT113), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1125), .A2(new_n1126), .B1(new_n1117), .B2(new_n1098), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1108), .A2(new_n1122), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(G301), .B1(new_n1048), .B2(new_n1059), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1093), .A2(new_n1105), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1042), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1039), .A2(KEYINPUT62), .A3(new_n1041), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(KEYINPUT127), .B(new_n929), .C1(new_n1129), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1131), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1033), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1139), .A2(new_n1001), .B1(new_n1037), .B2(KEYINPUT51), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1132), .B(new_n1040), .C1(new_n1140), .C2(new_n1034), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT62), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1138), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1106), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1127), .B1(new_n1144), .B2(new_n1000), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1122), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT127), .B1(new_n1146), .B2(new_n929), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n926), .B1(new_n1137), .B2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g723(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n852), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g725(.A1(new_n892), .A2(new_n1151), .ZN(G308));
  OR2_X1    g726(.A1(new_n892), .A2(new_n1151), .ZN(G225));
endmodule


