

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G2104), .A2(n580), .ZN(n884) );
  INV_X1 U551 ( .A(n730), .ZN(n747) );
  NOR2_X2 U552 ( .A1(G2105), .A2(n575), .ZN(n902) );
  NOR2_X1 U553 ( .A1(n737), .A2(n736), .ZN(n515) );
  INV_X1 U554 ( .A(KEYINPUT26), .ZN(n662) );
  XNOR2_X1 U555 ( .A(n693), .B(KEYINPUT96), .ZN(n694) );
  XNOR2_X1 U556 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U557 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U558 ( .A(n726), .B(KEYINPUT100), .ZN(n735) );
  INV_X1 U559 ( .A(n745), .ZN(n746) );
  NAND2_X1 U560 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U561 ( .A(n748), .B(KEYINPUT104), .ZN(n749) );
  NOR2_X1 U562 ( .A1(G651), .A2(n568), .ZN(n806) );
  XOR2_X1 U563 ( .A(KEYINPUT17), .B(n579), .Z(n903) );
  XNOR2_X1 U564 ( .A(n761), .B(KEYINPUT106), .ZN(n762) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n568) );
  INV_X1 U566 ( .A(G651), .ZN(n516) );
  NOR2_X1 U567 ( .A1(n568), .A2(n516), .ZN(n809) );
  NAND2_X1 U568 ( .A1(G72), .A2(n809), .ZN(n519) );
  NOR2_X1 U569 ( .A1(G543), .A2(n516), .ZN(n517) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n517), .Z(n805) );
  NAND2_X1 U571 ( .A1(G60), .A2(n805), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n519), .A2(n518), .ZN(n523) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n520) );
  XNOR2_X1 U574 ( .A(n520), .B(KEYINPUT64), .ZN(n810) );
  NAND2_X1 U575 ( .A1(G85), .A2(n810), .ZN(n521) );
  XNOR2_X1 U576 ( .A(KEYINPUT65), .B(n521), .ZN(n522) );
  NOR2_X1 U577 ( .A1(n523), .A2(n522), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n806), .A2(G47), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n525), .A2(n524), .ZN(G290) );
  NAND2_X1 U580 ( .A1(n810), .A2(G86), .ZN(n532) );
  NAND2_X1 U581 ( .A1(G61), .A2(n805), .ZN(n527) );
  NAND2_X1 U582 ( .A1(G48), .A2(n806), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n530) );
  NAND2_X1 U584 ( .A1(G73), .A2(n809), .ZN(n528) );
  XOR2_X1 U585 ( .A(KEYINPUT2), .B(n528), .Z(n529) );
  NOR2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n533), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U589 ( .A1(G62), .A2(n805), .ZN(n535) );
  NAND2_X1 U590 ( .A1(G88), .A2(n810), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U592 ( .A1(G75), .A2(n809), .ZN(n537) );
  NAND2_X1 U593 ( .A1(G50), .A2(n806), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U596 ( .A(KEYINPUT79), .B(n540), .ZN(G303) );
  NAND2_X1 U597 ( .A1(G90), .A2(n810), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT67), .B(n541), .Z(n543) );
  NAND2_X1 U599 ( .A1(n809), .A2(G77), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n544), .B(KEYINPUT9), .ZN(n546) );
  NAND2_X1 U602 ( .A1(G64), .A2(n805), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n806), .A2(G52), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT66), .B(n547), .Z(n548) );
  NOR2_X1 U606 ( .A1(n549), .A2(n548), .ZN(G171) );
  NAND2_X1 U607 ( .A1(G65), .A2(n805), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G53), .A2(n806), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U610 ( .A(KEYINPUT69), .B(n552), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G78), .A2(n809), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G91), .A2(n810), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT68), .B(n555), .Z(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(G299) );
  NAND2_X1 U616 ( .A1(G89), .A2(n810), .ZN(n558) );
  XNOR2_X1 U617 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G76), .A2(n809), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U621 ( .A1(G63), .A2(n805), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G51), .A2(n806), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G49), .A2(n806), .ZN(n570) );
  NAND2_X1 U629 ( .A1(G87), .A2(n568), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U631 ( .A1(n805), .A2(n571), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G74), .A2(G651), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT77), .B(n572), .Z(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(G288) );
  INV_X1 U635 ( .A(G2104), .ZN(n575) );
  INV_X1 U636 ( .A(G2105), .ZN(n580) );
  NOR2_X1 U637 ( .A1(n575), .A2(n580), .ZN(n599) );
  NAND2_X1 U638 ( .A1(n599), .A2(G113), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G101), .A2(n902), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT23), .B(n576), .Z(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n584) );
  NOR2_X1 U642 ( .A1(G2104), .A2(G2105), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G137), .A2(n903), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G125), .A2(n884), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n584), .A2(n583), .ZN(G160) );
  NAND2_X1 U647 ( .A1(G160), .A2(G40), .ZN(n637) );
  INV_X1 U648 ( .A(G1384), .ZN(n590) );
  AND2_X1 U649 ( .A1(G138), .A2(n590), .ZN(n585) );
  AND2_X1 U650 ( .A1(n903), .A2(n585), .ZN(n592) );
  NAND2_X1 U651 ( .A1(G114), .A2(n599), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G126), .A2(n884), .ZN(n586) );
  AND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G102), .A2(n902), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n783) );
  AND2_X1 U656 ( .A1(n590), .A2(n783), .ZN(n591) );
  OR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n635) );
  NOR2_X1 U658 ( .A1(n637), .A2(n635), .ZN(n593) );
  XOR2_X1 U659 ( .A(n593), .B(KEYINPUT83), .Z(n753) );
  INV_X1 U660 ( .A(n753), .ZN(n634) );
  NAND2_X1 U661 ( .A1(n903), .A2(G140), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n902), .A2(G104), .ZN(n594) );
  XOR2_X1 U663 ( .A(KEYINPUT85), .B(n594), .Z(n595) );
  NAND2_X1 U664 ( .A1(n596), .A2(n595), .ZN(n598) );
  XOR2_X1 U665 ( .A(KEYINPUT34), .B(KEYINPUT86), .Z(n597) );
  XNOR2_X1 U666 ( .A(n598), .B(n597), .ZN(n605) );
  NAND2_X1 U667 ( .A1(G116), .A2(n599), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G128), .A2(n884), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n603) );
  XOR2_X1 U670 ( .A(KEYINPUT35), .B(KEYINPUT87), .Z(n602) );
  XNOR2_X1 U671 ( .A(n603), .B(n602), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U673 ( .A(KEYINPUT36), .B(n606), .ZN(n914) );
  XOR2_X1 U674 ( .A(G2067), .B(KEYINPUT37), .Z(n607) );
  NOR2_X1 U675 ( .A1(n914), .A2(n607), .ZN(n958) );
  AND2_X1 U676 ( .A1(n914), .A2(n607), .ZN(n959) );
  NAND2_X1 U677 ( .A1(G117), .A2(n599), .ZN(n609) );
  NAND2_X1 U678 ( .A1(G129), .A2(n884), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n902), .A2(G105), .ZN(n610) );
  XOR2_X1 U681 ( .A(KEYINPUT38), .B(n610), .Z(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT89), .B(n613), .Z(n615) );
  NAND2_X1 U684 ( .A1(n903), .A2(G141), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n909) );
  NOR2_X1 U686 ( .A1(G1996), .A2(n909), .ZN(n952) );
  NAND2_X1 U687 ( .A1(G107), .A2(n599), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G131), .A2(n903), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U690 ( .A1(G95), .A2(n902), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G119), .A2(n884), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n895) );
  NAND2_X1 U694 ( .A1(G1991), .A2(n895), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(KEYINPUT88), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G1996), .A2(n909), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U698 ( .A(KEYINPUT90), .B(n625), .ZN(n971) );
  NOR2_X1 U699 ( .A1(G1986), .A2(G290), .ZN(n627) );
  NOR2_X1 U700 ( .A1(G1991), .A2(n895), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT105), .B(n626), .Z(n957) );
  NOR2_X1 U702 ( .A1(n627), .A2(n957), .ZN(n628) );
  NOR2_X1 U703 ( .A1(n971), .A2(n628), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n952), .A2(n629), .ZN(n630) );
  XOR2_X1 U705 ( .A(KEYINPUT39), .B(n630), .Z(n631) );
  NOR2_X1 U706 ( .A1(n959), .A2(n631), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n958), .A2(n632), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n760) );
  INV_X1 U709 ( .A(n635), .ZN(n636) );
  NOR2_X4 U710 ( .A1(n637), .A2(n636), .ZN(n677) );
  INV_X1 U711 ( .A(n677), .ZN(n661) );
  NAND2_X1 U712 ( .A1(G8), .A2(n661), .ZN(n737) );
  NOR2_X1 U713 ( .A1(G305), .A2(G1981), .ZN(n638) );
  XOR2_X1 U714 ( .A(n638), .B(KEYINPUT24), .Z(n639) );
  NOR2_X1 U715 ( .A1(n737), .A2(n639), .ZN(n750) );
  NOR2_X1 U716 ( .A1(G2090), .A2(G303), .ZN(n640) );
  XNOR2_X1 U717 ( .A(KEYINPUT102), .B(n640), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n641), .A2(G8), .ZN(n727) );
  INV_X1 U719 ( .A(n661), .ZN(n664) );
  NOR2_X1 U720 ( .A1(n664), .A2(G1961), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n642), .B(KEYINPUT91), .ZN(n644) );
  XNOR2_X1 U722 ( .A(G2078), .B(KEYINPUT25), .ZN(n1010) );
  NAND2_X1 U723 ( .A1(n677), .A2(n1010), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n697) );
  NAND2_X1 U725 ( .A1(n697), .A2(G171), .ZN(n691) );
  NAND2_X1 U726 ( .A1(G66), .A2(n805), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G92), .A2(n810), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U729 ( .A1(G79), .A2(n809), .ZN(n648) );
  NAND2_X1 U730 ( .A1(G54), .A2(n806), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U733 ( .A(KEYINPUT15), .B(n651), .ZN(n978) );
  INV_X1 U734 ( .A(n978), .ZN(n847) );
  NAND2_X1 U735 ( .A1(G56), .A2(n805), .ZN(n652) );
  XOR2_X1 U736 ( .A(KEYINPUT14), .B(n652), .Z(n658) );
  NAND2_X1 U737 ( .A1(G81), .A2(n810), .ZN(n653) );
  XNOR2_X1 U738 ( .A(n653), .B(KEYINPUT12), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G68), .A2(n809), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U741 ( .A(KEYINPUT13), .B(n656), .Z(n657) );
  NOR2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U743 ( .A1(n806), .A2(G43), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n800) );
  INV_X1 U745 ( .A(G1996), .ZN(n863) );
  NOR2_X1 U746 ( .A1(n661), .A2(n863), .ZN(n663) );
  XNOR2_X1 U747 ( .A(n663), .B(n662), .ZN(n666) );
  INV_X1 U748 ( .A(n664), .ZN(n707) );
  NAND2_X1 U749 ( .A1(n707), .A2(G1341), .ZN(n665) );
  NAND2_X1 U750 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U751 ( .A1(n800), .A2(n667), .ZN(n668) );
  OR2_X1 U752 ( .A1(n847), .A2(n668), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n847), .A2(n668), .ZN(n673) );
  NAND2_X1 U754 ( .A1(G1348), .A2(n707), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n677), .A2(G2067), .ZN(n669) );
  NAND2_X1 U756 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U757 ( .A(KEYINPUT93), .B(n671), .Z(n672) );
  NAND2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n677), .A2(G2072), .ZN(n676) );
  XNOR2_X1 U761 ( .A(n676), .B(KEYINPUT27), .ZN(n679) );
  INV_X1 U762 ( .A(G1956), .ZN(n980) );
  NOR2_X1 U763 ( .A1(n980), .A2(n677), .ZN(n678) );
  NOR2_X1 U764 ( .A1(n679), .A2(n678), .ZN(n683) );
  INV_X1 U765 ( .A(G299), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n683), .A2(n682), .ZN(n680) );
  NAND2_X1 U767 ( .A1(n681), .A2(n680), .ZN(n687) );
  NOR2_X1 U768 ( .A1(n683), .A2(n682), .ZN(n685) );
  XOR2_X1 U769 ( .A(KEYINPUT28), .B(KEYINPUT92), .Z(n684) );
  XNOR2_X1 U770 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n689) );
  XOR2_X1 U772 ( .A(KEYINPUT29), .B(KEYINPUT94), .Z(n688) );
  XNOR2_X1 U773 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n691), .A2(n690), .ZN(n715) );
  NOR2_X1 U775 ( .A1(G1966), .A2(n737), .ZN(n702) );
  NOR2_X1 U776 ( .A1(G2084), .A2(n707), .ZN(n701) );
  NOR2_X1 U777 ( .A1(n702), .A2(n701), .ZN(n692) );
  NAND2_X1 U778 ( .A1(G8), .A2(n692), .ZN(n695) );
  XOR2_X1 U779 ( .A(KEYINPUT30), .B(KEYINPUT95), .Z(n693) );
  NOR2_X1 U780 ( .A1(G168), .A2(n696), .ZN(n699) );
  NOR2_X1 U781 ( .A1(G171), .A2(n697), .ZN(n698) );
  NOR2_X1 U782 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U783 ( .A(KEYINPUT31), .B(n700), .Z(n716) );
  AND2_X1 U784 ( .A1(n715), .A2(n716), .ZN(n705) );
  AND2_X1 U785 ( .A1(G8), .A2(n701), .ZN(n703) );
  OR2_X1 U786 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U787 ( .A(n706), .B(KEYINPUT97), .ZN(n725) );
  INV_X1 U788 ( .A(G8), .ZN(n714) );
  NOR2_X1 U789 ( .A1(G2090), .A2(n707), .ZN(n708) );
  XOR2_X1 U790 ( .A(KEYINPUT98), .B(n708), .Z(n709) );
  NAND2_X1 U791 ( .A1(n709), .A2(G303), .ZN(n711) );
  NOR2_X1 U792 ( .A1(G1971), .A2(n737), .ZN(n710) );
  NOR2_X1 U793 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U794 ( .A(n712), .B(KEYINPUT99), .ZN(n713) );
  OR2_X1 U795 ( .A1(n714), .A2(n713), .ZN(n718) );
  AND2_X1 U796 ( .A1(n715), .A2(n718), .ZN(n717) );
  NAND2_X1 U797 ( .A1(n717), .A2(n716), .ZN(n722) );
  INV_X1 U798 ( .A(n718), .ZN(n720) );
  AND2_X1 U799 ( .A1(G286), .A2(G8), .ZN(n719) );
  OR2_X1 U800 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U801 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U802 ( .A(n723), .B(KEYINPUT32), .ZN(n724) );
  NAND2_X1 U803 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U804 ( .A1(n727), .A2(n735), .ZN(n728) );
  NAND2_X1 U805 ( .A1(n737), .A2(n728), .ZN(n729) );
  XNOR2_X1 U806 ( .A(n729), .B(KEYINPUT103), .ZN(n730) );
  NOR2_X1 U807 ( .A1(G1971), .A2(G303), .ZN(n731) );
  NOR2_X1 U808 ( .A1(G1976), .A2(G288), .ZN(n985) );
  NOR2_X1 U809 ( .A1(n731), .A2(n985), .ZN(n733) );
  INV_X1 U810 ( .A(KEYINPUT33), .ZN(n732) );
  AND2_X1 U811 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U812 ( .A1(n735), .A2(n734), .ZN(n743) );
  XOR2_X1 U813 ( .A(G305), .B(G1981), .Z(n998) );
  NAND2_X1 U814 ( .A1(G1976), .A2(G288), .ZN(n986) );
  INV_X1 U815 ( .A(n986), .ZN(n736) );
  NOR2_X1 U816 ( .A1(KEYINPUT33), .A2(n515), .ZN(n740) );
  NAND2_X1 U817 ( .A1(n985), .A2(KEYINPUT33), .ZN(n738) );
  NOR2_X1 U818 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U819 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U820 ( .A1(n998), .A2(n741), .ZN(n742) );
  NAND2_X1 U821 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U822 ( .A(n744), .B(KEYINPUT101), .ZN(n745) );
  NOR2_X1 U823 ( .A1(n750), .A2(n749), .ZN(n758) );
  XNOR2_X1 U824 ( .A(KEYINPUT82), .B(G1986), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n751), .B(G290), .ZN(n982) );
  NAND2_X1 U826 ( .A1(n982), .A2(n753), .ZN(n752) );
  XNOR2_X1 U827 ( .A(n752), .B(KEYINPUT84), .ZN(n756) );
  OR2_X1 U828 ( .A1(n971), .A2(n959), .ZN(n754) );
  NAND2_X1 U829 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U830 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U832 ( .A1(n760), .A2(n759), .ZN(n763) );
  INV_X1 U833 ( .A(KEYINPUT40), .ZN(n761) );
  XNOR2_X1 U834 ( .A(n763), .B(n762), .ZN(G329) );
  XOR2_X1 U835 ( .A(KEYINPUT107), .B(G2435), .Z(n765) );
  XNOR2_X1 U836 ( .A(G2430), .B(G2438), .ZN(n764) );
  XNOR2_X1 U837 ( .A(n765), .B(n764), .ZN(n772) );
  XOR2_X1 U838 ( .A(G2446), .B(G2454), .Z(n767) );
  XNOR2_X1 U839 ( .A(G2451), .B(G2443), .ZN(n766) );
  XNOR2_X1 U840 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U841 ( .A(n768), .B(G2427), .Z(n770) );
  XNOR2_X1 U842 ( .A(G1341), .B(G1348), .ZN(n769) );
  XNOR2_X1 U843 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U844 ( .A(n772), .B(n771), .ZN(n773) );
  AND2_X1 U845 ( .A1(n773), .A2(G14), .ZN(G401) );
  INV_X1 U846 ( .A(G171), .ZN(G301) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U848 ( .A1(G111), .A2(n599), .ZN(n775) );
  NAND2_X1 U849 ( .A1(G135), .A2(n903), .ZN(n774) );
  NAND2_X1 U850 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U851 ( .A1(n884), .A2(G123), .ZN(n776) );
  XOR2_X1 U852 ( .A(KEYINPUT18), .B(n776), .Z(n777) );
  NOR2_X1 U853 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U854 ( .A1(n902), .A2(G99), .ZN(n779) );
  NAND2_X1 U855 ( .A1(n780), .A2(n779), .ZN(n954) );
  XNOR2_X1 U856 ( .A(G2096), .B(n954), .ZN(n781) );
  OR2_X1 U857 ( .A1(G2100), .A2(n781), .ZN(G156) );
  INV_X1 U858 ( .A(G132), .ZN(G219) );
  INV_X1 U859 ( .A(G57), .ZN(G237) );
  INV_X1 U860 ( .A(G108), .ZN(G238) );
  INV_X1 U861 ( .A(G69), .ZN(G235) );
  AND2_X1 U862 ( .A1(n903), .A2(G138), .ZN(n784) );
  NOR2_X1 U863 ( .A1(n784), .A2(n783), .ZN(G164) );
  XOR2_X1 U864 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n786) );
  NAND2_X1 U865 ( .A1(G7), .A2(G661), .ZN(n785) );
  XOR2_X1 U866 ( .A(n786), .B(n785), .Z(n842) );
  NAND2_X1 U867 ( .A1(n842), .A2(G567), .ZN(n787) );
  XOR2_X1 U868 ( .A(KEYINPUT11), .B(n787), .Z(G234) );
  INV_X1 U869 ( .A(n800), .ZN(n989) );
  NAND2_X1 U870 ( .A1(n989), .A2(G860), .ZN(G153) );
  INV_X1 U871 ( .A(G868), .ZN(n824) );
  NAND2_X1 U872 ( .A1(n978), .A2(n824), .ZN(n788) );
  XNOR2_X1 U873 ( .A(n788), .B(KEYINPUT72), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G868), .A2(G301), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n790), .A2(n789), .ZN(G284) );
  NOR2_X1 U876 ( .A1(G286), .A2(n824), .ZN(n792) );
  NOR2_X1 U877 ( .A1(G868), .A2(G299), .ZN(n791) );
  NOR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(G297) );
  INV_X1 U879 ( .A(G559), .ZN(n793) );
  NOR2_X1 U880 ( .A1(G860), .A2(n793), .ZN(n794) );
  XNOR2_X1 U881 ( .A(KEYINPUT73), .B(n794), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n795), .A2(n847), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n796), .B(KEYINPUT74), .ZN(n797) );
  XNOR2_X1 U884 ( .A(KEYINPUT16), .B(n797), .ZN(G148) );
  NOR2_X1 U885 ( .A1(n978), .A2(n824), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(KEYINPUT75), .ZN(n799) );
  NOR2_X1 U887 ( .A1(G559), .A2(n799), .ZN(n802) );
  NOR2_X1 U888 ( .A1(G868), .A2(n800), .ZN(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U890 ( .A(KEYINPUT76), .B(n803), .ZN(G282) );
  NAND2_X1 U891 ( .A1(n847), .A2(G559), .ZN(n822) );
  XOR2_X1 U892 ( .A(n989), .B(n822), .Z(n804) );
  NOR2_X1 U893 ( .A1(n804), .A2(G860), .ZN(n815) );
  NAND2_X1 U894 ( .A1(G67), .A2(n805), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G55), .A2(n806), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n814) );
  NAND2_X1 U897 ( .A1(G80), .A2(n809), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G93), .A2(n810), .ZN(n811) );
  NAND2_X1 U899 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U900 ( .A1(n814), .A2(n813), .ZN(n825) );
  XOR2_X1 U901 ( .A(n815), .B(n825), .Z(G145) );
  XOR2_X1 U902 ( .A(n825), .B(G290), .Z(n818) );
  XOR2_X1 U903 ( .A(G303), .B(KEYINPUT19), .Z(n816) );
  XNOR2_X1 U904 ( .A(n816), .B(G288), .ZN(n817) );
  XNOR2_X1 U905 ( .A(n818), .B(n817), .ZN(n819) );
  XOR2_X1 U906 ( .A(n989), .B(n819), .Z(n821) );
  XOR2_X1 U907 ( .A(G305), .B(G299), .Z(n820) );
  XNOR2_X1 U908 ( .A(n821), .B(n820), .ZN(n846) );
  XNOR2_X1 U909 ( .A(n846), .B(n822), .ZN(n823) );
  NOR2_X1 U910 ( .A1(n824), .A2(n823), .ZN(n827) );
  NOR2_X1 U911 ( .A1(G868), .A2(n825), .ZN(n826) );
  NOR2_X1 U912 ( .A1(n827), .A2(n826), .ZN(G295) );
  NAND2_X1 U913 ( .A1(G2078), .A2(G2084), .ZN(n828) );
  XOR2_X1 U914 ( .A(KEYINPUT20), .B(n828), .Z(n829) );
  NAND2_X1 U915 ( .A1(G2090), .A2(n829), .ZN(n830) );
  XNOR2_X1 U916 ( .A(KEYINPUT21), .B(n830), .ZN(n831) );
  NAND2_X1 U917 ( .A1(n831), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U918 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U919 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U920 ( .A1(G235), .A2(G238), .ZN(n832) );
  NAND2_X1 U921 ( .A1(G120), .A2(n832), .ZN(n833) );
  NOR2_X1 U922 ( .A1(n833), .A2(G237), .ZN(n834) );
  XNOR2_X1 U923 ( .A(n834), .B(KEYINPUT81), .ZN(n924) );
  AND2_X1 U924 ( .A1(G567), .A2(n924), .ZN(n840) );
  NOR2_X1 U925 ( .A1(G220), .A2(G219), .ZN(n835) );
  XOR2_X1 U926 ( .A(KEYINPUT22), .B(n835), .Z(n836) );
  NOR2_X1 U927 ( .A1(G218), .A2(n836), .ZN(n837) );
  NAND2_X1 U928 ( .A1(G96), .A2(n837), .ZN(n925) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n925), .ZN(n838) );
  XOR2_X1 U930 ( .A(KEYINPUT80), .B(n838), .Z(n839) );
  NOR2_X1 U931 ( .A1(n840), .A2(n839), .ZN(G319) );
  INV_X1 U932 ( .A(G319), .ZN(n919) );
  NAND2_X1 U933 ( .A1(G483), .A2(G661), .ZN(n841) );
  NOR2_X1 U934 ( .A1(n919), .A2(n841), .ZN(n845) );
  NAND2_X1 U935 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n842), .ZN(G217) );
  INV_X1 U937 ( .A(n842), .ZN(G223) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U939 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n845), .A2(n844), .ZN(G188) );
  XOR2_X1 U942 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  XOR2_X1 U943 ( .A(n846), .B(G286), .Z(n849) );
  XOR2_X1 U944 ( .A(G301), .B(n847), .Z(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n850) );
  NOR2_X1 U946 ( .A1(G37), .A2(n850), .ZN(G397) );
  XOR2_X1 U947 ( .A(G2096), .B(G2090), .Z(n852) );
  XNOR2_X1 U948 ( .A(G2072), .B(G2067), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n862) );
  XOR2_X1 U950 ( .A(KEYINPUT111), .B(G2678), .Z(n854) );
  XNOR2_X1 U951 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U953 ( .A(G2100), .B(KEYINPUT112), .Z(n856) );
  XNOR2_X1 U954 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U956 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U959 ( .A(n862), .B(n861), .Z(G227) );
  XNOR2_X1 U960 ( .A(G1991), .B(n863), .ZN(n865) );
  XNOR2_X1 U961 ( .A(G1981), .B(G1966), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n875) );
  XOR2_X1 U963 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n867) );
  XNOR2_X1 U964 ( .A(G1986), .B(KEYINPUT41), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n871) );
  XNOR2_X1 U966 ( .A(n980), .B(G1961), .ZN(n869) );
  XNOR2_X1 U967 ( .A(G1976), .B(G1971), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U970 ( .A(KEYINPUT114), .B(G2474), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G124), .A2(n884), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U975 ( .A1(n599), .A2(G112), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G100), .A2(n902), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G136), .A2(n903), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U980 ( .A1(n882), .A2(n881), .ZN(G162) );
  XOR2_X1 U981 ( .A(G164), .B(G162), .Z(n883) );
  XNOR2_X1 U982 ( .A(n954), .B(n883), .ZN(n899) );
  NAND2_X1 U983 ( .A1(G115), .A2(n599), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G127), .A2(n884), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n887), .B(KEYINPUT47), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G103), .A2(n902), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n903), .A2(G139), .ZN(n890) );
  XOR2_X1 U990 ( .A(KEYINPUT118), .B(n890), .Z(n891) );
  NOR2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n962) );
  XNOR2_X1 U992 ( .A(n962), .B(KEYINPUT117), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n893), .B(KEYINPUT48), .ZN(n894) );
  XNOR2_X1 U994 ( .A(KEYINPUT119), .B(n894), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n895), .B(KEYINPUT46), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n899), .B(n898), .Z(n913) );
  NAND2_X1 U998 ( .A1(G118), .A2(n599), .ZN(n901) );
  NAND2_X1 U999 ( .A1(G130), .A2(n884), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n902), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(G142), .A2(n903), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n906), .B(KEYINPUT45), .Z(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(G160), .B(n911), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G397), .A2(n918), .ZN(n923) );
  NOR2_X1 U1014 ( .A1(n919), .A2(G401), .ZN(n920) );
  XOR2_X1 U1015 ( .A(KEYINPUT120), .B(n920), .Z(n921) );
  NOR2_X1 U1016 ( .A1(G395), .A2(n921), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(G225) );
  XNOR2_X1 U1018 ( .A(KEYINPUT121), .B(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1022 ( .A(n926), .B(KEYINPUT109), .Z(G325) );
  INV_X1 U1023 ( .A(G325), .ZN(G261) );
  INV_X1 U1024 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1025 ( .A(G16), .B(KEYINPUT126), .Z(n949) );
  XNOR2_X1 U1026 ( .A(KEYINPUT127), .B(G1966), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(n927), .B(G21), .ZN(n939) );
  XOR2_X1 U1028 ( .A(G20), .B(G1956), .Z(n931) );
  XNOR2_X1 U1029 ( .A(G1981), .B(G6), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G19), .B(G1341), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT59), .B(G1348), .Z(n932) );
  XNOR2_X1 U1034 ( .A(G4), .B(n932), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1036 ( .A(KEYINPUT60), .B(n935), .Z(n937) );
  XNOR2_X1 U1037 ( .A(G1961), .B(G5), .ZN(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G1971), .B(G22), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(G24), .B(G1986), .ZN(n940) );
  NOR2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n943) );
  XOR2_X1 U1043 ( .A(G1976), .B(G23), .Z(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(KEYINPUT58), .B(n944), .ZN(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(n947), .B(KEYINPUT61), .ZN(n948) );
  NAND2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n950), .ZN(n977) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n953), .Z(n969) );
  XNOR2_X1 U1053 ( .A(G160), .B(G2084), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n967) );
  XOR2_X1 U1058 ( .A(G2072), .B(n962), .Z(n964) );
  XOR2_X1 U1059 ( .A(G164), .B(G2078), .Z(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1061 ( .A(KEYINPUT50), .B(n965), .Z(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(KEYINPUT52), .B(n972), .ZN(n973) );
  INV_X1 U1066 ( .A(KEYINPUT55), .ZN(n1025) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n1025), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n974), .A2(G29), .ZN(n975) );
  XOR2_X1 U1069 ( .A(KEYINPUT122), .B(n975), .Z(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n1006) );
  XNOR2_X1 U1071 ( .A(KEYINPUT56), .B(G16), .ZN(n1004) );
  XOR2_X1 U1072 ( .A(G1348), .B(n978), .Z(n979) );
  XNOR2_X1 U1073 ( .A(n979), .B(KEYINPUT124), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G299), .B(n980), .Z(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n997) );
  XOR2_X1 U1077 ( .A(G301), .B(G1961), .Z(n995) );
  INV_X1 U1078 ( .A(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(n988), .B(KEYINPUT125), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G1341), .B(n989), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(G1971), .B(G303), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G168), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(n1000), .B(KEYINPUT57), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1028) );
  XNOR2_X1 U1093 ( .A(G2072), .B(G33), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(G2067), .B(G26), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1016) );
  XOR2_X1 U1096 ( .A(G1991), .B(G25), .Z(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(G28), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(G1996), .B(G32), .Z(n1012) );
  XNOR2_X1 U1099 ( .A(n1010), .B(G27), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1017), .B(KEYINPUT53), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(G2084), .B(KEYINPUT54), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(G34), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(KEYINPUT123), .B(G2090), .Z(n1021) );
  XNOR2_X1 U1108 ( .A(G35), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(n1025), .B(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(G29), .A2(n1026), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(n1029), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1114 ( .A(G150), .ZN(G311) );
endmodule

