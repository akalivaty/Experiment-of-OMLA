

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590;

  XNOR2_X1 U322 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U323 ( .A(n375), .B(n374), .Z(n290) );
  NOR2_X1 U324 ( .A1(n390), .A2(n577), .ZN(n391) );
  XNOR2_X1 U325 ( .A(n395), .B(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U326 ( .A(n397), .B(n396), .ZN(n529) );
  XNOR2_X1 U327 ( .A(n447), .B(KEYINPUT117), .ZN(n448) );
  XNOR2_X1 U328 ( .A(n376), .B(n290), .ZN(n377) );
  XNOR2_X1 U329 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U330 ( .A(n451), .B(G190GAT), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(G190GAT), .B(G134GAT), .Z(n368) );
  XOR2_X1 U333 ( .A(G120GAT), .B(G71GAT), .Z(n326) );
  XNOR2_X1 U334 ( .A(n368), .B(n326), .ZN(n293) );
  XOR2_X1 U335 ( .A(G127GAT), .B(KEYINPUT0), .Z(n292) );
  XNOR2_X1 U336 ( .A(G113GAT), .B(KEYINPUT84), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n443) );
  XNOR2_X1 U338 ( .A(n293), .B(n443), .ZN(n299) );
  XOR2_X1 U339 ( .A(G183GAT), .B(KEYINPUT17), .Z(n295) );
  XNOR2_X1 U340 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n408) );
  XOR2_X1 U342 ( .A(G15GAT), .B(n408), .Z(n297) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U345 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U346 ( .A(G176GAT), .B(G99GAT), .Z(n301) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(G43GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U349 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n303) );
  XNOR2_X1 U350 ( .A(KEYINPUT87), .B(KEYINPUT20), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(n307), .B(n306), .Z(n510) );
  INV_X1 U354 ( .A(n510), .ZN(n532) );
  XOR2_X1 U355 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n309) );
  XNOR2_X1 U356 ( .A(KEYINPUT68), .B(KEYINPUT71), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U358 ( .A(G113GAT), .B(G197GAT), .Z(n311) );
  XOR2_X1 U359 ( .A(G141GAT), .B(G22GAT), .Z(n417) );
  XOR2_X1 U360 ( .A(G169GAT), .B(G8GAT), .Z(n401) );
  XNOR2_X1 U361 ( .A(n417), .B(n401), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U363 ( .A(n313), .B(n312), .Z(n315) );
  NAND2_X1 U364 ( .A1(G229GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U366 ( .A(n316), .B(KEYINPUT30), .Z(n319) );
  XNOR2_X1 U367 ( .A(G15GAT), .B(G1GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n317), .B(KEYINPUT69), .ZN(n358) );
  XNOR2_X1 U369 ( .A(n358), .B(KEYINPUT29), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U371 ( .A(G29GAT), .B(KEYINPUT7), .Z(n321) );
  XNOR2_X1 U372 ( .A(G43GAT), .B(G36GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U374 ( .A(G50GAT), .B(KEYINPUT8), .Z(n322) );
  XOR2_X1 U375 ( .A(n323), .B(n322), .Z(n380) );
  XOR2_X1 U376 ( .A(n324), .B(n380), .Z(n574) );
  XNOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n325), .B(KEYINPUT73), .ZN(n362) );
  XNOR2_X1 U379 ( .A(n362), .B(n326), .ZN(n330) );
  INV_X1 U380 ( .A(n330), .ZN(n328) );
  AND2_X1 U381 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  INV_X1 U382 ( .A(n329), .ZN(n327) );
  NAND2_X1 U383 ( .A1(n328), .A2(n327), .ZN(n332) );
  NAND2_X1 U384 ( .A1(n330), .A2(n329), .ZN(n331) );
  NAND2_X1 U385 ( .A1(n332), .A2(n331), .ZN(n333) );
  XOR2_X1 U386 ( .A(n333), .B(KEYINPUT31), .Z(n336) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n334), .B(KEYINPUT75), .ZN(n367) );
  XNOR2_X1 U389 ( .A(n367), .B(KEYINPUT32), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U391 ( .A(KEYINPUT76), .B(KEYINPUT74), .Z(n338) );
  XNOR2_X1 U392 ( .A(KEYINPUT77), .B(KEYINPUT33), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n345) );
  XOR2_X1 U395 ( .A(G78GAT), .B(G148GAT), .Z(n342) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(G204GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n412) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(G92GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n343), .B(G64GAT), .ZN(n404) );
  XNOR2_X1 U400 ( .A(n412), .B(n404), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n577) );
  XOR2_X1 U402 ( .A(n577), .B(KEYINPUT41), .Z(n560) );
  NAND2_X1 U403 ( .A1(n574), .A2(n560), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n346), .B(KEYINPUT46), .ZN(n385) );
  XOR2_X1 U405 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n348) );
  XNOR2_X1 U406 ( .A(KEYINPUT81), .B(KEYINPUT15), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n366) );
  XOR2_X1 U408 ( .A(G78GAT), .B(G211GAT), .Z(n350) );
  XNOR2_X1 U409 ( .A(G183GAT), .B(G71GAT), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U411 ( .A(KEYINPUT80), .B(G64GAT), .Z(n352) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(G127GAT), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U414 ( .A(n354), .B(n353), .Z(n360) );
  XOR2_X1 U415 ( .A(G155GAT), .B(G22GAT), .Z(n356) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U420 ( .A(n361), .B(KEYINPUT82), .Z(n364) );
  XNOR2_X1 U421 ( .A(n362), .B(KEYINPUT12), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U423 ( .A(n366), .B(n365), .Z(n581) );
  INV_X1 U424 ( .A(KEYINPUT47), .ZN(n381) );
  XOR2_X1 U425 ( .A(n367), .B(G106GAT), .Z(n370) );
  XNOR2_X1 U426 ( .A(n368), .B(G218GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n378) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n372) );
  XNOR2_X1 U429 ( .A(G92GAT), .B(KEYINPUT78), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U431 ( .A(G162GAT), .B(n373), .ZN(n376) );
  XOR2_X1 U432 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n375) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n553) );
  OR2_X1 U435 ( .A1(n381), .A2(n553), .ZN(n382) );
  NOR2_X1 U436 ( .A1(n581), .A2(n382), .ZN(n383) );
  NAND2_X1 U437 ( .A1(n385), .A2(n383), .ZN(n388) );
  NOR2_X1 U438 ( .A1(n553), .A2(n581), .ZN(n384) );
  NAND2_X1 U439 ( .A1(n385), .A2(n384), .ZN(n386) );
  NAND2_X1 U440 ( .A1(n386), .A2(n381), .ZN(n387) );
  NAND2_X1 U441 ( .A1(n388), .A2(n387), .ZN(n394) );
  XOR2_X1 U442 ( .A(KEYINPUT36), .B(n553), .Z(n588) );
  INV_X1 U443 ( .A(n581), .ZN(n482) );
  NOR2_X1 U444 ( .A1(n588), .A2(n482), .ZN(n389) );
  XOR2_X1 U445 ( .A(KEYINPUT45), .B(n389), .Z(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT110), .B(n391), .ZN(n392) );
  INV_X1 U447 ( .A(n574), .ZN(n499) );
  XOR2_X1 U448 ( .A(n499), .B(KEYINPUT72), .Z(n556) );
  INV_X1 U449 ( .A(n556), .ZN(n454) );
  NAND2_X1 U450 ( .A1(n392), .A2(n454), .ZN(n393) );
  NAND2_X1 U451 ( .A1(n394), .A2(n393), .ZN(n397) );
  XNOR2_X1 U452 ( .A(KEYINPUT64), .B(KEYINPUT111), .ZN(n395) );
  XOR2_X1 U453 ( .A(KEYINPUT93), .B(G204GAT), .Z(n399) );
  XNOR2_X1 U454 ( .A(G36GAT), .B(G190GAT), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U456 ( .A(n401), .B(n400), .Z(n403) );
  NAND2_X1 U457 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U459 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U460 ( .A(G211GAT), .B(KEYINPUT21), .Z(n407) );
  XNOR2_X1 U461 ( .A(G197GAT), .B(G218GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n413) );
  XNOR2_X1 U463 ( .A(n408), .B(n413), .ZN(n409) );
  XOR2_X1 U464 ( .A(n410), .B(n409), .Z(n506) );
  INV_X1 U465 ( .A(n506), .ZN(n521) );
  NOR2_X1 U466 ( .A1(n529), .A2(n521), .ZN(n411) );
  XNOR2_X1 U467 ( .A(KEYINPUT54), .B(n411), .ZN(n571) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n426) );
  XOR2_X1 U469 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n415) );
  XNOR2_X1 U470 ( .A(G50GAT), .B(KEYINPUT88), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U472 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U475 ( .A(n420), .B(KEYINPUT89), .Z(n424) );
  XOR2_X1 U476 ( .A(G155GAT), .B(KEYINPUT2), .Z(n422) );
  XNOR2_X1 U477 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n442) );
  XNOR2_X1 U479 ( .A(n442), .B(KEYINPUT23), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n461) );
  XOR2_X1 U482 ( .A(G85GAT), .B(G134GAT), .Z(n428) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(G141GAT), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U485 ( .A(G57GAT), .B(G148GAT), .Z(n430) );
  XNOR2_X1 U486 ( .A(G1GAT), .B(G120GAT), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U488 ( .A(n432), .B(n431), .Z(n437) );
  XOR2_X1 U489 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n434) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U492 ( .A(KEYINPUT91), .B(n435), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U494 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n439) );
  XNOR2_X1 U495 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U497 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n503) );
  NOR2_X1 U500 ( .A1(n461), .A2(n503), .ZN(n446) );
  AND2_X1 U501 ( .A1(n571), .A2(n446), .ZN(n449) );
  INV_X1 U502 ( .A(KEYINPUT55), .ZN(n447) );
  NOR2_X1 U503 ( .A1(n532), .A2(n450), .ZN(n565) );
  NAND2_X1 U504 ( .A1(n565), .A2(n553), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n451) );
  INV_X1 U506 ( .A(n503), .ZN(n570) );
  NOR2_X1 U507 ( .A1(n454), .A2(n577), .ZN(n485) );
  XOR2_X1 U508 ( .A(n506), .B(KEYINPUT27), .Z(n464) );
  NOR2_X1 U509 ( .A1(n570), .A2(n464), .ZN(n455) );
  XOR2_X1 U510 ( .A(KEYINPUT94), .B(n455), .Z(n528) );
  XOR2_X1 U511 ( .A(n461), .B(KEYINPUT66), .Z(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT28), .B(n456), .Z(n514) );
  INV_X1 U513 ( .A(n514), .ZN(n530) );
  NAND2_X1 U514 ( .A1(n532), .A2(n530), .ZN(n457) );
  NOR2_X1 U515 ( .A1(n528), .A2(n457), .ZN(n469) );
  NOR2_X1 U516 ( .A1(n532), .A2(n521), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n461), .A2(n458), .ZN(n459) );
  XOR2_X1 U518 ( .A(n459), .B(KEYINPUT96), .Z(n460) );
  XNOR2_X1 U519 ( .A(KEYINPUT25), .B(n460), .ZN(n466) );
  XOR2_X1 U520 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n463) );
  NAND2_X1 U521 ( .A1(n461), .A2(n532), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(n573) );
  NOR2_X1 U523 ( .A1(n573), .A2(n464), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n467), .A2(n503), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n480) );
  XOR2_X1 U527 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n471) );
  OR2_X1 U528 ( .A1(n482), .A2(n553), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n471), .B(n470), .ZN(n472) );
  NOR2_X1 U530 ( .A1(n480), .A2(n472), .ZN(n501) );
  NAND2_X1 U531 ( .A1(n485), .A2(n501), .ZN(n478) );
  NOR2_X1 U532 ( .A1(n570), .A2(n478), .ZN(n473) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n473), .Z(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(n474), .ZN(G1324GAT) );
  NOR2_X1 U535 ( .A1(n521), .A2(n478), .ZN(n475) );
  XOR2_X1 U536 ( .A(G8GAT), .B(n475), .Z(G1325GAT) );
  NOR2_X1 U537 ( .A1(n532), .A2(n478), .ZN(n477) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n530), .A2(n478), .ZN(n479) );
  XOR2_X1 U541 ( .A(G22GAT), .B(n479), .Z(G1327GAT) );
  XNOR2_X1 U542 ( .A(KEYINPUT98), .B(KEYINPUT38), .ZN(n487) );
  NOR2_X1 U543 ( .A1(n480), .A2(n588), .ZN(n481) );
  NAND2_X1 U544 ( .A1(n482), .A2(n481), .ZN(n483) );
  XOR2_X1 U545 ( .A(KEYINPUT37), .B(n483), .Z(n484) );
  XNOR2_X1 U546 ( .A(KEYINPUT97), .B(n484), .ZN(n518) );
  NAND2_X1 U547 ( .A1(n518), .A2(n485), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n497) );
  NOR2_X1 U549 ( .A1(n497), .A2(n570), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n489) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U554 ( .A1(n521), .A2(n497), .ZN(n492) );
  XOR2_X1 U555 ( .A(G36GAT), .B(n492), .Z(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n494) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n496) );
  NOR2_X1 U559 ( .A1(n532), .A2(n497), .ZN(n495) );
  XOR2_X1 U560 ( .A(n496), .B(n495), .Z(G1330GAT) );
  NOR2_X1 U561 ( .A1(n530), .A2(n497), .ZN(n498) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n498), .Z(G1331GAT) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n505) );
  NAND2_X1 U564 ( .A1(n560), .A2(n499), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(KEYINPUT103), .ZN(n517) );
  NAND2_X1 U566 ( .A1(n501), .A2(n517), .ZN(n502) );
  XOR2_X1 U567 ( .A(KEYINPUT104), .B(n502), .Z(n513) );
  NAND2_X1 U568 ( .A1(n503), .A2(n513), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n508) );
  NAND2_X1 U571 ( .A1(n513), .A2(n506), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT107), .Z(n512) );
  NAND2_X1 U575 ( .A1(n513), .A2(n510), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U578 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U581 ( .A1(n570), .A2(n525), .ZN(n519) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n519), .Z(n520) );
  XNOR2_X1 U583 ( .A(KEYINPUT108), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n525), .ZN(n523) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n532), .A2(n525), .ZN(n524) );
  XOR2_X1 U588 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U589 ( .A1(n530), .A2(n525), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(n526), .Z(n527) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT112), .ZN(n534) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n542), .A2(n530), .ZN(n531) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n539), .A2(n556), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U599 ( .A1(n539), .A2(n560), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n539), .A2(n581), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U605 ( .A1(n539), .A2(n553), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n545) );
  INV_X1 U608 ( .A(n542), .ZN(n543) );
  NOR2_X1 U609 ( .A1(n573), .A2(n543), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n552), .A2(n574), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U614 ( .A1(n552), .A2(n560), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT115), .Z(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n581), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT116), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n565), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n565), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n581), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n568) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT122), .B(n569), .Z(n576) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n586) );
  NAND2_X1 U640 ( .A1(n586), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U643 ( .A1(n586), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT125), .Z(n583) );
  NAND2_X1 U647 ( .A1(n586), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n585) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n590) );
  INV_X1 U652 ( .A(n586), .ZN(n587) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U654 ( .A(n590), .B(n589), .Z(G1355GAT) );
endmodule

