

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749;

  AND2_X1 U367 ( .A1(n375), .A2(n373), .ZN(n372) );
  XNOR2_X1 U368 ( .A(n366), .B(G137), .ZN(n728) );
  INV_X2 U369 ( .A(G143), .ZN(n447) );
  NOR2_X1 U370 ( .A1(G953), .A2(G237), .ZN(n510) );
  INV_X1 U371 ( .A(n549), .ZN(n589) );
  OR2_X1 U372 ( .A1(n493), .A2(n374), .ZN(n373) );
  XNOR2_X1 U373 ( .A(n606), .B(KEYINPUT104), .ZN(n417) );
  XNOR2_X1 U374 ( .A(n402), .B(n503), .ZN(n723) );
  NOR2_X1 U375 ( .A1(n568), .A2(n645), .ZN(n391) );
  BUF_X1 U376 ( .A(n532), .Z(n563) );
  INV_X2 U377 ( .A(G953), .ZN(n494) );
  AND2_X2 U378 ( .A1(n630), .A2(n615), .ZN(n633) );
  AND2_X2 U379 ( .A1(n616), .A2(n615), .ZN(n618) );
  AND2_X2 U380 ( .A1(n408), .A2(n421), .ZN(n407) );
  XNOR2_X2 U381 ( .A(n423), .B(n611), .ZN(n704) );
  NAND2_X2 U382 ( .A1(n407), .A2(n406), .ZN(n423) );
  NOR2_X1 U383 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U384 ( .A(n425), .B(KEYINPUT35), .ZN(n747) );
  NOR2_X1 U385 ( .A1(n540), .A2(n538), .ZN(n539) );
  NOR2_X1 U386 ( .A1(n697), .A2(n387), .ZN(n379) );
  XNOR2_X1 U387 ( .A(n380), .B(n570), .ZN(n697) );
  XNOR2_X1 U388 ( .A(n578), .B(n351), .ZN(n599) );
  XNOR2_X1 U389 ( .A(n488), .B(n487), .ZN(n581) );
  XNOR2_X1 U390 ( .A(n518), .B(n349), .ZN(n528) );
  XNOR2_X1 U391 ( .A(n384), .B(n481), .ZN(n710) );
  XNOR2_X1 U392 ( .A(n480), .B(n482), .ZN(n384) );
  XNOR2_X1 U393 ( .A(n502), .B(n501), .ZN(n402) );
  XNOR2_X1 U394 ( .A(n497), .B(G134), .ZN(n366) );
  XNOR2_X1 U395 ( .A(n732), .B(G101), .ZN(n382) );
  XNOR2_X1 U396 ( .A(KEYINPUT16), .B(G122), .ZN(n501) );
  XNOR2_X2 U397 ( .A(n423), .B(n611), .ZN(n345) );
  AND2_X2 U398 ( .A1(n714), .A2(n734), .ZN(n354) );
  XNOR2_X2 U399 ( .A(n609), .B(KEYINPUT45), .ZN(n714) );
  XNOR2_X2 U400 ( .A(n447), .B(G128), .ZN(n497) );
  XOR2_X1 U401 ( .A(G131), .B(G140), .Z(n515) );
  INV_X1 U402 ( .A(G237), .ZN(n446) );
  NAND2_X1 U403 ( .A1(n393), .A2(n392), .ZN(n684) );
  AND2_X1 U404 ( .A1(n395), .A2(n394), .ZN(n393) );
  NOR2_X1 U405 ( .A1(n528), .A2(KEYINPUT103), .ZN(n396) );
  XNOR2_X1 U406 ( .A(n381), .B(n483), .ZN(n489) );
  NAND2_X1 U407 ( .A1(n681), .A2(n441), .ZN(n378) );
  XNOR2_X1 U408 ( .A(KEYINPUT15), .B(G902), .ZN(n610) );
  XNOR2_X1 U409 ( .A(n499), .B(KEYINPUT10), .ZN(n514) );
  XNOR2_X1 U410 ( .A(n386), .B(n385), .ZN(n521) );
  INV_X1 U411 ( .A(KEYINPUT8), .ZN(n385) );
  NAND2_X1 U412 ( .A1(n494), .A2(G234), .ZN(n386) );
  XNOR2_X1 U413 ( .A(n364), .B(n513), .ZN(n363) );
  XNOR2_X1 U414 ( .A(G122), .B(G104), .ZN(n513) );
  XNOR2_X1 U415 ( .A(n512), .B(n511), .ZN(n362) );
  XNOR2_X1 U416 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n512) );
  XNOR2_X1 U417 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n359) );
  XNOR2_X1 U418 ( .A(G113), .B(G143), .ZN(n360) );
  NOR2_X1 U419 ( .A1(n747), .A2(n587), .ZN(n430) );
  XNOR2_X1 U420 ( .A(n457), .B(n368), .ZN(n377) );
  INV_X1 U421 ( .A(KEYINPUT30), .ZN(n368) );
  INV_X1 U422 ( .A(G478), .ZN(n398) );
  NOR2_X1 U423 ( .A1(n526), .A2(n389), .ZN(n388) );
  NAND2_X1 U424 ( .A1(n435), .A2(n436), .ZN(n434) );
  XNOR2_X1 U425 ( .A(G116), .B(G113), .ZN(n450) );
  INV_X1 U426 ( .A(KEYINPUT3), .ZN(n449) );
  XNOR2_X1 U427 ( .A(G122), .B(KEYINPUT9), .ZN(n519) );
  XOR2_X1 U428 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n520) );
  XNOR2_X1 U429 ( .A(n470), .B(n469), .ZN(n620) );
  XNOR2_X1 U430 ( .A(n515), .B(n466), .ZN(n468) );
  XNOR2_X1 U431 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U432 ( .A1(n528), .A2(KEYINPUT103), .ZN(n394) );
  NAND2_X1 U433 ( .A1(n537), .A2(KEYINPUT103), .ZN(n395) );
  INV_X1 U434 ( .A(G902), .ZN(n471) );
  INV_X1 U435 ( .A(KEYINPUT90), .ZN(n464) );
  OR2_X1 U436 ( .A1(n610), .A2(KEYINPUT2), .ZN(n422) );
  NAND2_X1 U437 ( .A1(n610), .A2(KEYINPUT80), .ZN(n421) );
  NAND2_X1 U438 ( .A1(n420), .A2(KEYINPUT2), .ZN(n419) );
  NAND2_X1 U439 ( .A1(G234), .A2(G237), .ZN(n458) );
  NOR2_X1 U440 ( .A1(n710), .A2(G902), .ZN(n488) );
  XNOR2_X1 U441 ( .A(n470), .B(n442), .ZN(n612) );
  XNOR2_X1 U442 ( .A(n453), .B(n347), .ZN(n442) );
  XNOR2_X1 U443 ( .A(G110), .B(KEYINPUT23), .ZN(n476) );
  XNOR2_X1 U444 ( .A(n514), .B(n479), .ZN(n480) );
  XNOR2_X1 U445 ( .A(KEYINPUT79), .B(KEYINPUT91), .ZN(n479) );
  XOR2_X1 U446 ( .A(G140), .B(G128), .Z(n475) );
  XNOR2_X1 U447 ( .A(n361), .B(n358), .ZN(n516) );
  XNOR2_X1 U448 ( .A(n360), .B(n359), .ZN(n358) );
  XNOR2_X1 U449 ( .A(n363), .B(n362), .ZN(n361) );
  XNOR2_X1 U450 ( .A(n497), .B(n496), .ZN(n404) );
  XNOR2_X1 U451 ( .A(n530), .B(n529), .ZN(n696) );
  AND2_X1 U452 ( .A1(n681), .A2(n685), .ZN(n365) );
  NAND2_X1 U453 ( .A1(n372), .A2(n369), .ZN(n568) );
  NAND2_X1 U454 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X1 U455 ( .A1(n433), .A2(n432), .ZN(n588) );
  OR2_X1 U456 ( .A1(n528), .A2(n397), .ZN(n649) );
  AND2_X1 U457 ( .A1(n413), .A2(n603), .ZN(n412) );
  NAND2_X1 U458 ( .A1(n674), .A2(n414), .ZN(n413) );
  INV_X1 U459 ( .A(KEYINPUT65), .ZN(n414) );
  BUF_X1 U460 ( .A(n345), .Z(n709) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n705) );
  XNOR2_X1 U462 ( .A(n401), .B(n523), .ZN(n400) );
  XOR2_X1 U463 ( .A(G107), .B(G116), .Z(n522) );
  XNOR2_X1 U464 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U465 ( .A(n390), .B(KEYINPUT42), .ZN(n749) );
  NOR2_X1 U466 ( .A1(n696), .A2(n536), .ZN(n390) );
  INV_X1 U467 ( .A(n579), .ZN(n426) );
  XNOR2_X1 U468 ( .A(n524), .B(n398), .ZN(n537) );
  INV_X1 U469 ( .A(n537), .ZN(n397) );
  INV_X1 U470 ( .A(KEYINPUT2), .ZN(n424) );
  XOR2_X1 U471 ( .A(n507), .B(n506), .Z(n346) );
  XOR2_X1 U472 ( .A(n448), .B(KEYINPUT75), .Z(n347) );
  XOR2_X1 U473 ( .A(n477), .B(n476), .Z(n348) );
  INV_X1 U474 ( .A(n671), .ZN(n389) );
  INV_X1 U475 ( .A(n559), .ZN(n668) );
  XOR2_X1 U476 ( .A(n517), .B(G475), .Z(n349) );
  NAND2_X1 U477 ( .A1(n581), .A2(n671), .ZN(n669) );
  XNOR2_X1 U478 ( .A(n580), .B(KEYINPUT22), .ZN(n350) );
  XOR2_X1 U479 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n351) );
  AND2_X1 U480 ( .A1(n684), .A2(n681), .ZN(n352) );
  XOR2_X1 U481 ( .A(n628), .B(n627), .Z(n353) );
  AND2_X1 U482 ( .A1(n492), .A2(n559), .ZN(n591) );
  BUF_X1 U483 ( .A(n637), .Z(n355) );
  XNOR2_X1 U484 ( .A(n403), .B(n723), .ZN(n637) );
  XNOR2_X1 U485 ( .A(n405), .B(n404), .ZN(n403) );
  XNOR2_X1 U486 ( .A(n500), .B(n382), .ZN(n405) );
  BUF_X1 U487 ( .A(n599), .Z(n387) );
  NAND2_X2 U488 ( .A1(n357), .A2(n356), .ZN(n606) );
  NAND2_X1 U489 ( .A1(n431), .A2(n438), .ZN(n356) );
  NAND2_X1 U490 ( .A1(n434), .A2(n668), .ZN(n357) );
  NOR2_X1 U491 ( .A1(n599), .A2(n350), .ZN(n438) );
  NAND2_X1 U492 ( .A1(n510), .A2(G214), .ZN(n364) );
  NAND2_X1 U493 ( .A1(n537), .A2(n528), .ZN(n579) );
  NAND2_X1 U494 ( .A1(n365), .A2(n684), .ZN(n530) );
  NOR2_X1 U495 ( .A1(n688), .A2(n352), .ZN(n689) );
  XNOR2_X1 U496 ( .A(n366), .B(n522), .ZN(n399) );
  AND2_X1 U497 ( .A1(n493), .A2(n377), .ZN(n371) );
  XNOR2_X2 U498 ( .A(n597), .B(KEYINPUT106), .ZN(n493) );
  INV_X1 U499 ( .A(n377), .ZN(n463) );
  NAND2_X1 U500 ( .A1(n377), .A2(n367), .ZN(n376) );
  INV_X1 U501 ( .A(n378), .ZN(n367) );
  NOR2_X1 U502 ( .A1(n378), .A2(n509), .ZN(n370) );
  INV_X1 U503 ( .A(n509), .ZN(n374) );
  NAND2_X1 U504 ( .A1(n376), .A2(n509), .ZN(n375) );
  XNOR2_X1 U505 ( .A(n379), .B(KEYINPUT34), .ZN(n427) );
  NAND2_X1 U506 ( .A1(n591), .A2(n604), .ZN(n380) );
  NAND2_X1 U507 ( .A1(n489), .A2(G217), .ZN(n484) );
  NAND2_X1 U508 ( .A1(n610), .A2(G234), .ZN(n381) );
  XNOR2_X1 U509 ( .A(n382), .B(G146), .ZN(n418) );
  INV_X2 U510 ( .A(n563), .ZN(n543) );
  XNOR2_X2 U511 ( .A(n383), .B(KEYINPUT105), .ZN(n635) );
  NOR2_X2 U512 ( .A1(n411), .A2(n410), .ZN(n383) );
  NAND2_X1 U513 ( .A1(n427), .A2(n426), .ZN(n425) );
  XNOR2_X2 U514 ( .A(n543), .B(KEYINPUT38), .ZN(n681) );
  AND2_X2 U515 ( .A1(n492), .A2(n547), .ZN(n597) );
  NAND2_X1 U516 ( .A1(n415), .A2(n412), .ZN(n411) );
  NAND2_X1 U517 ( .A1(n396), .A2(n397), .ZN(n392) );
  NAND2_X1 U518 ( .A1(n409), .A2(n419), .ZN(n408) );
  XNOR2_X1 U519 ( .A(n391), .B(n525), .ZN(n742) );
  XNOR2_X1 U520 ( .A(n478), .B(n348), .ZN(n481) );
  NAND2_X1 U521 ( .A1(n603), .A2(n388), .ZN(n548) );
  NOR2_X2 U522 ( .A1(n742), .A2(n749), .ZN(n531) );
  NAND2_X1 U523 ( .A1(n521), .A2(G217), .ZN(n401) );
  XNOR2_X2 U524 ( .A(n467), .B(G104), .ZN(n502) );
  NAND2_X1 U525 ( .A1(n714), .A2(n734), .ZN(n409) );
  NAND2_X1 U526 ( .A1(n354), .A2(n422), .ZN(n406) );
  NOR2_X1 U527 ( .A1(n417), .A2(KEYINPUT65), .ZN(n410) );
  NAND2_X1 U528 ( .A1(n417), .A2(n416), .ZN(n415) );
  AND2_X1 U529 ( .A1(n596), .A2(KEYINPUT65), .ZN(n416) );
  XNOR2_X2 U530 ( .A(n728), .B(n418), .ZN(n470) );
  OR2_X1 U531 ( .A1(n610), .A2(KEYINPUT80), .ZN(n420) );
  XNOR2_X1 U532 ( .A(n354), .B(n424), .ZN(n702) );
  XNOR2_X2 U533 ( .A(n547), .B(KEYINPUT1), .ZN(n559) );
  XNOR2_X2 U534 ( .A(n473), .B(n472), .ZN(n547) );
  NAND2_X1 U535 ( .A1(n428), .A2(n608), .ZN(n609) );
  XNOR2_X1 U536 ( .A(n429), .B(n590), .ZN(n428) );
  NAND2_X1 U537 ( .A1(n635), .A2(n430), .ZN(n429) );
  INV_X1 U538 ( .A(n439), .ZN(n437) );
  NOR2_X1 U539 ( .A1(n439), .A2(n559), .ZN(n431) );
  NAND2_X1 U540 ( .A1(n438), .A2(n437), .ZN(n432) );
  INV_X1 U541 ( .A(n434), .ZN(n433) );
  NAND2_X1 U542 ( .A1(n599), .A2(n350), .ZN(n435) );
  NAND2_X1 U543 ( .A1(n439), .A2(n350), .ZN(n436) );
  NAND2_X1 U544 ( .A1(n684), .A2(n671), .ZN(n439) );
  NOR2_X1 U545 ( .A1(n463), .A2(n440), .ZN(n545) );
  NAND2_X1 U546 ( .A1(n493), .A2(n441), .ZN(n440) );
  INV_X1 U547 ( .A(n526), .ZN(n441) );
  XNOR2_X2 U548 ( .A(G110), .B(G107), .ZN(n467) );
  AND2_X1 U549 ( .A1(n542), .A2(n541), .ZN(n443) );
  XNOR2_X1 U550 ( .A(KEYINPUT62), .B(n612), .ZN(n444) );
  XNOR2_X1 U551 ( .A(n527), .B(KEYINPUT28), .ZN(n445) );
  AND2_X1 U552 ( .A1(n443), .A2(n554), .ZN(n555) );
  INV_X1 U553 ( .A(KEYINPUT48), .ZN(n557) );
  INV_X1 U554 ( .A(n674), .ZN(n596) );
  INV_X1 U555 ( .A(n713), .ZN(n615) );
  NAND2_X1 U556 ( .A1(n471), .A2(n446), .ZN(n504) );
  NAND2_X1 U557 ( .A1(n504), .A2(G214), .ZN(n685) );
  XNOR2_X2 U558 ( .A(KEYINPUT4), .B(KEYINPUT69), .ZN(n732) );
  XNOR2_X1 U559 ( .A(G131), .B(KEYINPUT5), .ZN(n448) );
  XNOR2_X1 U560 ( .A(n449), .B(G119), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n451), .B(n450), .ZN(n503) );
  NAND2_X1 U562 ( .A1(n510), .A2(G210), .ZN(n452) );
  XNOR2_X1 U563 ( .A(n503), .B(n452), .ZN(n453) );
  NAND2_X1 U564 ( .A1(n612), .A2(n471), .ZN(n456) );
  INV_X1 U565 ( .A(KEYINPUT94), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n454), .B(G472), .ZN(n455) );
  XNOR2_X2 U567 ( .A(n456), .B(n455), .ZN(n549) );
  NAND2_X1 U568 ( .A1(n685), .A2(n589), .ZN(n457) );
  XNOR2_X1 U569 ( .A(n458), .B(KEYINPUT14), .ZN(n459) );
  XNOR2_X1 U570 ( .A(KEYINPUT74), .B(n459), .ZN(n460) );
  NAND2_X1 U571 ( .A1(G952), .A2(n460), .ZN(n695) );
  NOR2_X1 U572 ( .A1(G953), .A2(n695), .ZN(n574) );
  NAND2_X1 U573 ( .A1(n460), .A2(G902), .ZN(n572) );
  OR2_X1 U574 ( .A1(n494), .A2(n572), .ZN(n461) );
  NOR2_X1 U575 ( .A1(G900), .A2(n461), .ZN(n462) );
  NOR2_X1 U576 ( .A1(n574), .A2(n462), .ZN(n526) );
  NAND2_X1 U577 ( .A1(G227), .A2(n494), .ZN(n465) );
  XNOR2_X1 U578 ( .A(n468), .B(n502), .ZN(n469) );
  NAND2_X1 U579 ( .A1(n620), .A2(n471), .ZN(n473) );
  XNOR2_X1 U580 ( .A(KEYINPUT70), .B(G469), .ZN(n472) );
  XNOR2_X1 U581 ( .A(G119), .B(G137), .ZN(n474) );
  XNOR2_X1 U582 ( .A(n475), .B(n474), .ZN(n482) );
  NAND2_X1 U583 ( .A1(G221), .A2(n521), .ZN(n478) );
  XOR2_X1 U584 ( .A(KEYINPUT24), .B(KEYINPUT71), .Z(n477) );
  XNOR2_X2 U585 ( .A(G146), .B(G125), .ZN(n499) );
  XOR2_X1 U586 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n485) );
  XOR2_X1 U587 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n483) );
  XNOR2_X1 U588 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U589 ( .A(n486), .B(KEYINPUT92), .ZN(n487) );
  NAND2_X1 U590 ( .A1(n489), .A2(G221), .ZN(n491) );
  INV_X1 U591 ( .A(KEYINPUT21), .ZN(n490) );
  XNOR2_X1 U592 ( .A(n491), .B(n490), .ZN(n671) );
  INV_X1 U593 ( .A(n669), .ZN(n492) );
  NAND2_X1 U594 ( .A1(n494), .A2(G224), .ZN(n495) );
  XNOR2_X1 U595 ( .A(n495), .B(KEYINPUT84), .ZN(n496) );
  XNOR2_X1 U596 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n498) );
  XNOR2_X1 U597 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U598 ( .A1(n637), .A2(n610), .ZN(n508) );
  NAND2_X1 U599 ( .A1(n504), .A2(G210), .ZN(n507) );
  INV_X1 U600 ( .A(KEYINPUT86), .ZN(n505) );
  XNOR2_X1 U601 ( .A(n505), .B(KEYINPUT87), .ZN(n506) );
  XNOR2_X2 U602 ( .A(n508), .B(n346), .ZN(n532) );
  XOR2_X1 U603 ( .A(KEYINPUT72), .B(KEYINPUT39), .Z(n509) );
  INV_X1 U604 ( .A(KEYINPUT100), .ZN(n511) );
  XNOR2_X1 U605 ( .A(n515), .B(n514), .ZN(n729) );
  XNOR2_X1 U606 ( .A(n516), .B(n729), .ZN(n628) );
  NOR2_X1 U607 ( .A1(G902), .A2(n628), .ZN(n518) );
  INV_X1 U608 ( .A(KEYINPUT13), .ZN(n517) );
  XNOR2_X1 U609 ( .A(n520), .B(n519), .ZN(n523) );
  NOR2_X1 U610 ( .A1(G902), .A2(n705), .ZN(n524) );
  NAND2_X1 U611 ( .A1(n528), .A2(n397), .ZN(n645) );
  XNOR2_X1 U612 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n525) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n527) );
  NAND2_X1 U614 ( .A1(n445), .A2(n547), .ZN(n536) );
  XNOR2_X1 U615 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n529) );
  XNOR2_X1 U616 ( .A(n531), .B(KEYINPUT46), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n532), .A2(n685), .ZN(n551) );
  INV_X1 U618 ( .A(KEYINPUT76), .ZN(n533) );
  XNOR2_X1 U619 ( .A(n533), .B(KEYINPUT19), .ZN(n534) );
  XNOR2_X1 U620 ( .A(n551), .B(n534), .ZN(n577) );
  BUF_X1 U621 ( .A(n577), .Z(n535) );
  NOR2_X2 U622 ( .A1(n536), .A2(n535), .ZN(n657) );
  NAND2_X1 U623 ( .A1(n649), .A2(n645), .ZN(n682) );
  NAND2_X1 U624 ( .A1(n657), .A2(n682), .ZN(n540) );
  XNOR2_X1 U625 ( .A(KEYINPUT47), .B(KEYINPUT68), .ZN(n538) );
  XNOR2_X1 U626 ( .A(n539), .B(KEYINPUT73), .ZN(n542) );
  NAND2_X1 U627 ( .A1(n540), .A2(KEYINPUT47), .ZN(n541) );
  NOR2_X1 U628 ( .A1(n579), .A2(n543), .ZN(n544) );
  NAND2_X1 U629 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U630 ( .A(KEYINPUT107), .B(n546), .ZN(n744) );
  XNOR2_X1 U631 ( .A(n559), .B(KEYINPUT85), .ZN(n583) );
  NOR2_X1 U632 ( .A1(n548), .A2(n645), .ZN(n550) );
  XNOR2_X1 U633 ( .A(n549), .B(KEYINPUT6), .ZN(n604) );
  NAND2_X1 U634 ( .A1(n550), .A2(n604), .ZN(n561) );
  NOR2_X1 U635 ( .A1(n561), .A2(n551), .ZN(n552) );
  XOR2_X1 U636 ( .A(KEYINPUT36), .B(n552), .Z(n553) );
  NOR2_X1 U637 ( .A1(n583), .A2(n553), .ZN(n664) );
  NOR2_X1 U638 ( .A1(n744), .A2(n664), .ZN(n554) );
  NAND2_X1 U639 ( .A1(n556), .A2(n555), .ZN(n558) );
  XNOR2_X1 U640 ( .A(n558), .B(n557), .ZN(n566) );
  NAND2_X1 U641 ( .A1(n685), .A2(n668), .ZN(n560) );
  NOR2_X1 U642 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U643 ( .A(n562), .B(KEYINPUT43), .ZN(n564) );
  NOR2_X1 U644 ( .A1(n564), .A2(n563), .ZN(n626) );
  INV_X1 U645 ( .A(n626), .ZN(n565) );
  NAND2_X1 U646 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U647 ( .A(n567), .B(KEYINPUT81), .ZN(n569) );
  OR2_X1 U648 ( .A1(n568), .A2(n649), .ZN(n666) );
  AND2_X2 U649 ( .A1(n569), .A2(n666), .ZN(n734) );
  XNOR2_X1 U650 ( .A(KEYINPUT83), .B(KEYINPUT33), .ZN(n570) );
  NOR2_X1 U651 ( .A1(G898), .A2(n494), .ZN(n571) );
  XOR2_X1 U652 ( .A(KEYINPUT88), .B(n571), .Z(n725) );
  NOR2_X1 U653 ( .A1(n725), .A2(n572), .ZN(n573) );
  OR2_X1 U654 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U655 ( .A(n575), .B(KEYINPUT89), .ZN(n576) );
  INV_X1 U656 ( .A(KEYINPUT66), .ZN(n580) );
  OR2_X1 U657 ( .A1(n604), .A2(n581), .ZN(n582) );
  NOR2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n588), .A2(n584), .ZN(n586) );
  XNOR2_X1 U660 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n585) );
  XNOR2_X1 U661 ( .A(n586), .B(n585), .ZN(n746) );
  INV_X1 U662 ( .A(n746), .ZN(n587) );
  BUF_X1 U663 ( .A(n589), .Z(n674) );
  INV_X1 U664 ( .A(n581), .ZN(n603) );
  INV_X1 U665 ( .A(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n674), .A2(n591), .ZN(n592) );
  XOR2_X1 U667 ( .A(KEYINPUT95), .B(n592), .Z(n677) );
  NOR2_X1 U668 ( .A1(n677), .A2(n387), .ZN(n595) );
  XNOR2_X1 U669 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n593) );
  XNOR2_X1 U670 ( .A(n593), .B(KEYINPUT96), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n595), .B(n594), .ZN(n662) );
  INV_X1 U672 ( .A(n662), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n598) );
  OR2_X1 U674 ( .A1(n387), .A2(n598), .ZN(n644) );
  NAND2_X1 U675 ( .A1(n600), .A2(n644), .ZN(n601) );
  NAND2_X1 U676 ( .A1(n601), .A2(n682), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT102), .ZN(n607) );
  NOR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n642) );
  AND2_X1 U680 ( .A1(n607), .A2(n642), .ZN(n608) );
  INV_X1 U681 ( .A(KEYINPUT64), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n345), .A2(G472), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(n444), .ZN(n616) );
  INV_X1 U684 ( .A(G952), .ZN(n614) );
  AND2_X1 U685 ( .A1(n614), .A2(G953), .ZN(n713) );
  INV_X1 U686 ( .A(KEYINPUT63), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n618), .B(n617), .ZN(G57) );
  NAND2_X1 U688 ( .A1(n704), .A2(G469), .ZN(n622) );
  XNOR2_X1 U689 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n619) );
  XNOR2_X1 U690 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X2 U691 ( .A1(n623), .A2(n713), .ZN(n625) );
  INV_X1 U692 ( .A(KEYINPUT117), .ZN(n624) );
  XNOR2_X1 U693 ( .A(n625), .B(n624), .ZN(G54) );
  XOR2_X1 U694 ( .A(G140), .B(n626), .Z(G42) );
  NAND2_X1 U695 ( .A1(n345), .A2(G475), .ZN(n629) );
  XOR2_X1 U696 ( .A(KEYINPUT118), .B(KEYINPUT59), .Z(n627) );
  XNOR2_X1 U697 ( .A(n629), .B(n353), .ZN(n630) );
  XNOR2_X1 U698 ( .A(KEYINPUT119), .B(KEYINPUT60), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n631), .B(KEYINPUT67), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n633), .B(n632), .ZN(G60) );
  XNOR2_X1 U701 ( .A(G110), .B(KEYINPUT114), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n635), .B(n634), .ZN(G12) );
  NAND2_X1 U703 ( .A1(n704), .A2(G210), .ZN(n639) );
  XNOR2_X1 U704 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n355), .B(n636), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X2 U707 ( .A1(n640), .A2(n713), .ZN(n641) );
  XNOR2_X1 U708 ( .A(n641), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U709 ( .A(G101), .B(KEYINPUT110), .ZN(n643) );
  XNOR2_X1 U710 ( .A(n643), .B(n642), .ZN(G3) );
  INV_X1 U711 ( .A(n644), .ZN(n650) );
  INV_X1 U712 ( .A(n645), .ZN(n659) );
  NAND2_X1 U713 ( .A1(n650), .A2(n659), .ZN(n646) );
  XNOR2_X1 U714 ( .A(n646), .B(G104), .ZN(G6) );
  XOR2_X1 U715 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n648) );
  XNOR2_X1 U716 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n654) );
  XNOR2_X1 U718 ( .A(G107), .B(KEYINPUT26), .ZN(n652) );
  INV_X1 U719 ( .A(n649), .ZN(n661) );
  NAND2_X1 U720 ( .A1(n661), .A2(n650), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(G9) );
  XOR2_X1 U723 ( .A(G128), .B(KEYINPUT29), .Z(n656) );
  NAND2_X1 U724 ( .A1(n657), .A2(n661), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n656), .B(n655), .ZN(G30) );
  NAND2_X1 U726 ( .A1(n657), .A2(n659), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n658), .B(G146), .ZN(G48) );
  NAND2_X1 U728 ( .A1(n659), .A2(n662), .ZN(n660) );
  XNOR2_X1 U729 ( .A(G113), .B(n660), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(G116), .ZN(G18) );
  XNOR2_X1 U732 ( .A(G125), .B(n664), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U734 ( .A(n666), .ZN(n667) );
  XOR2_X1 U735 ( .A(G134), .B(n667), .Z(G36) );
  XOR2_X1 U736 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n693) );
  NAND2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n670), .B(KEYINPUT50), .ZN(n676) );
  NOR2_X1 U739 ( .A1(n671), .A2(n581), .ZN(n672) );
  XOR2_X1 U740 ( .A(KEYINPUT49), .B(n672), .Z(n673) );
  NOR2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U744 ( .A(KEYINPUT51), .B(n679), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n696), .A2(n680), .ZN(n691) );
  AND2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n687) );
  INV_X1 U748 ( .A(n685), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n697), .A2(n689), .ZN(n690) );
  NOR2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U752 ( .A(n693), .B(n692), .Z(n694) );
  NOR2_X1 U753 ( .A1(n695), .A2(n694), .ZN(n699) );
  NOR2_X1 U754 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U755 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U756 ( .A1(n700), .A2(n494), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U758 ( .A(n703), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U759 ( .A1(n709), .A2(G478), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n705), .B(KEYINPUT120), .ZN(n706) );
  XNOR2_X1 U761 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n713), .A2(n708), .ZN(G63) );
  NAND2_X1 U763 ( .A1(n709), .A2(G217), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n710), .B(n711), .ZN(n712) );
  NOR2_X1 U765 ( .A1(n713), .A2(n712), .ZN(G66) );
  BUF_X1 U766 ( .A(n714), .Z(n715) );
  NAND2_X1 U767 ( .A1(n715), .A2(n494), .ZN(n721) );
  XOR2_X1 U768 ( .A(KEYINPUT61), .B(KEYINPUT122), .Z(n717) );
  NAND2_X1 U769 ( .A1(G224), .A2(G953), .ZN(n716) );
  XNOR2_X1 U770 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U771 ( .A(KEYINPUT121), .B(n718), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n719), .A2(G898), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n727) );
  XOR2_X1 U774 ( .A(G101), .B(KEYINPUT123), .Z(n722) );
  XNOR2_X1 U775 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U777 ( .A(n727), .B(n726), .Z(G69) );
  XNOR2_X1 U778 ( .A(n728), .B(KEYINPUT124), .ZN(n730) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U780 ( .A(n732), .B(n731), .ZN(n737) );
  INV_X1 U781 ( .A(n737), .ZN(n733) );
  XOR2_X1 U782 ( .A(n734), .B(n733), .Z(n735) );
  NOR2_X1 U783 ( .A1(G953), .A2(n735), .ZN(n736) );
  XNOR2_X1 U784 ( .A(KEYINPUT125), .B(n736), .ZN(n741) );
  XNOR2_X1 U785 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(G72) );
  BUF_X1 U789 ( .A(n742), .Z(n743) );
  XOR2_X1 U790 ( .A(n743), .B(G131), .Z(G33) );
  XNOR2_X1 U791 ( .A(G143), .B(n744), .ZN(n745) );
  XNOR2_X1 U792 ( .A(n745), .B(KEYINPUT115), .ZN(G45) );
  XNOR2_X1 U793 ( .A(G119), .B(n746), .ZN(G21) );
  XOR2_X1 U794 ( .A(G122), .B(n747), .Z(n748) );
  XNOR2_X1 U795 ( .A(KEYINPUT126), .B(n748), .ZN(G24) );
  XOR2_X1 U796 ( .A(G137), .B(n749), .Z(G39) );
endmodule

