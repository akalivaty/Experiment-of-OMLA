//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT66), .A2(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT66), .A2(G116), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n191), .A2(KEYINPUT67), .A3(G119), .A4(new_n192), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT66), .A2(G116), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT66), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(G116), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n193), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT2), .B(G113), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n202), .B(new_n193), .C1(new_n197), .C2(new_n200), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n197), .A2(new_n200), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n208), .A2(KEYINPUT68), .A3(new_n202), .A4(new_n193), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT65), .A3(G134), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n212), .B2(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n214), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G143), .B(G146), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G143), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(KEYINPUT64), .A3(G146), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(G143), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n226), .B1(new_n236), .B2(KEYINPUT1), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n228), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n229), .A2(KEYINPUT64), .A3(G146), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT64), .B1(new_n229), .B2(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n236), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n241), .A2(new_n244), .B1(new_n242), .B2(new_n225), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n220), .A2(new_n221), .A3(new_n214), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n223), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n224), .A2(new_n238), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT28), .B1(new_n210), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n210), .A2(new_n249), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n248), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n238), .A2(new_n223), .A3(new_n218), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n209), .A3(new_n207), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n252), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n209), .A4(new_n207), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT28), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n251), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT27), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n255), .A2(new_n268), .A3(KEYINPUT30), .ZN(new_n269));
  OR2_X1    g083(.A1(new_n268), .A2(KEYINPUT30), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(KEYINPUT30), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n253), .A2(new_n254), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n210), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n252), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n274), .A3(new_n267), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n261), .A2(new_n267), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n207), .A2(new_n209), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n271), .B1(new_n249), .B2(new_n270), .ZN(new_n279));
  INV_X1    g093(.A(new_n272), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n252), .A3(new_n266), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT31), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT71), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n281), .A2(new_n276), .A3(new_n252), .A4(new_n266), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n259), .A2(KEYINPUT28), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n252), .A2(new_n256), .A3(new_n257), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n250), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n285), .B1(new_n288), .B2(new_n266), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n273), .A2(new_n274), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n276), .B1(new_n291), .B2(new_n266), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n190), .B1(new_n284), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n267), .B1(new_n273), .B2(new_n274), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n295), .B(new_n296), .C1(new_n261), .C2(new_n267), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n252), .A2(new_n256), .A3(KEYINPUT72), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n210), .A2(new_n299), .A3(new_n249), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(KEYINPUT28), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n267), .A2(new_n295), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n251), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n301), .A2(KEYINPUT73), .A3(new_n251), .A4(new_n302), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n297), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G472), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n290), .B1(new_n289), .B2(new_n292), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n261), .A2(new_n267), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n311), .A2(new_n283), .A3(KEYINPUT71), .A4(new_n285), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n188), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n294), .B(new_n309), .C1(KEYINPUT32), .C2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G137), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(G221), .A3(G234), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n315), .B(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n196), .A2(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n226), .A2(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT74), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT24), .B(G110), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n226), .A2(KEYINPUT23), .A3(G119), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n196), .A2(G128), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n319), .B(new_n328), .C1(new_n329), .C2(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G110), .ZN(new_n331));
  INV_X1    g145(.A(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G125), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n335), .A3(KEYINPUT16), .ZN(new_n336));
  OR3_X1    g150(.A1(new_n334), .A2(KEYINPUT16), .A3(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G146), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(G146), .B1(new_n336), .B2(new_n337), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n327), .B(new_n331), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n337), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n232), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n338), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(KEYINPUT75), .A3(new_n327), .A4(new_n331), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n333), .A2(new_n335), .A3(new_n232), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n338), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n324), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT74), .B1(new_n319), .B2(new_n320), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n325), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n330), .A2(G110), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n318), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n318), .ZN(new_n358));
  AOI211_X1 g172(.A(new_n358), .B(new_n355), .C1(new_n343), .C2(new_n347), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G217), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(G234), .B2(new_n306), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT77), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n357), .A2(new_n359), .A3(G902), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n348), .A2(new_n356), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n358), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n355), .B1(new_n343), .B2(new_n347), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n318), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n306), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(new_n375), .A3(new_n362), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n365), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT9), .B(G234), .ZN(new_n379));
  OAI21_X1  g193(.A(G221), .B1(new_n379), .B2(G902), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n316), .A2(G227), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G104), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT79), .B1(new_n388), .B2(G107), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n386), .A2(G104), .ZN(new_n390));
  OAI211_X1 g204(.A(G101), .B(new_n387), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(new_n388), .B2(G107), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n386), .A3(G104), .ZN(new_n394));
  INV_X1    g208(.A(G101), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n388), .A2(G107), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n392), .A2(new_n394), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT1), .B1(new_n229), .B2(G146), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n229), .A2(G146), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n399), .A2(G128), .B1(new_n236), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n228), .B1(new_n401), .B2(KEYINPUT80), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n237), .A2(new_n225), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n398), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT10), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n248), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n392), .A2(new_n394), .A3(new_n396), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n395), .A2(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n412), .B2(new_n397), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT4), .B1(new_n410), .B2(new_n411), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n245), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n398), .A2(KEYINPUT10), .A3(new_n238), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n407), .A2(new_n408), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n227), .A2(new_n236), .A3(new_n400), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n399), .A2(G128), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n241), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n391), .A2(new_n397), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n405), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT12), .B1(new_n423), .B2(new_n248), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n425), .B(new_n408), .C1(new_n405), .C2(new_n422), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n417), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT81), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n429), .B(new_n417), .C1(new_n424), .C2(new_n426), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n384), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G469), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n415), .A2(new_n416), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n408), .B1(new_n433), .B2(new_n407), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n417), .A2(new_n384), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n431), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n424), .A2(new_n426), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(new_n435), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n415), .A2(new_n416), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n236), .A2(new_n400), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n419), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n418), .B1(new_n442), .B2(new_n403), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n401), .A2(KEYINPUT80), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n421), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(KEYINPUT10), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n248), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n384), .B1(new_n447), .B2(new_n417), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n432), .B(new_n306), .C1(new_n439), .C2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n432), .A2(new_n306), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n380), .B1(new_n437), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G214), .B1(G237), .B2(G902), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n201), .A2(KEYINPUT5), .ZN(new_n455));
  OAI21_X1  g269(.A(G113), .B1(new_n198), .B2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n204), .A3(new_n398), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n413), .A2(new_n414), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n459), .B(new_n460), .C1(new_n210), .C2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n245), .A2(new_n334), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT82), .B1(new_n245), .B2(new_n334), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n420), .A2(new_n334), .ZN(new_n467));
  INV_X1    g281(.A(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n465), .A2(new_n466), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n467), .ZN(new_n473));
  OAI22_X1  g287(.A1(new_n473), .A2(new_n463), .B1(new_n470), .B2(new_n469), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n462), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT83), .B(KEYINPUT8), .Z(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(new_n460), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n204), .A2(new_n398), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n455), .A2(KEYINPUT84), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n456), .B1(new_n455), .B2(KEYINPUT84), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n398), .B1(new_n458), .B2(new_n204), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n475), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n459), .B1(new_n210), .B2(new_n461), .ZN(new_n485));
  INV_X1    g299(.A(new_n460), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT6), .A3(new_n462), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n469), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n491), .A3(new_n486), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n484), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n484), .B2(new_n493), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n454), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n453), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G237), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n316), .A3(G214), .ZN(new_n500));
  AND2_X1   g314(.A1(KEYINPUT85), .A2(G143), .ZN(new_n501));
  NOR2_X1   g315(.A1(KEYINPUT85), .A2(G143), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n262), .B(G214), .C1(KEYINPUT85), .C2(G143), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G131), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT89), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n222), .A3(new_n504), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n510), .A3(G131), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n510), .B1(new_n505), .B2(G131), .ZN(new_n513));
  AOI211_X1 g327(.A(KEYINPUT89), .B(new_n222), .C1(new_n503), .C2(new_n504), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT17), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR3_X1    g329(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT90), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n346), .A2(KEYINPUT90), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n512), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G113), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n388), .ZN(new_n520));
  NAND2_X1  g334(.A1(KEYINPUT18), .A2(G131), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n503), .A2(new_n521), .A3(new_n504), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n333), .A2(new_n335), .A3(new_n232), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n232), .B1(new_n333), .B2(new_n335), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n333), .A2(new_n335), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G146), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n349), .A3(KEYINPUT87), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n521), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT86), .B1(new_n505), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n535), .B(new_n521), .C1(new_n503), .C2(new_n504), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n524), .B(new_n532), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n518), .A2(new_n520), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n508), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n513), .A2(new_n514), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n529), .B(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n338), .B1(new_n541), .B2(G146), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n522), .B(KEYINPUT88), .ZN(new_n544));
  OAI22_X1  g358(.A1(new_n540), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n520), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(G475), .A2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT20), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n538), .A2(new_n547), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n538), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n520), .B1(new_n518), .B2(new_n537), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(KEYINPUT91), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n306), .ZN(new_n561));
  OAI21_X1  g375(.A(G475), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G952), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n564), .A2(KEYINPUT95), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(KEYINPUT95), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n316), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(G234), .B2(G237), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT21), .B(G898), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n306), .B(new_n316), .C1(G234), .C2(G237), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n379), .A2(new_n361), .A3(G953), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n574));
  INV_X1    g388(.A(G116), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(G122), .ZN(new_n576));
  INV_X1    g390(.A(G122), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT92), .A3(G116), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n191), .A2(G122), .A3(new_n192), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n579), .B2(new_n580), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n386), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n580), .A2(KEYINPUT14), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n579), .B1(new_n580), .B2(KEYINPUT14), .ZN(new_n586));
  OAI21_X1  g400(.A(G107), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n229), .A2(G128), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n226), .A2(G143), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G134), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n589), .A3(new_n212), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n584), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT13), .ZN(new_n597));
  OAI21_X1  g411(.A(G134), .B1(new_n588), .B2(KEYINPUT13), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n226), .A2(G143), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT13), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n212), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n602), .B(KEYINPUT94), .C1(new_n601), .C2(new_n590), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n603), .A3(new_n592), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n579), .A2(new_n580), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT93), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(G107), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n584), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n573), .B1(new_n595), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n584), .A2(new_n608), .ZN(new_n611));
  INV_X1    g425(.A(new_n604), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n594), .A3(new_n572), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G478), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n616), .A2(KEYINPUT15), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n563), .A2(new_n571), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n314), .A2(new_n378), .A3(new_n498), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n310), .A2(new_n312), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n306), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n313), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n453), .A2(new_n377), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n571), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n454), .B(new_n630), .C1(new_n495), .C2(new_n496), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n595), .A2(new_n609), .A3(new_n573), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n572), .B1(new_n613), .B2(new_n594), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT33), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n610), .A2(new_n614), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(G478), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n616), .A2(new_n306), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n615), .B2(new_n616), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n563), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n629), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND3_X1  g459(.A1(new_n551), .A2(KEYINPUT96), .A3(new_n554), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n553), .B1(new_n552), .B2(new_n549), .ZN(new_n648));
  AOI211_X1 g462(.A(KEYINPUT20), .B(new_n550), .C1(new_n538), .C2(new_n547), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n562), .A3(new_n620), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n631), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n629), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n370), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n372), .A2(new_n657), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT97), .ZN(new_n662));
  INV_X1    g476(.A(new_n363), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n372), .B(new_n658), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT97), .B1(new_n665), .B2(new_n363), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n376), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n497), .A2(new_n453), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n627), .A2(new_n669), .A3(new_n621), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n568), .B1(new_n673), .B2(new_n570), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n652), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n314), .A2(new_n669), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  INV_X1    g491(.A(new_n380), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n428), .A2(new_n430), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n436), .B1(new_n679), .B2(new_n383), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G469), .ZN(new_n681));
  INV_X1    g495(.A(new_n417), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n383), .B1(new_n434), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n398), .A2(new_n238), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n248), .B1(new_n445), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n425), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n423), .A2(KEYINPUT12), .A3(new_n248), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n384), .A3(new_n417), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n450), .B1(new_n690), .B2(new_n432), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n678), .B1(new_n681), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n674), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT40), .Z(new_n695));
  OAI21_X1  g509(.A(new_n266), .B1(new_n273), .B2(new_n274), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n266), .B1(new_n298), .B2(new_n300), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n697), .A2(G902), .A3(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(new_n624), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n294), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n625), .A2(new_n187), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n189), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n484), .A2(new_n493), .ZN(new_n706));
  INV_X1    g520(.A(new_n494), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n484), .A2(new_n493), .A3(new_n494), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n710), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n648), .A2(new_n649), .ZN(new_n714));
  INV_X1    g528(.A(G475), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n518), .A2(new_n537), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n546), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n556), .A3(new_n538), .ZN(new_n718));
  AOI21_X1  g532(.A(G902), .B1(new_n558), .B2(KEYINPUT91), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n620), .B1(new_n714), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n668), .A3(new_n454), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n713), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n695), .A2(new_n705), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  INV_X1    g540(.A(new_n674), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n640), .B(new_n727), .C1(new_n714), .C2(new_n720), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n314), .A2(new_n669), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  OAI21_X1  g545(.A(new_n306), .B1(new_n439), .B2(new_n448), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n380), .A3(new_n449), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT99), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT99), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n736), .A3(new_n380), .A4(new_n449), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n735), .A2(KEYINPUT100), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT100), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n625), .A2(new_n190), .B1(new_n308), .B2(G472), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n377), .B1(new_n704), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n742), .A3(new_n642), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT41), .B(G113), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G15));
  INV_X1    g559(.A(KEYINPUT101), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n735), .A2(new_n737), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT100), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n735), .A2(KEYINPUT100), .A3(new_n737), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n314), .A2(new_n749), .A3(new_n378), .A4(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n653), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n746), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n740), .A2(new_n742), .A3(KEYINPUT101), .A4(new_n653), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G116), .ZN(G18));
  INV_X1    g570(.A(new_n454), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n708), .B2(new_n709), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n758), .A2(new_n735), .A3(new_n737), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n376), .A2(new_n667), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n314), .A2(new_n759), .A3(new_n621), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G119), .ZN(G21));
  INV_X1    g576(.A(new_n285), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n301), .A2(new_n251), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n764), .A2(new_n267), .B1(new_n282), .B2(KEYINPUT31), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n763), .B1(new_n765), .B2(KEYINPUT102), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT102), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n266), .B1(new_n301), .B2(new_n251), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(new_n292), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n188), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n626), .A2(new_n770), .A3(new_n377), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n758), .A2(new_n722), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n571), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n740), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NAND2_X1  g589(.A1(new_n728), .A2(KEYINPUT103), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT103), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n563), .A2(new_n777), .A3(new_n640), .A4(new_n727), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n306), .B1(new_n284), .B2(new_n293), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n765), .A2(KEYINPUT102), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n285), .A3(new_n769), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n780), .A2(G472), .B1(new_n782), .B2(new_n187), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n779), .A2(new_n783), .A3(new_n759), .A4(new_n760), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  AOI21_X1  g599(.A(new_n429), .B1(new_n688), .B2(new_n417), .ZN(new_n786));
  INV_X1    g600(.A(new_n430), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n383), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT104), .ZN(new_n789));
  INV_X1    g603(.A(new_n436), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n788), .A2(new_n789), .A3(G469), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n691), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n789), .B1(new_n680), .B2(G469), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n380), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n708), .A2(new_n454), .A3(new_n709), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n779), .A3(new_n314), .A4(new_n378), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT42), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n776), .A2(new_n778), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n795), .A3(new_n794), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT105), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n294), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n625), .A2(KEYINPUT105), .A3(new_n190), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n704), .A2(new_n803), .A3(new_n309), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n801), .A2(new_n805), .A3(KEYINPUT42), .A4(new_n378), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G131), .ZN(G33));
  NAND4_X1  g622(.A1(new_n796), .A2(new_n314), .A3(new_n378), .A4(new_n675), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G134), .ZN(G36));
  NOR2_X1   g624(.A1(new_n714), .A2(new_n720), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n640), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT43), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(KEYINPUT43), .A3(new_n640), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n668), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n313), .B2(new_n626), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT44), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT107), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n680), .A2(KEYINPUT45), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT45), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n431), .B2(new_n436), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(G469), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(KEYINPUT46), .A3(new_n451), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT46), .B1(new_n824), .B2(new_n451), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n449), .B(new_n825), .C1(new_n826), .C2(KEYINPUT106), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(KEYINPUT106), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n678), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n795), .B(KEYINPUT108), .Z(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n817), .B2(new_n818), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n820), .A2(new_n693), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G137), .ZN(G39));
  INV_X1    g648(.A(KEYINPUT47), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n829), .B2(new_n678), .ZN(new_n836));
  OAI211_X1 g650(.A(KEYINPUT47), .B(new_n380), .C1(new_n827), .C2(new_n828), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n314), .A2(new_n378), .A3(new_n728), .A4(new_n795), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G140), .ZN(G42));
  NAND2_X1  g655(.A1(new_n564), .A2(new_n316), .ZN(new_n842));
  INV_X1    g656(.A(new_n568), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n814), .B2(new_n815), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n771), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n758), .A2(new_n735), .A3(new_n737), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT117), .Z(new_n848));
  NOR2_X1   g662(.A1(new_n747), .A2(new_n795), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n805), .A2(new_n378), .A3(new_n844), .A4(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT48), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n377), .A2(new_n843), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n702), .A3(new_n704), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n641), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n567), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n848), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n733), .A2(new_n678), .A3(new_n449), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n836), .A2(new_n837), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n845), .A2(new_n831), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n626), .A2(new_n770), .A3(new_n668), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n844), .A3(new_n849), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n563), .A2(new_n640), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n863), .B1(new_n853), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n713), .A2(new_n757), .A3(new_n737), .A4(new_n735), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT116), .B1(new_n866), .B2(new_n845), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  OAI211_X1 g683(.A(KEYINPUT116), .B(new_n869), .C1(new_n866), .C2(new_n845), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n865), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n861), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n861), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n857), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n857), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n376), .A2(new_n667), .A3(new_n727), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n497), .A2(new_n880), .A3(new_n721), .ZN(new_n881));
  INV_X1    g695(.A(new_n793), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n452), .B1(new_n437), .B2(new_n789), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n678), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n313), .A2(KEYINPUT32), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n881), .B(new_n884), .C1(new_n701), .C2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n784), .A2(new_n676), .A3(new_n730), .A4(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT113), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n730), .A2(new_n886), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n692), .A2(new_n758), .A3(new_n760), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n704), .B2(new_n741), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n800), .A2(new_n846), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n892), .A2(new_n675), .B1(new_n893), .B2(new_n862), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT113), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n890), .A2(new_n894), .A3(new_n895), .A4(KEYINPUT52), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g711(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n887), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT115), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT115), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n887), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n642), .A2(KEYINPUT110), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT110), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n631), .B2(new_n641), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n904), .A2(new_n627), .A3(new_n628), .A4(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n743), .A2(new_n774), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n620), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT111), .B1(new_n563), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT111), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n811), .A2(new_n911), .A3(new_n620), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n631), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n627), .A2(new_n913), .A3(new_n628), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n622), .A2(new_n761), .A3(new_n914), .A4(new_n670), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n908), .A2(new_n755), .A3(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n796), .A2(new_n779), .A3(new_n783), .A4(new_n760), .ZN(new_n918));
  INV_X1    g732(.A(new_n795), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n620), .A2(new_n720), .A3(new_n674), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n920), .A2(new_n651), .A3(new_n760), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n314), .A2(new_n692), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n918), .A2(new_n809), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT112), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n918), .A2(new_n809), .A3(KEYINPUT112), .A4(new_n922), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n807), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n917), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT53), .B1(new_n903), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n918), .A2(new_n809), .A3(new_n922), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n930), .A2(KEYINPUT112), .B1(new_n806), .B2(new_n799), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n743), .A2(new_n774), .A3(new_n907), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n915), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n931), .A2(new_n755), .A3(new_n933), .A4(new_n925), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT53), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n887), .B(KEYINPUT52), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT54), .B1(new_n929), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n903), .A2(new_n928), .A3(KEYINPUT53), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n842), .B1(new_n879), .B2(new_n943), .ZN(new_n944));
  NOR4_X1   g758(.A1(new_n812), .A2(new_n377), .A3(new_n757), .A4(new_n678), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n733), .A2(new_n449), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT49), .Z(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n713), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n705), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT109), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n944), .A2(new_n950), .ZN(G75));
  NAND2_X1  g765(.A1(new_n939), .A2(new_n940), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(G210), .A3(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n490), .B(KEYINPUT55), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT120), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n488), .A2(new_n492), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT119), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n955), .B(new_n957), .Z(new_n958));
  XOR2_X1   g772(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n953), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n316), .A2(G952), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT56), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n958), .B1(new_n953), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(G51));
  XNOR2_X1  g780(.A(new_n450), .B(KEYINPUT57), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n941), .B1(new_n939), .B2(new_n940), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n683), .A2(new_n689), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n939), .A2(new_n940), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n973), .A2(new_n306), .A3(new_n824), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n961), .B1(new_n972), .B2(new_n974), .ZN(G54));
  NAND2_X1  g789(.A1(KEYINPUT58), .A2(G475), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT122), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n952), .A2(G902), .A3(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(new_n548), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n548), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n979), .A2(new_n980), .A3(new_n961), .ZN(G60));
  NAND2_X1  g795(.A1(new_n634), .A2(new_n636), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n638), .B(KEYINPUT59), .Z(new_n983));
  OAI211_X1 g797(.A(new_n982), .B(new_n983), .C1(new_n968), .C2(new_n969), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n962), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n982), .B1(new_n943), .B2(new_n983), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n939), .B2(new_n940), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(new_n360), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n665), .ZN(new_n992));
  XNOR2_X1  g806(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n991), .A2(new_n992), .A3(new_n962), .A4(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n962), .B1(new_n990), .B2(new_n360), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n661), .B(new_n989), .C1(new_n939), .C2(new_n940), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n994), .A2(new_n998), .ZN(G66));
  OAI21_X1  g813(.A(G953), .B1(new_n569), .B2(new_n468), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT124), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n917), .B2(new_n316), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT125), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n957), .B1(G898), .B2(new_n316), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  NAND2_X1  g819(.A1(new_n805), .A2(new_n378), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(new_n772), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n830), .A2(new_n693), .A3(new_n1007), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n784), .A2(new_n676), .A3(new_n730), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n807), .A2(new_n809), .A3(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n833), .A2(new_n840), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n269), .A2(new_n272), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT126), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(new_n541), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1014), .A2(new_n316), .ZN(new_n1015));
  AOI22_X1  g829(.A1(new_n1011), .A2(new_n1015), .B1(new_n673), .B2(G953), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n725), .A2(new_n1009), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT62), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n910), .A2(new_n641), .A3(new_n912), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n694), .A2(new_n795), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n742), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1019), .A2(new_n833), .A3(new_n840), .A4(new_n1022), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1023), .A2(new_n316), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1016), .B1(new_n1024), .B2(new_n1014), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1014), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n316), .B1(G227), .B2(G900), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n1016), .B(new_n1030), .C1(new_n1024), .C2(new_n1014), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(new_n1031), .ZN(G72));
  NAND2_X1  g846(.A1(G472), .A2(G902), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n1033), .B(KEYINPUT63), .Z(new_n1034));
  OAI21_X1  g848(.A(new_n1034), .B1(new_n1023), .B2(new_n917), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n961), .B1(new_n1035), .B2(new_n697), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1034), .B1(new_n1011), .B2(new_n917), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n291), .A3(new_n267), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n282), .A2(new_n296), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1034), .B(new_n1039), .C1(new_n929), .C2(new_n937), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n1036), .A2(new_n1038), .A3(new_n1040), .ZN(G57));
endmodule


