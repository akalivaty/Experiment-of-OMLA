//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OR3_X1    g003(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n202), .A2(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT89), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n206), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(new_n205), .B2(new_n210), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n211), .A2(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n209), .B1(new_n214), .B2(new_n204), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT90), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT90), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n209), .B(new_n217), .C1(new_n214), .C2(new_n204), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT91), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G1gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT91), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n221), .B(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G1gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT92), .B(new_n220), .C1(new_n223), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n222), .B1(new_n226), .B2(G1gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G8gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G1gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(G8gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n230), .A2(new_n233), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n238), .A3(KEYINPUT93), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n216), .A2(new_n229), .A3(new_n218), .A4(new_n237), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT93), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n216), .A2(new_n245), .A3(new_n218), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n237), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n215), .A2(new_n245), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n243), .A2(new_n244), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(KEYINPUT94), .A2(KEYINPUT18), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n219), .A2(new_n238), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n243), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n244), .B(KEYINPUT13), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n251), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n243), .A2(new_n244), .A3(new_n249), .A4(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n252), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G113gat), .B(G141gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G197gat), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT11), .B(G169gat), .Z(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n252), .A2(new_n256), .A3(new_n265), .A4(new_n258), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G190gat), .B(G218gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(G232gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT41), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G99gat), .A2(G106gat), .ZN(new_n274));
  INV_X1    g073(.A(G85gat), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  AOI22_X1  g075(.A1(KEYINPUT8), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT98), .ZN(new_n278));
  NAND2_X1  g077(.A1(G85gat), .A2(G92gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT7), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G99gat), .B(G106gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n278), .A2(new_n282), .A3(new_n280), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(KEYINPUT99), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT99), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n281), .A2(new_n287), .A3(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n273), .B1(new_n219), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT100), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n246), .A2(new_n248), .A3(new_n288), .A4(new_n286), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n270), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n295), .ZN(new_n297));
  INV_X1    g096(.A(new_n270), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n271), .A2(new_n272), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT97), .ZN(new_n302));
  XOR2_X1   g101(.A(G134gat), .B(G162gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(KEYINPUT101), .Z(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n304), .A2(KEYINPUT101), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n296), .A2(new_n299), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G183gat), .B(G211gat), .Z(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(G71gat), .A2(G78gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT9), .ZN(new_n314));
  XNOR2_X1  g113(.A(G57gat), .B(G64gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(G71gat), .A2(G78gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n313), .A2(KEYINPUT95), .ZN(new_n319));
  OR3_X1    g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n316), .B2(new_n319), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT21), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G231gat), .A2(G233gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G127gat), .B(G155gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT20), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n329), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n312), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n247), .B1(new_n324), .B2(new_n323), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  NAND3_X1  g136(.A1(new_n331), .A2(new_n312), .A3(new_n332), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n334), .B2(new_n338), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n310), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G230gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n286), .A2(new_n323), .A3(new_n288), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT10), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n284), .A2(new_n322), .A3(new_n285), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n289), .A2(KEYINPUT10), .A3(new_n322), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n347), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G120gat), .B(G148gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G176gat), .B(G204gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  OR2_X1    g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n355), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  XNOR2_X1  g159(.A(G197gat), .B(G204gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(G211gat), .A2(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(KEYINPUT22), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G211gat), .ZN(new_n365));
  INV_X1    g164(.A(G218gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n362), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n364), .B(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n360), .B1(new_n369), .B2(KEYINPUT29), .ZN(new_n370));
  NAND2_X1  g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT76), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(G155gat), .A3(G162gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G155gat), .ZN(new_n376));
  INV_X1    g175(.A(G162gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n371), .A2(KEYINPUT2), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G141gat), .B(G148gat), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n375), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n371), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n378), .A2(KEYINPUT78), .A3(new_n371), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n379), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G141gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(G148gat), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT77), .B(G141gat), .Z(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(G148gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n382), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n370), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n389), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT77), .B(G141gat), .ZN(new_n395));
  INV_X1    g194(.A(G148gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n397), .A2(new_n379), .A3(new_n386), .A4(new_n385), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(new_n360), .A3(new_n382), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n369), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n393), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G228gat), .ZN(new_n406));
  INV_X1    g205(.A(G233gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n368), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n364), .B(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n399), .A2(new_n401), .ZN(new_n412));
  OAI221_X1 g211(.A(new_n393), .B1(new_n406), .B2(new_n407), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n415), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n409), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(G22gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n416), .A2(new_n421), .A3(new_n418), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G120gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G113gat), .ZN(new_n428));
  INV_X1    g227(.A(G113gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(G120gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT1), .ZN(new_n432));
  INV_X1    g231(.A(G134gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G127gat), .ZN(new_n434));
  INV_X1    g233(.A(G127gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G134gat), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n431), .A2(new_n432), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n436), .ZN(new_n438));
  XNOR2_X1  g237(.A(G113gat), .B(G120gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n438), .B1(new_n439), .B2(KEYINPUT1), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT4), .B1(new_n392), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n441), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n443), .A2(new_n398), .A3(new_n444), .A4(new_n382), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n441), .A3(new_n399), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n392), .A2(new_n441), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(new_n398), .A3(new_n382), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n447), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n445), .A2(KEYINPUT79), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n442), .A2(KEYINPUT79), .A3(new_n445), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n455), .A2(KEYINPUT5), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n449), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G1gat), .B(G29gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT0), .ZN(new_n464));
  XNOR2_X1  g263(.A(G57gat), .B(G85gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n464), .B(new_n465), .Z(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n457), .A2(new_n466), .A3(new_n461), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n462), .A2(KEYINPUT6), .A3(new_n467), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475));
  INV_X1    g274(.A(G169gat), .ZN(new_n476));
  INV_X1    g275(.A(G176gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT23), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(G169gat), .B2(G176gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(G169gat), .A2(G176gat), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G183gat), .A2(G190gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT24), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G183gat), .ZN(new_n486));
  INV_X1    g285(.A(G190gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n485), .A2(KEYINPUT65), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT65), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n493), .A2(new_n496), .A3(new_n488), .A4(new_n489), .ZN(new_n497));
  AND4_X1   g296(.A1(KEYINPUT25), .A2(new_n478), .A3(new_n480), .A4(new_n481), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n491), .A2(new_n492), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n483), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n486), .A2(KEYINPUT27), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT27), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G183gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n503), .A3(new_n487), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT28), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n500), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT67), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT26), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT26), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(new_n476), .A3(new_n477), .A4(KEYINPUT67), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n481), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G183gat), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n514), .A2(new_n505), .A3(new_n506), .A4(new_n487), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n508), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n499), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n475), .B1(new_n517), .B2(KEYINPUT29), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n518), .B(new_n411), .C1(new_n517), .C2(new_n475), .ZN(new_n519));
  INV_X1    g318(.A(new_n490), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n492), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n497), .A2(new_n498), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n513), .A3(new_n515), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n526), .A2(new_n401), .B1(G226gat), .B2(G233gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n517), .A2(new_n475), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n369), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G64gat), .B(G92gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  NAND3_X1  g331(.A1(new_n519), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT75), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT30), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n529), .ZN(new_n539));
  INV_X1    g338(.A(new_n532), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n474), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT69), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT68), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n441), .B1(new_n499), .B2(new_n516), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT25), .A4(new_n481), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n489), .B1(G183gat), .B2(G190gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(KEYINPUT65), .B2(new_n485), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n550), .B2(new_n496), .ZN(new_n551));
  INV_X1    g350(.A(new_n492), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n482), .B2(new_n490), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n443), .B(new_n525), .C1(new_n551), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n546), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI211_X1 g357(.A(KEYINPUT68), .B(new_n556), .C1(new_n547), .C2(new_n554), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n544), .B(new_n545), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G15gat), .B(G43gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(G71gat), .B(G99gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT32), .B1(new_n558), .B2(new_n559), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n554), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n443), .B1(new_n524), .B2(new_n525), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n557), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT68), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n546), .A3(new_n557), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n544), .B1(new_n572), .B2(new_n545), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT70), .B1(new_n566), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n563), .B1(new_n572), .B2(KEYINPUT32), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n545), .B1(new_n558), .B2(new_n559), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT69), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT70), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n575), .A2(new_n577), .A3(new_n578), .A4(new_n560), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n547), .A2(new_n556), .A3(new_n554), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT73), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(KEYINPUT73), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT34), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n585), .B1(new_n556), .B2(KEYINPUT72), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(new_n586), .A3(new_n583), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(KEYINPUT74), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT71), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n563), .A2(new_n545), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n565), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n572), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n590), .A2(KEYINPUT74), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n580), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n591), .B1(new_n580), .B2(new_n597), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n426), .B(new_n543), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT35), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n536), .A2(new_n602), .A3(new_n538), .A4(new_n541), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n473), .A2(KEYINPUT84), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT84), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n472), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n426), .B(new_n607), .C1(new_n598), .C2(new_n599), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT86), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n580), .A2(new_n597), .ZN(new_n611));
  INV_X1    g410(.A(new_n591), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n580), .A2(new_n591), .A3(new_n597), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n615), .A2(KEYINPUT86), .A3(new_n426), .A4(new_n607), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n610), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n519), .A2(new_n529), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n618), .B1(new_n519), .B2(new_n529), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n532), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT83), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n625), .A2(new_n627), .A3(new_n533), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(KEYINPUT85), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT85), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(new_n622), .B2(new_n532), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n631), .A3(new_n619), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT38), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n628), .A2(new_n604), .A3(new_n606), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n458), .A2(new_n449), .ZN(new_n636));
  INV_X1    g435(.A(new_n459), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n635), .B(new_n455), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n638), .A2(new_n466), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n455), .B1(new_n636), .B2(new_n637), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n452), .A2(new_n453), .A3(new_n447), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT39), .B1(new_n641), .B2(KEYINPUT82), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(KEYINPUT82), .B2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(KEYINPUT40), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n468), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT40), .B1(new_n639), .B2(new_n644), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n425), .B1(new_n648), .B2(new_n542), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n423), .A2(KEYINPUT81), .A3(new_n424), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT81), .B1(new_n423), .B2(new_n424), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n543), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n634), .A2(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n598), .A2(new_n599), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT36), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n615), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n654), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n617), .A2(KEYINPUT87), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT87), .B1(new_n617), .B2(new_n659), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n269), .B(new_n359), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n473), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n234), .ZN(G1324gat));
  INV_X1    g463(.A(new_n269), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n617), .A2(new_n659), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT87), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n617), .A2(new_n659), .A3(KEYINPUT87), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n665), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  NAND4_X1  g470(.A1(new_n670), .A2(new_n542), .A3(new_n359), .A4(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n542), .ZN(new_n673));
  OAI21_X1  g472(.A(G8gat), .B1(new_n662), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n672), .ZN(new_n675));
  MUX2_X1   g474(.A(new_n672), .B(new_n675), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n658), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G15gat), .B1(new_n662), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n670), .A2(new_n680), .A3(new_n615), .A4(new_n359), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(G1326gat));
  INV_X1    g481(.A(new_n652), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n662), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT43), .B(G22gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n310), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n660), .B2(new_n661), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n309), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n687), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n339), .A2(new_n340), .ZN(new_n692));
  INV_X1    g491(.A(new_n358), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n665), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n689), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G29gat), .B1(new_n696), .B2(new_n473), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n694), .A2(new_n310), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n269), .B(new_n699), .C1(new_n660), .C2(new_n661), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n473), .A2(G29gat), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n700), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n701), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n697), .A2(new_n703), .A3(new_n705), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n708));
  NOR4_X1   g507(.A1(new_n694), .A2(new_n310), .A3(G36gat), .A4(new_n673), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n670), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n269), .B(new_n709), .C1(new_n660), .C2(new_n661), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT102), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n707), .B1(new_n713), .B2(KEYINPUT46), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(KEYINPUT46), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n710), .A2(new_n712), .A3(KEYINPUT103), .A4(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G36gat), .B1(new_n696), .B2(new_n673), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n714), .A2(new_n715), .A3(new_n717), .A4(new_n718), .ZN(G1329gat));
  XNOR2_X1  g518(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n689), .A2(new_n677), .A3(new_n691), .A4(new_n695), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(G43gat), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n655), .A2(G43gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT105), .B1(new_n700), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n670), .A2(new_n726), .A3(new_n699), .A4(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n720), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n721), .A2(G43gat), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n730), .B(KEYINPUT47), .C1(new_n700), .C2(new_n724), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1330gat));
  OAI21_X1  g531(.A(G50gat), .B1(new_n696), .B2(new_n426), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n683), .A2(G50gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n704), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT48), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n689), .A2(new_n652), .A3(new_n691), .A4(new_n695), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n737), .A2(G50gat), .B1(new_n704), .B2(new_n734), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(KEYINPUT48), .B2(new_n738), .ZN(G1331gat));
  NOR3_X1   g538(.A1(new_n342), .A2(new_n269), .A3(new_n693), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n666), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n473), .B(KEYINPUT106), .Z(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g545(.A1(new_n741), .A2(new_n673), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  NOR2_X1   g550(.A1(new_n741), .A2(new_n655), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n753));
  INV_X1    g552(.A(G71gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n752), .B2(KEYINPUT108), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n678), .A2(new_n754), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n742), .B2(new_n757), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n741), .A2(KEYINPUT107), .A3(new_n754), .A4(new_n678), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n753), .A2(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT50), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n762));
  OAI221_X1 g561(.A(new_n762), .B1(new_n758), .B2(new_n759), .C1(new_n753), .C2(new_n755), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n742), .A2(new_n652), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n341), .A2(new_n269), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n358), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT109), .Z(new_n769));
  NAND3_X1  g568(.A1(new_n689), .A2(new_n691), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n473), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n666), .A2(new_n309), .A3(new_n767), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n310), .B1(new_n617), .B2(new_n659), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(KEYINPUT110), .A3(new_n776), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n358), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n474), .A2(new_n275), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n771), .B1(new_n781), .B2(new_n782), .ZN(G1336gat));
  NAND4_X1  g582(.A1(new_n689), .A2(new_n542), .A3(new_n691), .A4(new_n769), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n777), .A2(new_n276), .A3(new_n542), .A4(new_n358), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1337gat));
  OAI21_X1  g591(.A(G99gat), .B1(new_n770), .B2(new_n678), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n655), .A2(G99gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n781), .B2(new_n794), .ZN(G1338gat));
  NOR3_X1   g594(.A1(new_n693), .A2(G106gat), .A3(new_n426), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n772), .A2(new_n773), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n775), .B2(new_n767), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT112), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n777), .A2(new_n802), .A3(new_n796), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n689), .A2(new_n425), .A3(new_n691), .A4(new_n769), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(G106gat), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n689), .A2(new_n652), .A3(new_n691), .A4(new_n769), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n807), .A2(G106gat), .B1(new_n777), .B2(new_n796), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n804), .A2(new_n806), .B1(new_n801), .B2(new_n808), .ZN(G1339gat));
  NOR4_X1   g608(.A1(new_n692), .A2(new_n309), .A3(new_n269), .A4(new_n358), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n348), .A2(new_n349), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n343), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n348), .A2(new_n344), .A3(new_n349), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n812), .A2(KEYINPUT113), .A3(KEYINPUT54), .A4(new_n813), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n355), .B1(new_n350), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n357), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n255), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n243), .A2(new_n253), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n244), .B1(new_n243), .B2(new_n249), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n263), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n268), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n268), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n821), .A2(new_n824), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n341), .B1(new_n833), .B2(new_n309), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n821), .A2(new_n269), .A3(new_n824), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n268), .A2(new_n828), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n836), .A2(new_n358), .B1(new_n306), .B2(new_n308), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n810), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n615), .A2(new_n673), .A3(new_n426), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n839), .A2(new_n743), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT115), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n429), .A3(new_n269), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n833), .A2(new_n309), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n838), .A3(new_n692), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n310), .A2(new_n665), .A3(new_n341), .A4(new_n693), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n655), .B(new_n652), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n473), .A2(new_n542), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n665), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n843), .A2(new_n850), .ZN(G1340gat));
  NAND3_X1  g650(.A1(new_n842), .A2(new_n427), .A3(new_n358), .ZN(new_n852));
  OAI21_X1  g651(.A(G120gat), .B1(new_n849), .B2(new_n693), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n849), .B2(new_n692), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n841), .A2(new_n435), .A3(new_n341), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n857), .B(new_n858), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n841), .A2(new_n433), .A3(new_n309), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n849), .B2(new_n310), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n846), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n677), .A2(new_n542), .A3(new_n426), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n744), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n269), .A2(new_n388), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT118), .Z(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n865), .A2(new_n872), .A3(new_n425), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n678), .A2(new_n848), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n683), .B1(new_n845), .B2(new_n846), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n872), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n874), .A2(new_n878), .A3(new_n665), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n871), .B1(new_n879), .B2(new_n390), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n871), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OAI221_X1 g683(.A(new_n871), .B1(new_n882), .B2(new_n881), .C1(new_n879), .C2(new_n390), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1344gat));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n396), .A3(new_n358), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT57), .B1(new_n839), .B2(new_n426), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n865), .A2(new_n872), .A3(new_n652), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n693), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n889), .A2(KEYINPUT119), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(G148gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n888), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n873), .B(new_n876), .C1(new_n872), .C2(new_n877), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI211_X1 g698(.A(KEYINPUT59), .B(new_n396), .C1(new_n899), .C2(new_n358), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n887), .B1(new_n897), .B2(new_n900), .ZN(G1345gat));
  NAND4_X1  g700(.A1(new_n865), .A2(new_n866), .A3(new_n341), .A4(new_n744), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n376), .B1(new_n902), .B2(KEYINPUT120), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n341), .A2(G155gat), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n903), .A2(new_n904), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n906), .B(new_n907), .ZN(G1346gat));
  NAND3_X1  g707(.A1(new_n868), .A2(new_n377), .A3(new_n309), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n898), .B2(new_n310), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G162gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n898), .A2(new_n910), .A3(new_n310), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(G1347gat));
  NAND3_X1  g713(.A1(new_n615), .A2(new_n542), .A3(new_n426), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n839), .A2(new_n474), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n269), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n743), .A2(new_n542), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT123), .Z(new_n919));
  NAND2_X1  g718(.A1(new_n847), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n665), .A2(new_n476), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(G1348gat));
  OAI21_X1  g722(.A(G176gat), .B1(new_n920), .B2(new_n693), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n916), .A2(new_n477), .A3(new_n358), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n920), .B2(new_n692), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n916), .A2(new_n514), .A3(new_n341), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n916), .A2(new_n487), .A3(new_n309), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n921), .A2(new_n309), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(G190gat), .ZN(new_n934));
  AOI211_X1 g733(.A(KEYINPUT61), .B(new_n487), .C1(new_n921), .C2(new_n309), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(G1351gat));
  AND2_X1   g735(.A1(new_n889), .A2(new_n890), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n678), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT125), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n919), .A2(new_n940), .A3(new_n678), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n937), .A2(new_n269), .A3(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT124), .B(G197gat), .Z(new_n944));
  NOR2_X1   g743(.A1(new_n839), .A2(new_n474), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n677), .A2(new_n673), .A3(new_n426), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n269), .A2(new_n944), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n943), .A2(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  XNOR2_X1  g748(.A(KEYINPUT126), .B(G204gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n947), .A2(new_n693), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n358), .A3(new_n942), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1353gat));
  NAND4_X1  g754(.A1(new_n945), .A2(new_n365), .A3(new_n341), .A4(new_n946), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n937), .A2(new_n341), .A3(new_n942), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  AND3_X1   g759(.A1(new_n937), .A2(new_n309), .A3(new_n942), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n309), .A2(new_n366), .ZN(new_n962));
  OAI22_X1  g761(.A1(new_n961), .A2(new_n366), .B1(new_n947), .B2(new_n962), .ZN(G1355gat));
endmodule


