

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736;

  XNOR2_X1 U371 ( .A(n380), .B(KEYINPUT22), .ZN(n517) );
  XNOR2_X1 U372 ( .A(n458), .B(n457), .ZN(n618) );
  XNOR2_X1 U373 ( .A(n424), .B(n414), .ZN(n441) );
  XNOR2_X1 U374 ( .A(KEYINPUT4), .B(KEYINPUT67), .ZN(n440) );
  OR2_X2 U375 ( .A1(n694), .A2(n515), .ZN(n366) );
  INV_X1 U376 ( .A(G953), .ZN(n712) );
  XNOR2_X2 U377 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n390) );
  NOR2_X1 U378 ( .A1(n517), .A2(n386), .ZN(n385) );
  INV_X1 U379 ( .A(G101), .ZN(n378) );
  XNOR2_X1 U380 ( .A(n551), .B(KEYINPUT112), .ZN(n736) );
  OR2_X1 U381 ( .A1(n517), .A2(n671), .ZN(n510) );
  NOR2_X1 U382 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U383 ( .A(n439), .B(KEYINPUT41), .ZN(n693) );
  XNOR2_X1 U384 ( .A(n449), .B(n448), .ZN(n564) );
  XNOR2_X1 U385 ( .A(n351), .B(G107), .ZN(n711) );
  XNOR2_X1 U386 ( .A(n378), .B(KEYINPUT71), .ZN(n429) );
  NOR2_X1 U387 ( .A1(n389), .A2(G953), .ZN(n388) );
  INV_X2 U388 ( .A(G143), .ZN(n362) );
  NOR2_X2 U389 ( .A1(n592), .A2(n721), .ZN(n593) );
  NAND2_X2 U390 ( .A1(n591), .A2(n590), .ZN(n721) );
  XNOR2_X2 U391 ( .A(G146), .B(G125), .ZN(n423) );
  INV_X1 U392 ( .A(n538), .ZN(n373) );
  XOR2_X1 U393 ( .A(G131), .B(G140), .Z(n443) );
  INV_X1 U394 ( .A(G224), .ZN(n389) );
  INV_X1 U395 ( .A(KEYINPUT30), .ZN(n370) );
  AND2_X1 U396 ( .A1(n468), .A2(n467), .ZN(n538) );
  NOR2_X1 U397 ( .A1(G900), .A2(n464), .ZN(n465) );
  INV_X1 U398 ( .A(KEYINPUT90), .ZN(n360) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n452) );
  XOR2_X1 U400 ( .A(G131), .B(KEYINPUT98), .Z(n451) );
  XNOR2_X1 U401 ( .A(n440), .B(G137), .ZN(n442) );
  XNOR2_X1 U402 ( .A(n430), .B(n393), .ZN(n456) );
  XNOR2_X1 U403 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U404 ( .A(G116), .B(G113), .ZN(n428) );
  XNOR2_X1 U405 ( .A(n423), .B(KEYINPUT10), .ZN(n479) );
  XNOR2_X1 U406 ( .A(n711), .B(KEYINPUT72), .ZN(n445) );
  NOR2_X1 U407 ( .A1(n557), .A2(n556), .ZN(n581) );
  INV_X1 U408 ( .A(G902), .ZN(n459) );
  INV_X1 U409 ( .A(n564), .ZN(n377) );
  AND2_X1 U410 ( .A1(n686), .A2(n554), .ZN(n439) );
  INV_X1 U411 ( .A(n520), .ZN(n515) );
  XNOR2_X1 U412 ( .A(n501), .B(n500), .ZN(n565) );
  XNOR2_X1 U413 ( .A(G478), .B(n421), .ZN(n527) );
  OR2_X1 U414 ( .A1(n634), .A2(G902), .ZN(n492) );
  NOR2_X1 U415 ( .A1(G237), .A2(G902), .ZN(n434) );
  XNOR2_X1 U416 ( .A(G902), .B(KEYINPUT89), .ZN(n433) );
  XOR2_X1 U417 ( .A(KEYINPUT12), .B(G104), .Z(n402) );
  XNOR2_X1 U418 ( .A(G143), .B(G113), .ZN(n401) );
  XOR2_X1 U419 ( .A(G122), .B(KEYINPUT11), .Z(n400) );
  NAND2_X1 U420 ( .A1(G234), .A2(G237), .ZN(n461) );
  NAND2_X1 U421 ( .A1(n372), .A2(n369), .ZN(n540) );
  XNOR2_X1 U422 ( .A(n371), .B(n370), .ZN(n369) );
  AND2_X1 U423 ( .A1(n539), .A2(n373), .ZN(n372) );
  AND2_X1 U424 ( .A1(n512), .A2(n511), .ZN(n670) );
  XNOR2_X1 U425 ( .A(G128), .B(KEYINPUT78), .ZN(n480) );
  XNOR2_X1 U426 ( .A(G140), .B(KEYINPUT23), .ZN(n477) );
  XNOR2_X1 U427 ( .A(KEYINPUT24), .B(G137), .ZN(n476) );
  XOR2_X1 U428 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n417) );
  XNOR2_X1 U429 ( .A(G116), .B(G107), .ZN(n409) );
  XOR2_X1 U430 ( .A(KEYINPUT100), .B(G122), .Z(n410) );
  XNOR2_X1 U431 ( .A(KEYINPUT7), .B(KEYINPUT102), .ZN(n411) );
  INV_X1 U432 ( .A(G134), .ZN(n414) );
  XNOR2_X1 U433 ( .A(n445), .B(n387), .ZN(n447) );
  XNOR2_X1 U434 ( .A(n444), .B(n446), .ZN(n387) );
  INV_X1 U435 ( .A(KEYINPUT34), .ZN(n365) );
  AND2_X1 U436 ( .A1(n670), .A2(n377), .ZN(n539) );
  XNOR2_X1 U437 ( .A(n356), .B(n392), .ZN(n391) );
  INV_X1 U438 ( .A(KEYINPUT0), .ZN(n392) );
  INV_X1 U439 ( .A(KEYINPUT64), .ZN(n358) );
  AND2_X1 U440 ( .A1(n606), .A2(G953), .ZN(n703) );
  INV_X1 U441 ( .A(KEYINPUT42), .ZN(n374) );
  OR2_X1 U442 ( .A1(n693), .A2(n376), .ZN(n375) );
  NAND2_X1 U443 ( .A1(n355), .A2(n377), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n367), .B(KEYINPUT40), .ZN(n542) );
  NAND2_X1 U445 ( .A1(n368), .A2(n395), .ZN(n367) );
  XNOR2_X1 U446 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n734) );
  INV_X1 U448 ( .A(KEYINPUT32), .ZN(n383) );
  NAND2_X1 U449 ( .A1(n379), .A2(n352), .ZN(n645) );
  INV_X1 U450 ( .A(n510), .ZN(n379) );
  XOR2_X1 U451 ( .A(G110), .B(G104), .Z(n351) );
  AND2_X2 U452 ( .A1(n601), .A2(n657), .ZN(n633) );
  AND2_X1 U453 ( .A1(n669), .A2(n666), .ZN(n352) );
  XNOR2_X1 U454 ( .A(KEYINPUT105), .B(n516), .ZN(n353) );
  XOR2_X1 U455 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n354) );
  XOR2_X1 U456 ( .A(n497), .B(n496), .Z(n355) );
  XNOR2_X1 U457 ( .A(KEYINPUT87), .B(KEYINPUT66), .ZN(n356) );
  XNOR2_X1 U458 ( .A(KEYINPUT35), .B(KEYINPUT79), .ZN(n357) );
  XNOR2_X1 U459 ( .A(n600), .B(n358), .ZN(n601) );
  NAND2_X1 U460 ( .A1(n633), .A2(G472), .ZN(n620) );
  XNOR2_X1 U461 ( .A(n359), .B(n423), .ZN(n426) );
  XNOR2_X1 U462 ( .A(n388), .B(n390), .ZN(n359) );
  XNOR2_X1 U463 ( .A(n361), .B(n360), .ZN(n463) );
  NAND2_X1 U464 ( .A1(n466), .A2(G902), .ZN(n361) );
  XNOR2_X2 U465 ( .A(n718), .B(G146), .ZN(n458) );
  XNOR2_X2 U466 ( .A(n441), .B(n442), .ZN(n718) );
  XNOR2_X2 U467 ( .A(n362), .B(G128), .ZN(n424) );
  XNOR2_X2 U468 ( .A(n363), .B(n357), .ZN(n731) );
  NAND2_X1 U469 ( .A1(n364), .A2(n546), .ZN(n363) );
  XNOR2_X1 U470 ( .A(n366), .B(n365), .ZN(n364) );
  INV_X1 U471 ( .A(n542), .ZN(n735) );
  INV_X1 U472 ( .A(n589), .ZN(n368) );
  NAND2_X1 U473 ( .A1(n537), .A2(n554), .ZN(n371) );
  XNOR2_X2 U474 ( .A(n375), .B(n374), .ZN(n536) );
  NAND2_X1 U475 ( .A1(n508), .A2(n520), .ZN(n380) );
  NAND2_X1 U476 ( .A1(n385), .A2(n353), .ZN(n384) );
  NOR2_X1 U477 ( .A1(n594), .A2(n721), .ZN(n599) );
  NOR2_X2 U478 ( .A1(n437), .A2(n680), .ZN(n686) );
  AND2_X2 U479 ( .A1(n381), .A2(n731), .ZN(n519) );
  NOR2_X1 U480 ( .A1(n734), .A2(n382), .ZN(n381) );
  INV_X1 U481 ( .A(n645), .ZN(n382) );
  INV_X1 U482 ( .A(n518), .ZN(n386) );
  XNOR2_X2 U483 ( .A(n506), .B(n391), .ZN(n520) );
  XOR2_X2 U484 ( .A(n586), .B(KEYINPUT38), .Z(n680) );
  INV_X2 U485 ( .A(n558), .ZN(n586) );
  NOR2_X2 U486 ( .A1(n565), .A2(n505), .ZN(n506) );
  XNOR2_X1 U487 ( .A(G119), .B(KEYINPUT3), .ZN(n393) );
  AND2_X1 U488 ( .A1(G227), .A2(n712), .ZN(n394) );
  AND2_X1 U489 ( .A1(n527), .A2(n526), .ZN(n395) );
  AND2_X1 U490 ( .A1(n570), .A2(n569), .ZN(n396) );
  XOR2_X1 U491 ( .A(n585), .B(KEYINPUT109), .Z(n397) );
  NOR2_X1 U492 ( .A1(n729), .A2(n563), .ZN(n398) );
  NOR2_X1 U493 ( .A1(n396), .A2(n573), .ZN(n574) );
  XNOR2_X1 U494 ( .A(n443), .B(n394), .ZN(n444) );
  NAND2_X1 U495 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U496 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n499) );
  XNOR2_X1 U498 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U499 ( .A(KEYINPUT19), .ZN(n500) );
  XNOR2_X1 U500 ( .A(n408), .B(G475), .ZN(n525) );
  INV_X1 U501 ( .A(n525), .ZN(n526) );
  XNOR2_X1 U502 ( .A(n443), .B(n479), .ZN(n719) );
  NAND2_X1 U503 ( .A1(G214), .A2(n452), .ZN(n399) );
  XNOR2_X1 U504 ( .A(n400), .B(n399), .ZN(n404) );
  XNOR2_X1 U505 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U506 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U507 ( .A(n719), .B(n405), .ZN(n603) );
  NOR2_X1 U508 ( .A1(G902), .A2(n603), .ZN(n407) );
  XNOR2_X1 U509 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n406) );
  XNOR2_X1 U510 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U511 ( .A(n410), .B(n409), .ZN(n413) );
  XNOR2_X1 U512 ( .A(n354), .B(n411), .ZN(n412) );
  XNOR2_X1 U513 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U514 ( .A(n415), .B(n441), .Z(n420) );
  NAND2_X1 U515 ( .A1(G234), .A2(n712), .ZN(n416) );
  XNOR2_X1 U516 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U517 ( .A(n418), .B(KEYINPUT82), .ZN(n475) );
  NAND2_X1 U518 ( .A1(n475), .A2(G217), .ZN(n419) );
  XNOR2_X1 U519 ( .A(n420), .B(n419), .ZN(n700) );
  NOR2_X1 U520 ( .A1(n700), .A2(G902), .ZN(n421) );
  NAND2_X1 U521 ( .A1(n525), .A2(n527), .ZN(n422) );
  XOR2_X1 U522 ( .A(KEYINPUT104), .B(n422), .Z(n682) );
  INV_X1 U523 ( .A(n682), .ZN(n437) );
  XOR2_X1 U524 ( .A(n424), .B(n440), .Z(n425) );
  XNOR2_X1 U525 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U526 ( .A(n427), .B(n445), .ZN(n432) );
  XOR2_X1 U527 ( .A(G122), .B(KEYINPUT16), .Z(n431) );
  XNOR2_X1 U528 ( .A(n431), .B(n456), .ZN(n710) );
  XNOR2_X1 U529 ( .A(n432), .B(n710), .ZN(n625) );
  XNOR2_X1 U530 ( .A(n433), .B(KEYINPUT15), .ZN(n595) );
  NOR2_X1 U531 ( .A1(n625), .A2(n595), .ZN(n436) );
  XOR2_X1 U532 ( .A(KEYINPUT74), .B(n434), .Z(n438) );
  NAND2_X1 U533 ( .A1(G210), .A2(n438), .ZN(n435) );
  BUF_X1 U534 ( .A(n499), .Z(n558) );
  NAND2_X1 U535 ( .A1(n438), .A2(G214), .ZN(n554) );
  XNOR2_X1 U536 ( .A(G101), .B(KEYINPUT91), .ZN(n446) );
  XNOR2_X1 U537 ( .A(n458), .B(n447), .ZN(n612) );
  NOR2_X1 U538 ( .A1(n612), .A2(G902), .ZN(n449) );
  XNOR2_X1 U539 ( .A(KEYINPUT70), .B(G469), .ZN(n448) );
  XNOR2_X1 U540 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n450) );
  XNOR2_X1 U541 ( .A(n451), .B(n450), .ZN(n454) );
  NAND2_X1 U542 ( .A1(n452), .A2(G210), .ZN(n453) );
  NAND2_X1 U543 ( .A1(n618), .A2(n459), .ZN(n460) );
  XNOR2_X2 U544 ( .A(n460), .B(G472), .ZN(n537) );
  BUF_X1 U545 ( .A(n537), .Z(n522) );
  XOR2_X1 U546 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n462) );
  XNOR2_X1 U547 ( .A(n462), .B(n461), .ZN(n466) );
  NAND2_X1 U548 ( .A1(G953), .A2(n463), .ZN(n502) );
  XNOR2_X1 U549 ( .A(KEYINPUT106), .B(n502), .ZN(n464) );
  XNOR2_X1 U550 ( .A(n465), .B(KEYINPUT107), .ZN(n468) );
  NAND2_X1 U551 ( .A1(G952), .A2(n466), .ZN(n692) );
  NOR2_X1 U552 ( .A1(n692), .A2(G953), .ZN(n504) );
  INV_X1 U553 ( .A(n504), .ZN(n467) );
  INV_X1 U554 ( .A(G234), .ZN(n469) );
  OR2_X1 U555 ( .A1(n595), .A2(n469), .ZN(n471) );
  XOR2_X1 U556 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n470) );
  XNOR2_X1 U557 ( .A(n471), .B(n470), .ZN(n487) );
  NAND2_X1 U558 ( .A1(n487), .A2(G221), .ZN(n474) );
  INV_X1 U559 ( .A(KEYINPUT95), .ZN(n472) );
  XNOR2_X1 U560 ( .A(n472), .B(KEYINPUT21), .ZN(n473) );
  XNOR2_X1 U561 ( .A(n474), .B(n473), .ZN(n665) );
  NOR2_X1 U562 ( .A1(n538), .A2(n665), .ZN(n493) );
  NAND2_X1 U563 ( .A1(n475), .A2(G221), .ZN(n486) );
  XNOR2_X1 U564 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U565 ( .A(n479), .B(n478), .ZN(n484) );
  XNOR2_X1 U566 ( .A(n480), .B(G110), .ZN(n482) );
  XNOR2_X1 U567 ( .A(KEYINPUT92), .B(G119), .ZN(n481) );
  XNOR2_X1 U568 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U569 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n486), .B(n485), .ZN(n634) );
  NAND2_X1 U571 ( .A1(n487), .A2(G217), .ZN(n490) );
  XNOR2_X1 U572 ( .A(KEYINPUT77), .B(KEYINPUT94), .ZN(n488) );
  XNOR2_X1 U573 ( .A(n488), .B(KEYINPUT25), .ZN(n489) );
  XNOR2_X1 U574 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U575 ( .A(n492), .B(n491), .ZN(n512) );
  INV_X1 U576 ( .A(n512), .ZN(n666) );
  NAND2_X1 U577 ( .A1(n493), .A2(n666), .ZN(n494) );
  XNOR2_X1 U578 ( .A(n494), .B(KEYINPUT69), .ZN(n555) );
  NAND2_X1 U579 ( .A1(n522), .A2(n555), .ZN(n497) );
  INV_X1 U580 ( .A(KEYINPUT113), .ZN(n495) );
  XNOR2_X1 U581 ( .A(n495), .B(KEYINPUT28), .ZN(n496) );
  XOR2_X1 U582 ( .A(G137), .B(n536), .Z(G39) );
  XOR2_X2 U583 ( .A(KEYINPUT6), .B(n537), .Z(n553) );
  INV_X1 U584 ( .A(KEYINPUT1), .ZN(n498) );
  XNOR2_X1 U585 ( .A(n564), .B(n498), .ZN(n513) );
  INV_X1 U586 ( .A(n513), .ZN(n582) );
  INV_X1 U587 ( .A(n582), .ZN(n671) );
  NAND2_X1 U588 ( .A1(n499), .A2(n554), .ZN(n501) );
  NOR2_X1 U589 ( .A1(G898), .A2(n502), .ZN(n503) );
  NOR2_X1 U590 ( .A1(n504), .A2(n503), .ZN(n505) );
  INV_X1 U591 ( .A(KEYINPUT96), .ZN(n507) );
  XNOR2_X1 U592 ( .A(n665), .B(n507), .ZN(n511) );
  AND2_X1 U593 ( .A1(n682), .A2(n511), .ZN(n508) );
  NOR2_X1 U594 ( .A1(n386), .A2(n510), .ZN(n509) );
  AND2_X1 U595 ( .A1(n509), .A2(n512), .ZN(n532) );
  XOR2_X1 U596 ( .A(G101), .B(n532), .Z(G3) );
  INV_X1 U597 ( .A(n522), .ZN(n669) );
  NAND2_X1 U598 ( .A1(n513), .A2(n670), .ZN(n523) );
  INV_X1 U599 ( .A(n553), .ZN(n518) );
  NOR2_X2 U600 ( .A1(n523), .A2(n518), .ZN(n514) );
  XNOR2_X1 U601 ( .A(n514), .B(KEYINPUT33), .ZN(n694) );
  NOR2_X1 U602 ( .A1(n525), .A2(n527), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n671), .A2(n666), .ZN(n516) );
  XNOR2_X1 U604 ( .A(n519), .B(KEYINPUT44), .ZN(n534) );
  NAND2_X1 U605 ( .A1(n539), .A2(n520), .ZN(n521) );
  NOR2_X1 U606 ( .A1(n522), .A2(n521), .ZN(n641) );
  NOR2_X1 U607 ( .A1(n669), .A2(n523), .ZN(n676) );
  NAND2_X1 U608 ( .A1(n520), .A2(n676), .ZN(n524) );
  XNOR2_X1 U609 ( .A(KEYINPUT31), .B(n524), .ZN(n652) );
  NOR2_X1 U610 ( .A1(n641), .A2(n652), .ZN(n530) );
  NOR2_X1 U611 ( .A1(n526), .A2(n527), .ZN(n651) );
  NOR2_X1 U612 ( .A1(n651), .A2(n395), .ZN(n529) );
  INV_X1 U613 ( .A(KEYINPUT103), .ZN(n528) );
  XNOR2_X1 U614 ( .A(n529), .B(n528), .ZN(n679) );
  NOR2_X1 U615 ( .A1(n530), .A2(n679), .ZN(n531) );
  NOR2_X1 U616 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U617 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X2 U618 ( .A(n535), .B(KEYINPUT45), .ZN(n704) );
  NAND2_X1 U619 ( .A1(n704), .A2(KEYINPUT2), .ZN(n592) );
  INV_X1 U620 ( .A(n536), .ZN(n543) );
  XNOR2_X1 U621 ( .A(KEYINPUT76), .B(n540), .ZN(n547) );
  NOR2_X1 U622 ( .A1(n547), .A2(n680), .ZN(n541) );
  XNOR2_X1 U623 ( .A(n541), .B(KEYINPUT39), .ZN(n589) );
  NAND2_X1 U624 ( .A1(n543), .A2(n542), .ZN(n545) );
  INV_X1 U625 ( .A(KEYINPUT46), .ZN(n544) );
  XNOR2_X1 U626 ( .A(n545), .B(n544), .ZN(n578) );
  INV_X1 U627 ( .A(n546), .ZN(n550) );
  NOR2_X1 U628 ( .A1(n547), .A2(n586), .ZN(n548) );
  XNOR2_X1 U629 ( .A(n548), .B(KEYINPUT111), .ZN(n549) );
  INV_X1 U630 ( .A(KEYINPUT81), .ZN(n552) );
  XNOR2_X1 U631 ( .A(n736), .B(n552), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n395), .A2(n553), .ZN(n557) );
  INV_X1 U633 ( .A(n554), .ZN(n684) );
  NAND2_X1 U634 ( .A1(n581), .A2(n558), .ZN(n560) );
  XOR2_X1 U635 ( .A(KEYINPUT114), .B(KEYINPUT36), .Z(n559) );
  NAND2_X1 U636 ( .A1(n561), .A2(n671), .ZN(n562) );
  XNOR2_X1 U637 ( .A(KEYINPUT115), .B(n562), .ZN(n729) );
  NOR2_X1 U638 ( .A1(KEYINPUT80), .A2(KEYINPUT47), .ZN(n563) );
  NOR2_X1 U639 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U640 ( .A1(n566), .A2(n355), .ZN(n648) );
  INV_X1 U641 ( .A(KEYINPUT47), .ZN(n567) );
  NAND2_X1 U642 ( .A1(n648), .A2(n567), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n568), .A2(KEYINPUT80), .ZN(n570) );
  INV_X1 U644 ( .A(n679), .ZN(n569) );
  NAND2_X1 U645 ( .A1(n679), .A2(KEYINPUT80), .ZN(n571) );
  NAND2_X1 U646 ( .A1(n648), .A2(n571), .ZN(n572) );
  AND2_X1 U647 ( .A1(n572), .A2(KEYINPUT47), .ZN(n573) );
  NAND2_X1 U648 ( .A1(n398), .A2(n574), .ZN(n575) );
  NOR2_X1 U649 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n580) );
  INV_X1 U651 ( .A(KEYINPUT48), .ZN(n579) );
  XNOR2_X1 U652 ( .A(n580), .B(n579), .ZN(n591) );
  XNOR2_X1 U653 ( .A(KEYINPUT108), .B(n581), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U655 ( .A(n584), .B(KEYINPUT43), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n397), .A2(n586), .ZN(n587) );
  XNOR2_X1 U657 ( .A(n587), .B(KEYINPUT110), .ZN(n732) );
  INV_X1 U658 ( .A(n651), .ZN(n588) );
  OR2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n654) );
  AND2_X1 U660 ( .A1(n732), .A2(n654), .ZN(n590) );
  XNOR2_X1 U661 ( .A(n593), .B(KEYINPUT75), .ZN(n657) );
  NAND2_X1 U662 ( .A1(n704), .A2(n595), .ZN(n594) );
  XNOR2_X1 U663 ( .A(n595), .B(KEYINPUT84), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n596), .A2(KEYINPUT2), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT65), .ZN(n598) );
  NOR2_X1 U666 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n633), .A2(G475), .ZN(n605) );
  XOR2_X1 U668 ( .A(KEYINPUT88), .B(KEYINPUT59), .Z(n602) );
  XNOR2_X1 U669 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U670 ( .A(n605), .B(n604), .ZN(n607) );
  INV_X1 U671 ( .A(G952), .ZN(n606) );
  NOR2_X2 U672 ( .A1(n607), .A2(n703), .ZN(n609) );
  XNOR2_X1 U673 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n608) );
  XNOR2_X1 U674 ( .A(n609), .B(n608), .ZN(G60) );
  NAND2_X1 U675 ( .A1(n633), .A2(G469), .ZN(n614) );
  XOR2_X1 U676 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n610) );
  XNOR2_X1 U677 ( .A(n610), .B(KEYINPUT58), .ZN(n611) );
  XNOR2_X1 U678 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U679 ( .A(n614), .B(n613), .ZN(n615) );
  NOR2_X2 U680 ( .A1(n615), .A2(n703), .ZN(n617) );
  INV_X1 U681 ( .A(KEYINPUT123), .ZN(n616) );
  XNOR2_X1 U682 ( .A(n617), .B(n616), .ZN(G54) );
  XOR2_X1 U683 ( .A(KEYINPUT62), .B(n618), .Z(n619) );
  XNOR2_X1 U684 ( .A(n620), .B(n619), .ZN(n621) );
  NOR2_X2 U685 ( .A1(n621), .A2(n703), .ZN(n624) );
  XNOR2_X1 U686 ( .A(KEYINPUT116), .B(KEYINPUT63), .ZN(n622) );
  XNOR2_X1 U687 ( .A(n622), .B(KEYINPUT85), .ZN(n623) );
  XNOR2_X1 U688 ( .A(n624), .B(n623), .ZN(G57) );
  NAND2_X1 U689 ( .A1(n633), .A2(G210), .ZN(n630) );
  BUF_X1 U690 ( .A(n625), .Z(n628) );
  XNOR2_X1 U691 ( .A(KEYINPUT86), .B(KEYINPUT54), .ZN(n626) );
  XOR2_X1 U692 ( .A(n626), .B(KEYINPUT55), .Z(n627) );
  XNOR2_X1 U693 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U694 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U695 ( .A1(n631), .A2(n703), .ZN(n632) );
  XNOR2_X1 U696 ( .A(n632), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U697 ( .A1(n633), .A2(G217), .ZN(n635) );
  XNOR2_X1 U698 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X1 U699 ( .A1(n636), .A2(n703), .ZN(G66) );
  NAND2_X1 U700 ( .A1(n641), .A2(n395), .ZN(n637) );
  XNOR2_X1 U701 ( .A(n637), .B(G104), .ZN(G6) );
  XOR2_X1 U702 ( .A(KEYINPUT27), .B(KEYINPUT118), .Z(n639) );
  XNOR2_X1 U703 ( .A(G107), .B(KEYINPUT117), .ZN(n638) );
  XNOR2_X1 U704 ( .A(n639), .B(n638), .ZN(n640) );
  XOR2_X1 U705 ( .A(KEYINPUT26), .B(n640), .Z(n643) );
  NAND2_X1 U706 ( .A1(n641), .A2(n651), .ZN(n642) );
  XNOR2_X1 U707 ( .A(n643), .B(n642), .ZN(G9) );
  XOR2_X1 U708 ( .A(G110), .B(KEYINPUT119), .Z(n644) );
  XNOR2_X1 U709 ( .A(n645), .B(n644), .ZN(G12) );
  XOR2_X1 U710 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  NAND2_X1 U711 ( .A1(n648), .A2(n651), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(G30) );
  NAND2_X1 U713 ( .A1(n648), .A2(n395), .ZN(n649) );
  XNOR2_X1 U714 ( .A(n649), .B(G146), .ZN(G48) );
  NAND2_X1 U715 ( .A1(n652), .A2(n395), .ZN(n650) );
  XNOR2_X1 U716 ( .A(n650), .B(G113), .ZN(G15) );
  NAND2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U718 ( .A(n653), .B(G116), .ZN(G18) );
  INV_X1 U719 ( .A(n654), .ZN(n655) );
  XOR2_X1 U720 ( .A(G134), .B(n655), .Z(n656) );
  XNOR2_X1 U721 ( .A(KEYINPUT120), .B(n656), .ZN(G36) );
  INV_X1 U722 ( .A(n657), .ZN(n663) );
  NOR2_X1 U723 ( .A1(KEYINPUT2), .A2(n705), .ZN(n658) );
  XNOR2_X1 U724 ( .A(n658), .B(KEYINPUT83), .ZN(n661) );
  INV_X1 U725 ( .A(KEYINPUT2), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n721), .A2(n659), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n664), .A2(G953), .ZN(n698) );
  NAND2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U731 ( .A(KEYINPUT49), .B(n667), .Z(n668) );
  NAND2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n674) );
  NOR2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U734 ( .A(n672), .B(KEYINPUT50), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U737 ( .A(KEYINPUT51), .B(n677), .Z(n678) );
  NOR2_X1 U738 ( .A1(n693), .A2(n678), .ZN(n689) );
  NOR2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U741 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U742 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U743 ( .A1(n694), .A2(n687), .ZN(n688) );
  NOR2_X1 U744 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U746 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U747 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U748 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U749 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U750 ( .A(KEYINPUT53), .B(n699), .Z(G75) );
  NAND2_X1 U751 ( .A1(n633), .A2(G478), .ZN(n701) );
  XNOR2_X1 U752 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U753 ( .A1(n703), .A2(n702), .ZN(G63) );
  BUF_X1 U754 ( .A(n704), .Z(n705) );
  NAND2_X1 U755 ( .A1(n712), .A2(n705), .ZN(n709) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n706) );
  XNOR2_X1 U757 ( .A(KEYINPUT61), .B(n706), .ZN(n707) );
  NAND2_X1 U758 ( .A1(n707), .A2(G898), .ZN(n708) );
  NAND2_X1 U759 ( .A1(n709), .A2(n708), .ZN(n716) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(n714) );
  NOR2_X1 U761 ( .A1(G898), .A2(n712), .ZN(n713) );
  NOR2_X1 U762 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U763 ( .A(n716), .B(n715), .ZN(n717) );
  XOR2_X1 U764 ( .A(KEYINPUT125), .B(n717), .Z(G69) );
  XOR2_X1 U765 ( .A(KEYINPUT126), .B(n718), .Z(n720) );
  XOR2_X1 U766 ( .A(n720), .B(n719), .Z(n724) );
  XNOR2_X1 U767 ( .A(n721), .B(n724), .ZN(n722) );
  NOR2_X1 U768 ( .A1(n722), .A2(G953), .ZN(n723) );
  XNOR2_X1 U769 ( .A(KEYINPUT127), .B(n723), .ZN(n728) );
  XOR2_X1 U770 ( .A(G227), .B(n724), .Z(n725) );
  NAND2_X1 U771 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n726), .A2(G953), .ZN(n727) );
  NAND2_X1 U773 ( .A1(n728), .A2(n727), .ZN(G72) );
  XNOR2_X1 U774 ( .A(G125), .B(n729), .ZN(n730) );
  XNOR2_X1 U775 ( .A(n730), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U776 ( .A(n731), .B(G122), .ZN(G24) );
  XOR2_X1 U777 ( .A(G140), .B(n732), .Z(n733) );
  XNOR2_X1 U778 ( .A(KEYINPUT121), .B(n733), .ZN(G42) );
  XOR2_X1 U779 ( .A(G119), .B(n734), .Z(G21) );
  XOR2_X1 U780 ( .A(G131), .B(n735), .Z(G33) );
  XOR2_X1 U781 ( .A(G143), .B(n736), .Z(G45) );
endmodule

