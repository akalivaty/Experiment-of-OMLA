

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764;

  AND2_X1 U379 ( .A1(n574), .A2(n573), .ZN(n597) );
  BUF_X1 U380 ( .A(n678), .Z(n359) );
  XNOR2_X1 U381 ( .A(n555), .B(n554), .ZN(n663) );
  OR2_X1 U382 ( .A1(n678), .A2(n575), .ZN(n553) );
  XNOR2_X1 U383 ( .A(n499), .B(KEYINPUT1), .ZN(n678) );
  XNOR2_X1 U384 ( .A(n422), .B(n421), .ZN(n499) );
  XOR2_X1 U385 ( .A(G110), .B(KEYINPUT77), .Z(n433) );
  XNOR2_X2 U386 ( .A(n681), .B(KEYINPUT6), .ZN(n545) );
  NAND2_X1 U387 ( .A1(n609), .A2(KEYINPUT90), .ZN(n603) );
  AND2_X2 U388 ( .A1(n617), .A2(n753), .ZN(n609) );
  XNOR2_X1 U389 ( .A(G116), .B(G131), .ZN(n369) );
  XOR2_X1 U390 ( .A(G131), .B(G140), .Z(n447) );
  XNOR2_X1 U391 ( .A(n578), .B(n577), .ZN(n659) );
  NOR2_X2 U392 ( .A1(n570), .A2(KEYINPUT65), .ZN(n567) );
  NAND2_X2 U393 ( .A1(n612), .A2(n611), .ZN(n619) );
  NOR2_X2 U394 ( .A1(n553), .A2(n589), .ZN(n555) );
  XNOR2_X2 U395 ( .A(n365), .B(KEYINPUT3), .ZN(n367) );
  XNOR2_X2 U396 ( .A(n367), .B(n366), .ZN(n427) );
  INV_X2 U397 ( .A(G953), .ZN(n754) );
  NOR2_X1 U398 ( .A1(n593), .A2(n643), .ZN(n595) );
  OR2_X1 U399 ( .A1(n659), .A2(n646), .ZN(n586) );
  XNOR2_X2 U400 ( .A(n599), .B(n598), .ZN(n617) );
  XNOR2_X1 U401 ( .A(n429), .B(KEYINPUT10), .ZN(n446) );
  XNOR2_X1 U402 ( .A(n360), .B(KEYINPUT93), .ZN(n596) );
  NAND2_X1 U403 ( .A1(n595), .A2(n594), .ZN(n360) );
  XOR2_X2 U404 ( .A(G122), .B(G104), .Z(n448) );
  NOR2_X2 U405 ( .A1(n495), .A2(n494), .ZN(n525) );
  INV_X1 U406 ( .A(G101), .ZN(n414) );
  AND2_X1 U407 ( .A1(n626), .A2(G953), .ZN(n738) );
  XNOR2_X1 U408 ( .A(n446), .B(n389), .ZN(n392) );
  XNOR2_X1 U409 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n410) );
  XNOR2_X1 U410 ( .A(n471), .B(KEYINPUT41), .ZN(n690) );
  XNOR2_X1 U411 ( .A(n480), .B(KEYINPUT39), .ZN(n529) );
  BUF_X1 U412 ( .A(n575), .Z(n679) );
  XNOR2_X1 U413 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U414 ( .A(n727), .B(KEYINPUT120), .ZN(n728) );
  INV_X1 U415 ( .A(n731), .ZN(n726) );
  BUF_X1 U416 ( .A(n620), .Z(n623) );
  INV_X1 U417 ( .A(n635), .ZN(n565) );
  AND2_X1 U418 ( .A1(n546), .A2(n589), .ZN(n361) );
  XOR2_X2 U419 ( .A(KEYINPUT4), .B(KEYINPUT64), .Z(n362) );
  XOR2_X1 U420 ( .A(n370), .B(n369), .Z(n363) );
  XNOR2_X1 U421 ( .A(n527), .B(KEYINPUT38), .ZN(n692) );
  NOR2_X1 U422 ( .A1(n508), .A2(n481), .ZN(n364) );
  INV_X1 U423 ( .A(KEYINPUT44), .ZN(n564) );
  NOR2_X1 U424 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U425 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U426 ( .A(n485), .B(KEYINPUT46), .ZN(n522) );
  XNOR2_X1 U427 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U428 ( .A(n420), .B(n709), .ZN(n421) );
  NOR2_X1 U429 ( .A1(n695), .A2(n694), .ZN(n471) );
  INV_X1 U430 ( .A(n513), .ZN(n650) );
  BUF_X1 U431 ( .A(n650), .Z(n654) );
  XNOR2_X1 U432 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X2 U433 ( .A(G119), .B(G113), .ZN(n365) );
  XNOR2_X1 U434 ( .A(G101), .B(KEYINPUT75), .ZN(n366) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n450) );
  NAND2_X1 U436 ( .A1(n450), .A2(G210), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n427), .B(n368), .ZN(n371) );
  XOR2_X1 U438 ( .A(KEYINPUT5), .B(KEYINPUT100), .Z(n370) );
  XNOR2_X1 U439 ( .A(n371), .B(n363), .ZN(n377) );
  XNOR2_X1 U440 ( .A(G137), .B(n362), .ZN(n376) );
  INV_X1 U441 ( .A(G143), .ZN(n372) );
  NAND2_X1 U442 ( .A1(G128), .A2(n372), .ZN(n375) );
  INV_X1 U443 ( .A(G128), .ZN(n373) );
  NAND2_X1 U444 ( .A1(n373), .A2(G143), .ZN(n374) );
  NAND2_X1 U445 ( .A1(n375), .A2(n374), .ZN(n434) );
  XNOR2_X1 U446 ( .A(n434), .B(G134), .ZN(n459) );
  XNOR2_X1 U447 ( .A(n376), .B(n459), .ZN(n752) );
  XNOR2_X1 U448 ( .A(n752), .B(G146), .ZN(n419) );
  XNOR2_X1 U449 ( .A(n377), .B(n419), .ZN(n637) );
  INV_X1 U450 ( .A(G902), .ZN(n442) );
  NAND2_X1 U451 ( .A1(n637), .A2(n442), .ZN(n378) );
  INV_X1 U452 ( .A(G472), .ZN(n636) );
  XNOR2_X2 U453 ( .A(n378), .B(n636), .ZN(n681) );
  INV_X1 U454 ( .A(n681), .ZN(n580) );
  XNOR2_X1 U455 ( .A(G902), .B(KEYINPUT15), .ZN(n606) );
  NAND2_X1 U456 ( .A1(n606), .A2(G234), .ZN(n380) );
  INV_X1 U457 ( .A(KEYINPUT20), .ZN(n379) );
  XNOR2_X1 U458 ( .A(n380), .B(n379), .ZN(n402) );
  INV_X1 U459 ( .A(G221), .ZN(n381) );
  OR2_X1 U460 ( .A1(n402), .A2(n381), .ZN(n382) );
  XNOR2_X1 U461 ( .A(n382), .B(KEYINPUT21), .ZN(n675) );
  XOR2_X1 U462 ( .A(KEYINPUT14), .B(KEYINPUT98), .Z(n384) );
  NAND2_X1 U463 ( .A1(G234), .A2(G237), .ZN(n383) );
  XOR2_X1 U464 ( .A(n384), .B(n383), .Z(n385) );
  NAND2_X1 U465 ( .A1(G952), .A2(n385), .ZN(n705) );
  NOR2_X1 U466 ( .A1(n705), .A2(G953), .ZN(n532) );
  AND2_X1 U467 ( .A1(n385), .A2(G953), .ZN(n386) );
  NAND2_X1 U468 ( .A1(G902), .A2(n386), .ZN(n533) );
  NOR2_X1 U469 ( .A1(G900), .A2(n533), .ZN(n387) );
  NOR2_X1 U470 ( .A1(n532), .A2(n387), .ZN(n478) );
  NOR2_X1 U471 ( .A1(n675), .A2(n478), .ZN(n388) );
  XNOR2_X1 U472 ( .A(KEYINPUT72), .B(n388), .ZN(n408) );
  XNOR2_X2 U473 ( .A(G146), .B(G125), .ZN(n429) );
  XNOR2_X1 U474 ( .A(G140), .B(KEYINPUT76), .ZN(n389) );
  AND2_X1 U475 ( .A1(G234), .A2(n754), .ZN(n390) );
  XNOR2_X1 U476 ( .A(KEYINPUT8), .B(n390), .ZN(n465) );
  NAND2_X1 U477 ( .A1(n465), .A2(G221), .ZN(n391) );
  XNOR2_X1 U478 ( .A(n392), .B(n391), .ZN(n400) );
  XNOR2_X1 U479 ( .A(G119), .B(KEYINPUT24), .ZN(n394) );
  XNOR2_X1 U480 ( .A(G137), .B(G128), .ZN(n393) );
  XNOR2_X1 U481 ( .A(n394), .B(n393), .ZN(n398) );
  XNOR2_X1 U482 ( .A(G110), .B(KEYINPUT81), .ZN(n396) );
  XNOR2_X1 U483 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n395) );
  XNOR2_X1 U484 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U485 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U486 ( .A(n400), .B(n399), .ZN(n734) );
  INV_X1 U487 ( .A(n734), .ZN(n401) );
  NAND2_X1 U488 ( .A1(n401), .A2(n442), .ZN(n407) );
  INV_X1 U489 ( .A(G217), .ZN(n732) );
  OR2_X1 U490 ( .A1(n402), .A2(n732), .ZN(n405) );
  INV_X1 U491 ( .A(KEYINPUT99), .ZN(n403) );
  XNOR2_X1 U492 ( .A(n403), .B(KEYINPUT25), .ZN(n404) );
  XNOR2_X1 U493 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U494 ( .A(n407), .B(n406), .ZN(n543) );
  NAND2_X1 U495 ( .A1(n408), .A2(n543), .ZN(n409) );
  XNOR2_X1 U496 ( .A(n409), .B(KEYINPUT71), .ZN(n492) );
  NAND2_X1 U497 ( .A1(n580), .A2(n492), .ZN(n411) );
  XNOR2_X1 U498 ( .A(n411), .B(n410), .ZN(n424) );
  XOR2_X1 U499 ( .A(n447), .B(n433), .Z(n413) );
  XNOR2_X1 U500 ( .A(G104), .B(G107), .ZN(n412) );
  XNOR2_X1 U501 ( .A(n413), .B(n412), .ZN(n417) );
  NAND2_X1 U502 ( .A1(G227), .A2(n754), .ZN(n415) );
  XNOR2_X1 U503 ( .A(n418), .B(n419), .ZN(n713) );
  NOR2_X1 U504 ( .A1(G902), .A2(n713), .ZN(n422) );
  XNOR2_X1 U505 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n420) );
  INV_X1 U506 ( .A(G469), .ZN(n709) );
  BUF_X2 U507 ( .A(n499), .Z(n581) );
  XOR2_X1 U508 ( .A(n581), .B(KEYINPUT108), .Z(n423) );
  NAND2_X1 U509 ( .A1(n424), .A2(n423), .ZN(n502) );
  INV_X1 U510 ( .A(G122), .ZN(n633) );
  XNOR2_X1 U511 ( .A(n448), .B(KEYINPUT16), .ZN(n426) );
  INV_X1 U512 ( .A(G116), .ZN(n425) );
  XNOR2_X1 U513 ( .A(n425), .B(G107), .ZN(n464) );
  XNOR2_X1 U514 ( .A(n426), .B(n464), .ZN(n428) );
  XNOR2_X1 U515 ( .A(n428), .B(n427), .ZN(n743) );
  XOR2_X1 U516 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n431) );
  INV_X1 U517 ( .A(n429), .ZN(n430) );
  XNOR2_X1 U518 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U519 ( .A(n433), .B(n432), .ZN(n439) );
  XNOR2_X1 U520 ( .A(n362), .B(n434), .ZN(n437) );
  NAND2_X1 U521 ( .A1(G224), .A2(n754), .ZN(n435) );
  XNOR2_X1 U522 ( .A(n435), .B(KEYINPUT82), .ZN(n436) );
  XNOR2_X1 U523 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U524 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U525 ( .A(n743), .B(n440), .ZN(n620) );
  NAND2_X1 U526 ( .A1(n620), .A2(n606), .ZN(n444) );
  INV_X1 U527 ( .A(G237), .ZN(n441) );
  NAND2_X1 U528 ( .A1(n442), .A2(n441), .ZN(n445) );
  NAND2_X1 U529 ( .A1(n445), .A2(G210), .ZN(n443) );
  XNOR2_X2 U530 ( .A(n444), .B(n443), .ZN(n503) );
  BUF_X1 U531 ( .A(n503), .Z(n527) );
  NAND2_X1 U532 ( .A1(n445), .A2(G214), .ZN(n691) );
  NAND2_X1 U533 ( .A1(n692), .A2(n691), .ZN(n695) );
  XNOR2_X1 U534 ( .A(n447), .B(n446), .ZN(n750) );
  XNOR2_X1 U535 ( .A(G113), .B(G143), .ZN(n449) );
  XNOR2_X1 U536 ( .A(n449), .B(n448), .ZN(n454) );
  XOR2_X1 U537 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n452) );
  NAND2_X1 U538 ( .A1(G214), .A2(n450), .ZN(n451) );
  XNOR2_X1 U539 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U540 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U541 ( .A(n750), .B(n455), .ZN(n719) );
  NOR2_X1 U542 ( .A1(G902), .A2(n719), .ZN(n457) );
  XNOR2_X1 U543 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n456) );
  XNOR2_X1 U544 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U545 ( .A(G475), .ZN(n718) );
  XNOR2_X1 U546 ( .A(n458), .B(n718), .ZN(n508) );
  INV_X1 U547 ( .A(n459), .ZN(n463) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n461) );
  XNOR2_X1 U549 ( .A(G122), .B(KEYINPUT9), .ZN(n460) );
  XNOR2_X1 U550 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U551 ( .A(n463), .B(n462), .ZN(n469) );
  XOR2_X1 U552 ( .A(n464), .B(KEYINPUT103), .Z(n467) );
  NAND2_X1 U553 ( .A1(G217), .A2(n465), .ZN(n466) );
  XNOR2_X1 U554 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U555 ( .A(n469), .B(n468), .ZN(n727) );
  NOR2_X1 U556 ( .A1(G902), .A2(n727), .ZN(n470) );
  XNOR2_X1 U557 ( .A(n470), .B(G478), .ZN(n509) );
  NAND2_X1 U558 ( .A1(n508), .A2(n509), .ZN(n694) );
  NOR2_X1 U559 ( .A1(n502), .A2(n690), .ZN(n472) );
  XNOR2_X1 U560 ( .A(KEYINPUT42), .B(n472), .ZN(n764) );
  INV_X1 U561 ( .A(n764), .ZN(n484) );
  OR2_X2 U562 ( .A1(n543), .A2(n675), .ZN(n474) );
  INV_X1 U563 ( .A(KEYINPUT69), .ZN(n473) );
  XNOR2_X2 U564 ( .A(n474), .B(n473), .ZN(n575) );
  NOR2_X1 U565 ( .A1(n581), .A2(n679), .ZN(n475) );
  AND2_X1 U566 ( .A1(n475), .A2(n692), .ZN(n479) );
  NAND2_X1 U567 ( .A1(n580), .A2(n691), .ZN(n476) );
  XNOR2_X1 U568 ( .A(KEYINPUT30), .B(n476), .ZN(n477) );
  NOR2_X1 U569 ( .A1(n478), .A2(n477), .ZN(n489) );
  NAND2_X1 U570 ( .A1(n479), .A2(n489), .ZN(n480) );
  INV_X1 U571 ( .A(n509), .ZN(n481) );
  AND2_X1 U572 ( .A1(n529), .A2(n364), .ZN(n482) );
  XNOR2_X1 U573 ( .A(n482), .B(KEYINPUT40), .ZN(n762) );
  INV_X1 U574 ( .A(n762), .ZN(n483) );
  INV_X1 U575 ( .A(n581), .ZN(n486) );
  INV_X1 U576 ( .A(n527), .ZN(n496) );
  NAND2_X1 U577 ( .A1(n486), .A2(n496), .ZN(n487) );
  NOR2_X1 U578 ( .A1(n487), .A2(n679), .ZN(n488) );
  NAND2_X1 U579 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U580 ( .A(n490), .B(KEYINPUT107), .ZN(n491) );
  NOR2_X1 U581 ( .A1(n508), .A2(n509), .ZN(n561) );
  NAND2_X1 U582 ( .A1(n491), .A2(n561), .ZN(n653) );
  NAND2_X1 U583 ( .A1(n492), .A2(n545), .ZN(n493) );
  XNOR2_X1 U584 ( .A(n493), .B(KEYINPUT106), .ZN(n495) );
  NAND2_X1 U585 ( .A1(n364), .A2(n691), .ZN(n494) );
  NAND2_X1 U586 ( .A1(n525), .A2(n496), .ZN(n498) );
  XOR2_X1 U587 ( .A(KEYINPUT36), .B(KEYINPUT94), .Z(n497) );
  XNOR2_X1 U588 ( .A(n498), .B(n497), .ZN(n501) );
  INV_X1 U589 ( .A(KEYINPUT96), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n359), .B(n500), .ZN(n546) );
  NAND2_X1 U591 ( .A1(n501), .A2(n546), .ZN(n662) );
  NAND2_X1 U592 ( .A1(n653), .A2(n662), .ZN(n519) );
  INV_X1 U593 ( .A(n502), .ZN(n507) );
  INV_X1 U594 ( .A(n503), .ZN(n504) );
  NAND2_X1 U595 ( .A1(n504), .A2(n691), .ZN(n506) );
  XNOR2_X1 U596 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n505) );
  XNOR2_X2 U597 ( .A(n506), .B(n505), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n507), .A2(n537), .ZN(n513) );
  INV_X1 U599 ( .A(n508), .ZN(n510) );
  NOR2_X1 U600 ( .A1(n510), .A2(n509), .ZN(n658) );
  NOR2_X1 U601 ( .A1(n658), .A2(n364), .ZN(n696) );
  INV_X1 U602 ( .A(n696), .ZN(n585) );
  NAND2_X1 U603 ( .A1(n650), .A2(n585), .ZN(n511) );
  NAND2_X1 U604 ( .A1(n511), .A2(KEYINPUT88), .ZN(n512) );
  XNOR2_X1 U605 ( .A(n512), .B(KEYINPUT47), .ZN(n517) );
  INV_X1 U606 ( .A(KEYINPUT88), .ZN(n515) );
  NAND2_X1 U607 ( .A1(n513), .A2(n585), .ZN(n514) );
  NAND2_X1 U608 ( .A1(n515), .A2(n514), .ZN(n516) );
  NAND2_X1 U609 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U610 ( .A(KEYINPUT70), .B(n520), .Z(n521) );
  NOR2_X1 U611 ( .A1(n522), .A2(n521), .ZN(n524) );
  INV_X1 U612 ( .A(KEYINPUT48), .ZN(n523) );
  XNOR2_X1 U613 ( .A(n524), .B(n523), .ZN(n616) );
  NAND2_X1 U614 ( .A1(n525), .A2(n359), .ZN(n526) );
  XNOR2_X1 U615 ( .A(KEYINPUT43), .B(n526), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n528), .A2(n527), .ZN(n629) );
  NAND2_X1 U617 ( .A1(n658), .A2(n529), .ZN(n530) );
  XNOR2_X1 U618 ( .A(n530), .B(KEYINPUT110), .ZN(n763) );
  NAND2_X1 U619 ( .A1(n629), .A2(n763), .ZN(n531) );
  NOR2_X2 U620 ( .A1(n616), .A2(n531), .ZN(n753) );
  INV_X1 U621 ( .A(n532), .ZN(n535) );
  OR2_X1 U622 ( .A1(n533), .A2(G898), .ZN(n534) );
  NAND2_X1 U623 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U624 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U625 ( .A(n538), .B(KEYINPUT0), .ZN(n556) );
  OR2_X1 U626 ( .A1(n694), .A2(n675), .ZN(n539) );
  OR2_X2 U627 ( .A1(n556), .A2(n539), .ZN(n542) );
  XNOR2_X1 U628 ( .A(KEYINPUT80), .B(KEYINPUT22), .ZN(n540) );
  XNOR2_X1 U629 ( .A(n540), .B(KEYINPUT67), .ZN(n541) );
  XNOR2_X1 U630 ( .A(n542), .B(n541), .ZN(n592) );
  BUF_X1 U631 ( .A(n543), .Z(n544) );
  NAND2_X1 U632 ( .A1(n592), .A2(n544), .ZN(n552) );
  INV_X1 U633 ( .A(n552), .ZN(n547) );
  INV_X1 U634 ( .A(n545), .ZN(n589) );
  NAND2_X1 U635 ( .A1(n547), .A2(n361), .ZN(n550) );
  XNOR2_X1 U636 ( .A(KEYINPUT84), .B(KEYINPUT32), .ZN(n548) );
  XNOR2_X1 U637 ( .A(n548), .B(KEYINPUT66), .ZN(n549) );
  XNOR2_X2 U638 ( .A(n550), .B(n549), .ZN(n631) );
  NAND2_X1 U639 ( .A1(n359), .A2(n681), .ZN(n551) );
  OR2_X1 U640 ( .A1(n552), .A2(n551), .ZN(n630) );
  NAND2_X1 U641 ( .A1(n631), .A2(n630), .ZN(n570) );
  XNOR2_X1 U642 ( .A(KEYINPUT78), .B(KEYINPUT33), .ZN(n554) );
  BUF_X2 U643 ( .A(n556), .Z(n579) );
  NOR2_X1 U644 ( .A1(n663), .A2(n579), .ZN(n560) );
  XNOR2_X1 U645 ( .A(KEYINPUT83), .B(KEYINPUT34), .ZN(n558) );
  INV_X1 U646 ( .A(KEYINPUT79), .ZN(n557) );
  XOR2_X1 U647 ( .A(n558), .B(n557), .Z(n559) );
  XNOR2_X1 U648 ( .A(n560), .B(n559), .ZN(n562) );
  NAND2_X1 U649 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X2 U650 ( .A(n563), .B(KEYINPUT35), .ZN(n635) );
  NAND2_X1 U651 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U652 ( .A1(n567), .A2(n566), .ZN(n572) );
  INV_X1 U653 ( .A(KEYINPUT65), .ZN(n568) );
  NAND2_X1 U654 ( .A1(n568), .A2(KEYINPUT44), .ZN(n569) );
  NAND2_X1 U655 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U656 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U657 ( .A1(n564), .A2(KEYINPUT65), .ZN(n573) );
  OR2_X1 U658 ( .A1(n681), .A2(n575), .ZN(n576) );
  OR2_X2 U659 ( .A1(n678), .A2(n576), .ZN(n674) );
  NOR2_X2 U660 ( .A1(n674), .A2(n579), .ZN(n578) );
  XNOR2_X1 U661 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n577) );
  INV_X1 U662 ( .A(n579), .ZN(n584) );
  OR2_X1 U663 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U664 ( .A1(n582), .A2(n679), .ZN(n583) );
  AND2_X1 U665 ( .A1(n584), .A2(n583), .ZN(n646) );
  NAND2_X1 U666 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U667 ( .A(n587), .B(KEYINPUT105), .ZN(n593) );
  INV_X1 U668 ( .A(n544), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n359), .A2(n588), .ZN(n590) );
  NOR2_X1 U670 ( .A1(n590), .A2(n545), .ZN(n591) );
  AND2_X1 U671 ( .A1(n592), .A2(n591), .ZN(n643) );
  NAND2_X1 U672 ( .A1(n635), .A2(KEYINPUT44), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U674 ( .A(KEYINPUT92), .B(KEYINPUT45), .ZN(n598) );
  INV_X1 U675 ( .A(KEYINPUT2), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n600), .A2(KEYINPUT91), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n606), .A2(n601), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n608) );
  NAND2_X1 U679 ( .A1(KEYINPUT2), .A2(KEYINPUT91), .ZN(n604) );
  AND2_X1 U680 ( .A1(n604), .A2(KEYINPUT90), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n612) );
  INV_X1 U683 ( .A(n609), .ZN(n666) );
  INV_X1 U684 ( .A(KEYINPUT90), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n666), .A2(n610), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n763), .A2(KEYINPUT2), .ZN(n613) );
  XNOR2_X1 U687 ( .A(KEYINPUT85), .B(n613), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n614), .A2(n629), .ZN(n615) );
  NOR2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n665) );
  BUF_X1 U690 ( .A(n617), .Z(n618) );
  NAND2_X1 U691 ( .A1(n665), .A2(n618), .ZN(n667) );
  NAND2_X2 U692 ( .A1(n619), .A2(n667), .ZN(n731) );
  NAND2_X1 U693 ( .A1(n726), .A2(G210), .ZN(n625) );
  XOR2_X1 U694 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n621) );
  XOR2_X1 U695 ( .A(n621), .B(KEYINPUT86), .Z(n622) );
  XNOR2_X1 U696 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n627) );
  INV_X1 U698 ( .A(G952), .ZN(n626) );
  NOR2_X2 U699 ( .A1(n627), .A2(n738), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U701 ( .A(n629), .B(G140), .ZN(G42) );
  XNOR2_X1 U702 ( .A(n630), .B(G110), .ZN(G12) );
  XNOR2_X1 U703 ( .A(G119), .B(KEYINPUT127), .ZN(n632) );
  XOR2_X1 U704 ( .A(n632), .B(n631), .Z(G21) );
  XNOR2_X1 U705 ( .A(n633), .B(KEYINPUT126), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(G24) );
  NOR2_X1 U707 ( .A1(n731), .A2(n636), .ZN(n639) );
  XNOR2_X1 U708 ( .A(n637), .B(KEYINPUT62), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U710 ( .A1(n640), .A2(n738), .ZN(n642) );
  XNOR2_X1 U711 ( .A(KEYINPUT95), .B(KEYINPUT63), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(G57) );
  XOR2_X1 U713 ( .A(G101), .B(n643), .Z(G3) );
  XOR2_X1 U714 ( .A(G104), .B(KEYINPUT111), .Z(n645) );
  NAND2_X1 U715 ( .A1(n646), .A2(n364), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n648) );
  NAND2_X1 U718 ( .A1(n646), .A2(n658), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U720 ( .A(G107), .B(n649), .ZN(G9) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .Z(n652) );
  NAND2_X1 U722 ( .A1(n654), .A2(n658), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(G30) );
  XNOR2_X1 U724 ( .A(G143), .B(n653), .ZN(G45) );
  NAND2_X1 U725 ( .A1(n654), .A2(n364), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n655), .B(KEYINPUT112), .ZN(n656) );
  XNOR2_X1 U727 ( .A(G146), .B(n656), .ZN(G48) );
  NAND2_X1 U728 ( .A1(n659), .A2(n364), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(G113), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n660), .B(G116), .ZN(G18) );
  XOR2_X1 U732 ( .A(G125), .B(KEYINPUT37), .Z(n661) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(G27) );
  NOR2_X1 U734 ( .A1(n690), .A2(n663), .ZN(n664) );
  NOR2_X1 U735 ( .A1(n664), .A2(G953), .ZN(n673) );
  NOR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n671) );
  INV_X1 U737 ( .A(n667), .ZN(n669) );
  XNOR2_X1 U738 ( .A(KEYINPUT87), .B(KEYINPUT2), .ZN(n668) );
  NOR2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n707) );
  INV_X1 U742 ( .A(n674), .ZN(n686) );
  NAND2_X1 U743 ( .A1(n544), .A2(n675), .ZN(n677) );
  XOR2_X1 U744 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n676) );
  XNOR2_X1 U745 ( .A(n677), .B(n676), .ZN(n684) );
  NAND2_X1 U746 ( .A1(n679), .A2(n359), .ZN(n680) );
  XNOR2_X1 U747 ( .A(KEYINPUT50), .B(n680), .ZN(n682) );
  NAND2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U751 ( .A(n687), .B(KEYINPUT114), .Z(n688) );
  XNOR2_X1 U752 ( .A(KEYINPUT51), .B(n688), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U758 ( .A1(n663), .A2(n699), .ZN(n700) );
  NOR2_X1 U759 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U760 ( .A(n702), .B(KEYINPUT115), .Z(n703) );
  XNOR2_X1 U761 ( .A(KEYINPUT52), .B(n703), .ZN(n704) );
  NOR2_X1 U762 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U763 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n708), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U765 ( .A1(n731), .A2(n709), .ZN(n715) );
  XOR2_X1 U766 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n711) );
  XNOR2_X1 U767 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n710) );
  XNOR2_X1 U768 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U769 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U770 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n738), .A2(n716), .ZN(n717) );
  XNOR2_X1 U772 ( .A(KEYINPUT118), .B(n717), .ZN(G54) );
  NOR2_X1 U773 ( .A1(n731), .A2(n718), .ZN(n723) );
  XNOR2_X1 U774 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n721) );
  XNOR2_X1 U775 ( .A(n719), .B(KEYINPUT97), .ZN(n720) );
  XNOR2_X1 U776 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n738), .A2(n724), .ZN(n725) );
  XNOR2_X1 U779 ( .A(KEYINPUT60), .B(n725), .ZN(G60) );
  NAND2_X1 U780 ( .A1(n726), .A2(G478), .ZN(n729) );
  NOR2_X1 U781 ( .A1(n738), .A2(n730), .ZN(G63) );
  BUF_X1 U782 ( .A(n731), .Z(n733) );
  NOR2_X1 U783 ( .A1(n733), .A2(n732), .ZN(n736) );
  XNOR2_X1 U784 ( .A(n734), .B(KEYINPUT121), .ZN(n735) );
  XNOR2_X1 U785 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U786 ( .A1(n738), .A2(n737), .ZN(G66) );
  NAND2_X1 U787 ( .A1(n618), .A2(n754), .ZN(n742) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n739) );
  XNOR2_X1 U789 ( .A(KEYINPUT61), .B(n739), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n740), .A2(G898), .ZN(n741) );
  NAND2_X1 U791 ( .A1(n742), .A2(n741), .ZN(n747) );
  XOR2_X1 U792 ( .A(n743), .B(G110), .Z(n745) );
  NOR2_X1 U793 ( .A1(n754), .A2(G898), .ZN(n744) );
  NOR2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U795 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U796 ( .A(KEYINPUT122), .B(n748), .ZN(G69) );
  XNOR2_X1 U797 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n749) );
  XNOR2_X1 U798 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(n756) );
  XNOR2_X1 U800 ( .A(n756), .B(n753), .ZN(n755) );
  NAND2_X1 U801 ( .A1(n755), .A2(n754), .ZN(n761) );
  XNOR2_X1 U802 ( .A(n756), .B(G227), .ZN(n757) );
  XNOR2_X1 U803 ( .A(n757), .B(KEYINPUT125), .ZN(n758) );
  NAND2_X1 U804 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U805 ( .A1(n759), .A2(G953), .ZN(n760) );
  NAND2_X1 U806 ( .A1(n761), .A2(n760), .ZN(G72) );
  XOR2_X1 U807 ( .A(G131), .B(n762), .Z(G33) );
  XNOR2_X1 U808 ( .A(G134), .B(n763), .ZN(G36) );
  XOR2_X1 U809 ( .A(G137), .B(n764), .Z(G39) );
endmodule

