//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT64), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n460), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT64), .B(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n459), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(G160));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n466), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n459), .B1(new_n467), .B2(new_n458), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(KEYINPUT65), .ZN(new_n481));
  OAI21_X1  g056(.A(G2105), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n482), .A2(KEYINPUT66), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(KEYINPUT66), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT67), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n479), .A2(new_n481), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(new_n491), .B2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT68), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n459), .B(new_n496), .C1(new_n467), .C2(new_n458), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n500), .A2(KEYINPUT69), .A3(new_n459), .A4(new_n496), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n473), .A2(new_n503), .A3(new_n496), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n470), .A2(G102), .A3(G2104), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G126), .ZN(new_n508));
  INV_X1    g083(.A(G114), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n480), .A2(new_n508), .B1(new_n509), .B2(new_n461), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n510), .B2(G2105), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G62), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(KEYINPUT70), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n519), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n523), .A2(new_n529), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT6), .B(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n532), .A2(new_n534), .A3(G543), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n533), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n516), .A2(new_n518), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT7), .Z(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G168));
  AND2_X1   g120(.A1(new_n536), .A2(G52), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n519), .A2(new_n533), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n547), .A2(new_n514), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n546), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n552), .A2(new_n514), .B1(new_n553), .B2(new_n549), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(G43), .B2(new_n536), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  XOR2_X1   g133(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n536), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(new_n549), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n539), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n565), .A2(G91), .B1(G651), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n564), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  XNOR2_X1  g146(.A(new_n544), .B(KEYINPUT73), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  NAND2_X1  g149(.A1(new_n536), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n565), .A2(G87), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT74), .Z(new_n581));
  AND3_X1   g156(.A1(new_n516), .A2(new_n518), .A3(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G48), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n539), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(new_n533), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n565), .A2(G85), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(KEYINPUT75), .B(G47), .ZN(new_n591));
  OAI221_X1 g166(.A(new_n589), .B1(new_n514), .B2(new_n590), .C1(new_n535), .C2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n535), .B2(KEYINPUT76), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(KEYINPUT76), .B2(new_n535), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n565), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n549), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n539), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n596), .A2(new_n599), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n611), .B2(KEYINPUT77), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(KEYINPUT77), .B2(new_n609), .ZN(G297));
  XOR2_X1   g188(.A(G297), .B(KEYINPUT78), .Z(G280));
  INV_X1    g189(.A(new_n604), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  OR2_X1    g192(.A1(new_n555), .A2(G868), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n604), .A2(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n485), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n491), .A2(G135), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n470), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n467), .A2(new_n470), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(new_n472), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n631), .A2(new_n632), .B1(new_n633), .B2(G2100), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n632), .B2(new_n631), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n633), .A2(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n627), .A2(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(G2427), .B(G2430), .Z(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT80), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(KEYINPUT17), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n658), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n662), .B(new_n664), .C1(new_n665), .C2(new_n661), .ZN(new_n666));
  OR3_X1    g241(.A1(new_n664), .A2(KEYINPUT18), .A3(new_n660), .ZN(new_n667));
  OAI21_X1  g242(.A(KEYINPUT18), .B1(new_n664), .B2(new_n660), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT82), .B(G2096), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n676), .B1(new_n682), .B2(KEYINPUT84), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(KEYINPUT84), .B2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n677), .A2(new_n679), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n676), .B2(new_n681), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n676), .A2(KEYINPUT85), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT86), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n690), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(KEYINPUT99), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  MUX2_X1   g276(.A(new_n700), .B(new_n701), .S(KEYINPUT91), .Z(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G1971), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n578), .A2(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G16), .B2(G23), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n699), .A2(G6), .ZN(new_n709));
  INV_X1    g284(.A(G305), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n699), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT32), .B(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT90), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n711), .B(new_n713), .Z(new_n714));
  NOR3_X1   g289(.A1(new_n707), .A2(new_n708), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n702), .A2(G1971), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n703), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT89), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT34), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n485), .A2(G119), .ZN(new_n723));
  OR3_X1    g298(.A1(KEYINPUT87), .A2(G95), .A3(G2105), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(new_n470), .B2(G107), .ZN(new_n725));
  OR2_X1    g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(KEYINPUT87), .B2(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n491), .A2(G131), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT88), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n723), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n722), .B1(new_n734), .B2(new_n721), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT35), .B(G1991), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G24), .B(G290), .S(G16), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1986), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n719), .A2(new_n720), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n720), .B1(new_n719), .B2(new_n740), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G162), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G35), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(KEYINPUT29), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n747), .A2(G2090), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT97), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n721), .A2(G33), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT25), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n491), .B2(G139), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n473), .A2(G127), .ZN(new_n756));
  NAND2_X1  g331(.A1(G115), .A2(G2104), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n470), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(new_n721), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G2072), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n491), .A2(G141), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  INV_X1    g339(.A(G105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n765), .C2(new_n628), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G129), .B2(new_n485), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G29), .B2(G32), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT24), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G160), .B2(new_n721), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n769), .A2(new_n770), .B1(G2084), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n761), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT94), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n721), .A2(G26), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n485), .A2(G128), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n781));
  INV_X1    g356(.A(G116), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G2105), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n491), .B2(G140), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(new_n721), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n779), .B(new_n787), .S(KEYINPUT28), .Z(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n699), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT23), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n610), .B2(new_n699), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G27), .A2(G29), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G164), .B2(G29), .ZN(new_n798));
  INV_X1    g373(.A(G2078), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n615), .A2(G16), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G4), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1348), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G1961), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n699), .A2(G5), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G171), .B2(new_n699), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT96), .Z(new_n808));
  AOI21_X1  g383(.A(new_n804), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n805), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n769), .A2(new_n770), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n555), .A2(new_n699), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n699), .B2(G19), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT92), .B(G1341), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT31), .B(G11), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT30), .B(G28), .Z(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G29), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n813), .B2(new_n814), .ZN(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G21), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G168), .B2(G16), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT95), .B(G1966), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n775), .A2(G2084), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n815), .A2(new_n819), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n802), .A2(new_n803), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n626), .B2(new_n721), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n810), .A2(new_n811), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n790), .A2(new_n796), .A3(new_n800), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(G2090), .B1(new_n747), .B2(new_n748), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n750), .A2(new_n778), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n698), .B1(new_n744), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n743), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n741), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n778), .A2(new_n831), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n835), .A2(KEYINPUT99), .A3(new_n750), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n837), .ZN(G311));
  NAND3_X1  g413(.A1(new_n835), .A2(new_n750), .A3(new_n836), .ZN(G150));
  INV_X1    g414(.A(G55), .ZN(new_n840));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n535), .A2(new_n840), .B1(new_n841), .B2(new_n549), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT101), .ZN(new_n843));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n539), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n847));
  OAI21_X1  g422(.A(G651), .B1(new_n846), .B2(KEYINPUT100), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(KEYINPUT102), .B2(new_n555), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n555), .A2(KEYINPUT102), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT103), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n615), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n849), .A2(G860), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT104), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(G145));
  NOR2_X1   g440(.A1(new_n785), .A2(new_n512), .ZN(new_n866));
  AOI21_X1  g441(.A(G164), .B1(new_n780), .B2(new_n784), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n755), .A2(new_n758), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n759), .B1(new_n866), .B2(new_n867), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(new_n767), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n767), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n485), .A2(G130), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  INV_X1    g450(.A(G118), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(G2105), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(new_n491), .B2(G142), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n631), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(new_n631), .A3(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n733), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n880), .A2(new_n730), .A3(new_n732), .A4(new_n881), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT105), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT105), .B1(new_n883), .B2(new_n884), .ZN(new_n887));
  OAI22_X1  g462(.A1(new_n872), .A2(new_n873), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n870), .A2(new_n871), .ZN(new_n890));
  INV_X1    g465(.A(new_n767), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n870), .A2(new_n871), .A3(new_n767), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n889), .A2(new_n892), .A3(new_n893), .A4(new_n885), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n626), .B(G160), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G162), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n872), .B2(new_n873), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n901));
  INV_X1    g476(.A(new_n883), .ZN(new_n902));
  INV_X1    g477(.A(new_n884), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n897), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n888), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n888), .A2(new_n906), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT107), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n898), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g489(.A1(new_n849), .A2(new_n605), .ZN(new_n915));
  XNOR2_X1  g490(.A(G299), .B(new_n615), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT41), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n916), .B(KEYINPUT108), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n855), .B(new_n619), .ZN(new_n919));
  MUX2_X1   g494(.A(new_n917), .B(new_n918), .S(new_n919), .Z(new_n920));
  XNOR2_X1  g495(.A(G166), .B(G305), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n578), .B(G290), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n921), .B(new_n922), .Z(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n920), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n915), .B1(new_n925), .B2(new_n605), .ZN(G295));
  OAI21_X1  g501(.A(new_n915), .B1(new_n925), .B2(new_n605), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n928));
  NOR2_X1   g503(.A1(G171), .A2(new_n544), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(G286), .B2(G171), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n853), .A2(new_n854), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n853), .B2(new_n854), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n928), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n917), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n932), .A2(new_n933), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n938), .A2(new_n916), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n923), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n916), .ZN(new_n941));
  INV_X1    g516(.A(new_n923), .ZN(new_n942));
  INV_X1    g517(.A(new_n933), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n931), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n935), .B1(new_n944), .B2(new_n928), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n941), .B(new_n942), .C1(new_n945), .C2(new_n917), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  AOI211_X1 g524(.A(new_n918), .B(new_n935), .C1(new_n944), .C2(new_n928), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n938), .A2(new_n917), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n923), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n947), .A3(new_n946), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n953), .B2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n953), .B2(KEYINPUT43), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n957), .A2(KEYINPUT110), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT110), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G397));
  INV_X1    g536(.A(new_n476), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT111), .B(G40), .Z(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n962), .B(new_n964), .C1(new_n468), .C2(G2105), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  INV_X1    g541(.A(new_n504), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n503), .B1(new_n497), .B2(new_n498), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n501), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n509), .A2(new_n461), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n466), .B2(G126), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n506), .B1(new_n971), .B2(new_n470), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n966), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT45), .B(new_n966), .C1(new_n969), .C2(new_n972), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT56), .B(G2072), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT120), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n981), .B(new_n966), .C1(new_n969), .C2(new_n972), .ZN(new_n982));
  INV_X1    g557(.A(new_n965), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n977), .A2(new_n979), .B1(new_n984), .B2(new_n795), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n986));
  XOR2_X1   g561(.A(G299), .B(new_n986), .Z(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n505), .B2(new_n511), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n984), .A2(new_n803), .B1(new_n991), .B2(new_n789), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(new_n604), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n985), .A2(new_n987), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n988), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n985), .A2(new_n987), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(KEYINPUT61), .A3(new_n994), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT61), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n985), .A2(new_n987), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n999), .B2(new_n988), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT60), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n992), .B(new_n615), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n997), .B(new_n1000), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n973), .A2(new_n974), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n983), .A3(new_n976), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT58), .B(G1341), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n1005), .A2(G1996), .B1(new_n991), .B2(new_n1006), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1007), .A2(new_n555), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1008), .A2(KEYINPUT59), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(KEYINPUT59), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n992), .A2(new_n1001), .A3(new_n615), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n995), .B1(new_n1003), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT125), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1005), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n975), .A2(KEYINPUT113), .A3(new_n976), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n799), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1020), .A2(new_n1021), .B1(new_n805), .B2(new_n984), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n1005), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(G171), .B(KEYINPUT54), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n976), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1004), .A2(G40), .A3(G160), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1029), .B(new_n1023), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1027), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1022), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G166), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT55), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1971), .ZN(new_n1041));
  AND4_X1   g616(.A1(KEYINPUT113), .A2(new_n1004), .A3(new_n983), .A4(new_n976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT113), .B1(new_n975), .B2(new_n976), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n983), .B1(new_n989), .B2(new_n981), .ZN(new_n1046));
  INV_X1    g621(.A(new_n982), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT114), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G2090), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n965), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n982), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1044), .A2(new_n1045), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G8), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1045), .B1(new_n1044), .B2(new_n1053), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1040), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1971), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n984), .A2(G2090), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1039), .B(G8), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n991), .A2(new_n1037), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n578), .A2(G1976), .ZN(new_n1062));
  INV_X1    g637(.A(G1976), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(G288), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n990), .A2(G8), .A3(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1067));
  XNOR2_X1  g642(.A(G305), .B(G1981), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(KEYINPUT49), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1065), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1060), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1057), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT115), .B1(new_n1077), .B2(new_n1058), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(G8), .A3(new_n1054), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1072), .B1(new_n1079), .B2(new_n1040), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT124), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1036), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT116), .B1(new_n984), .B2(G2084), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n1084));
  INV_X1    g659(.A(G2084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1050), .A2(new_n1084), .A3(new_n1085), .A4(new_n982), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1005), .A2(new_n822), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(G8), .A3(new_n544), .ZN(new_n1089));
  OAI21_X1  g664(.A(G8), .B1(new_n1088), .B2(new_n544), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT51), .B(G8), .C1(new_n1088), .C2(new_n544), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1091), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1089), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1016), .B1(new_n1082), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1036), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1057), .A2(KEYINPUT124), .A3(new_n1073), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT124), .B1(new_n1057), .B2(new_n1073), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1097), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(KEYINPUT125), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1015), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1060), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1070), .A2(new_n1063), .A3(new_n578), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(G1981), .B2(G305), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1105), .A2(new_n1071), .B1(new_n1107), .B2(new_n1061), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1088), .A2(G8), .A3(new_n572), .ZN(new_n1109));
  OAI21_X1  g684(.A(G8), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1040), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1073), .A2(KEYINPUT63), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT63), .B1(new_n1080), .B2(new_n1109), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g690(.A(KEYINPUT117), .B(KEYINPUT63), .C1(new_n1080), .C2(new_n1109), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1108), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT118), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1097), .A2(KEYINPUT62), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1076), .A2(new_n1081), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1097), .A2(KEYINPUT62), .ZN(new_n1121));
  AOI21_X1  g696(.A(G301), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1124), .B(new_n1108), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1104), .A2(new_n1118), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n767), .B(G1996), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1004), .A2(new_n965), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n785), .B(new_n789), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(new_n1129), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(KEYINPUT112), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(KEYINPUT112), .B2(new_n1132), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n733), .A2(new_n736), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n733), .A2(new_n736), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1129), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(G290), .B(G1986), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1128), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1126), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT46), .ZN(new_n1142));
  OR3_X1    g717(.A1(new_n1129), .A2(new_n1142), .A3(G1996), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1142), .B1(new_n1129), .B2(G1996), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1131), .A2(new_n767), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1143), .B(new_n1144), .C1(new_n1145), .C2(new_n1129), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT126), .Z(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT47), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n786), .A2(new_n789), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1129), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1129), .A2(G1986), .A3(G290), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT48), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1138), .A2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1148), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1141), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g731(.A(G229), .ZN(new_n1158));
  NAND3_X1  g732(.A1(new_n1158), .A2(new_n672), .A3(G319), .ZN(new_n1159));
  NOR2_X1   g733(.A1(G401), .A2(new_n1159), .ZN(new_n1160));
  AND4_X1   g734(.A1(KEYINPUT127), .A2(new_n954), .A3(new_n913), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1162));
  OAI21_X1  g736(.A(new_n908), .B1(new_n905), .B2(new_n907), .ZN(new_n1163));
  NAND3_X1  g737(.A1(new_n910), .A2(KEYINPUT107), .A3(new_n911), .ZN(new_n1164));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g739(.A(new_n1162), .B1(new_n1165), .B2(new_n898), .ZN(new_n1166));
  AOI21_X1  g740(.A(KEYINPUT127), .B1(new_n1166), .B2(new_n954), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n1161), .A2(new_n1167), .ZN(G308));
  NAND3_X1  g742(.A1(new_n954), .A2(new_n913), .A3(new_n1160), .ZN(new_n1169));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n1166), .A2(KEYINPUT127), .A3(new_n954), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1172), .ZN(G225));
endmodule


