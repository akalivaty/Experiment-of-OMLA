//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g0008(.A(G250), .B1(G257), .B2(G264), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n210), .A2(KEYINPUT0), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n216), .B1(KEYINPUT0), .B2(new_n210), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n212), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  AND2_X1   g0049(.A1(G58), .A2(G68), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G58), .A2(G68), .ZN(new_n251));
  OAI21_X1  g0051(.A(G20), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G159), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n204), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n218), .B1(new_n258), .B2(KEYINPUT7), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT7), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n211), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n255), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n249), .B1(new_n265), .B2(KEYINPUT16), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT16), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(new_n262), .B2(new_n211), .ZN(new_n268));
  NOR4_X1   g0068(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT7), .A4(G20), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n268), .A2(new_n269), .A3(new_n218), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n270), .B2(new_n255), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n203), .B2(G20), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n248), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n274), .A2(new_n277), .B1(new_n273), .B2(new_n276), .ZN(new_n278));
  INV_X1    g0078(.A(G200), .ZN(new_n279));
  OR2_X1    g0079(.A1(G223), .A2(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G226), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G1698), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n280), .B(new_n282), .C1(new_n260), .C2(new_n261), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G87), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n292), .A3(G274), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(G232), .A3(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n279), .B1(new_n287), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n292), .B1(new_n283), .B2(new_n284), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n272), .A2(KEYINPUT76), .A3(new_n278), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT17), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n278), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n266), .B2(new_n271), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n307), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n302), .ZN(new_n308));
  INV_X1    g0108(.A(new_n255), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n260), .A2(new_n261), .A3(G20), .ZN(new_n310));
  OAI21_X1  g0110(.A(G68), .B1(new_n310), .B2(new_n263), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n262), .A2(new_n211), .A3(new_n263), .ZN(new_n312));
  OAI211_X1 g0112(.A(KEYINPUT16), .B(new_n309), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n248), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n256), .A2(new_n257), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT64), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT7), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n310), .A2(new_n263), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(G68), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT16), .B1(new_n322), .B2(new_n309), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n278), .B1(new_n314), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n298), .A2(new_n299), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n298), .A2(new_n299), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT75), .A2(KEYINPUT18), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT75), .A2(KEYINPUT18), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n324), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n329), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n326), .B1(new_n335), .B2(G169), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n331), .B1(new_n307), .B2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n305), .A2(new_n308), .A3(new_n334), .A4(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n276), .A2(new_n218), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT12), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n203), .A2(G20), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n277), .A2(G68), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT74), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(KEYINPUT74), .A3(new_n343), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n211), .A2(G33), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n220), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n248), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n346), .A2(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  INV_X1    g0156(.A(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n281), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G232), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n358), .B(new_n360), .C1(new_n260), .C2(new_n261), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n292), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(KEYINPUT73), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n292), .A2(new_n294), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n293), .B1(new_n219), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n356), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g0171(.A(KEYINPUT13), .B(new_n369), .C1(new_n365), .C2(new_n366), .ZN(new_n372));
  OAI21_X1  g0172(.A(G169), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n373), .A2(KEYINPUT14), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT14), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(G169), .C1(new_n371), .C2(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n367), .A2(new_n370), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n367), .A2(new_n356), .A3(new_n370), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(G179), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n355), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(G190), .A3(new_n379), .ZN(new_n383));
  OAI21_X1  g0183(.A(G200), .B1(new_n371), .B2(new_n372), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(new_n354), .ZN(new_n385));
  INV_X1    g0185(.A(new_n253), .ZN(new_n386));
  XOR2_X1   g0186(.A(KEYINPUT8), .B(G58), .Z(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT70), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT70), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n273), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n386), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n349), .A2(new_n392), .B1(new_n220), .B2(new_n211), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n248), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n342), .A2(G77), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n277), .A2(new_n396), .B1(new_n220), .B2(new_n276), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT71), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n394), .A2(new_n400), .A3(new_n397), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(G232), .A2(G1698), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n357), .A2(G238), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n315), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n286), .C1(G107), .C2(new_n315), .ZN(new_n406));
  INV_X1    g0206(.A(new_n368), .ZN(new_n407));
  INV_X1    g0207(.A(G274), .ZN(new_n408));
  INV_X1    g0208(.A(new_n212), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(new_n291), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n407), .A2(G244), .B1(new_n290), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(G179), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n328), .B2(new_n412), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n402), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n402), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT69), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n412), .B2(new_n300), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n406), .A2(new_n411), .A3(KEYINPUT69), .A4(G190), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n418), .A2(new_n419), .B1(G200), .B2(new_n412), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n415), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n339), .A2(new_n382), .A3(new_n385), .A4(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT68), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n315), .A2(KEYINPUT67), .A3(G222), .A4(new_n357), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT67), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n357), .A2(G222), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n262), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n357), .B1(new_n256), .B2(new_n257), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(G223), .B1(new_n262), .B2(G77), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n286), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n293), .B1(new_n281), .B2(new_n368), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n423), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n292), .B1(new_n428), .B2(new_n430), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n436), .A2(KEYINPUT68), .A3(new_n433), .ZN(new_n437));
  OAI21_X1  g0237(.A(G190), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n432), .A2(new_n423), .A3(new_n434), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT68), .B1(new_n436), .B2(new_n433), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(G200), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G50), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n203), .B2(G20), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n277), .A2(new_n443), .B1(new_n442), .B2(new_n276), .ZN(new_n444));
  INV_X1    g0244(.A(G33), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n319), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n387), .ZN(new_n447));
  INV_X1    g0247(.A(G58), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(new_n448), .A3(new_n218), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(G20), .B1(G150), .B2(new_n253), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT9), .B(new_n444), .C1(new_n451), .C2(new_n249), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT9), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n249), .B1(new_n447), .B2(new_n450), .ZN(new_n454));
  INV_X1    g0254(.A(new_n444), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n438), .A2(new_n441), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT72), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n438), .A2(new_n460), .A3(new_n458), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT10), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n439), .A2(new_n440), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n457), .B1(new_n464), .B2(G190), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n441), .C1(new_n460), .C2(KEYINPUT10), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n454), .A2(new_n455), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n464), .B2(new_n325), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G169), .B2(new_n464), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n463), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n422), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT78), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT78), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(G33), .A3(G283), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n357), .A2(G244), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n256), .B2(new_n257), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n478), .B2(KEYINPUT4), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n221), .A2(G1698), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(KEYINPUT4), .C1(new_n261), .C2(new_n260), .ZN(new_n481));
  OAI211_X1 g0281(.A(G250), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n286), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n289), .A2(G1), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G257), .A3(new_n292), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n203), .A2(G45), .ZN(new_n491));
  OR2_X1    g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n486), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n410), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n484), .A2(new_n300), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n490), .A2(new_n494), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n262), .B2(new_n477), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(new_n476), .A3(new_n481), .A4(new_n482), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n500), .B2(new_n286), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n496), .B1(new_n501), .B2(G200), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT77), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n320), .A2(new_n321), .A3(G107), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  AND2_X1   g0305(.A1(G97), .A2(G107), .ZN(new_n506));
  NOR2_X1   g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(KEYINPUT6), .A3(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(new_n319), .B1(G77), .B2(new_n253), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n249), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n275), .A2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n203), .A2(G33), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n275), .A2(new_n515), .A3(new_n212), .A4(new_n247), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n517), .B2(G97), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n503), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n268), .A2(new_n269), .A3(new_n509), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n509), .A2(KEYINPUT6), .A3(G97), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n505), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n524), .A2(new_n211), .B1(new_n220), .B2(new_n386), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n248), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(KEYINPUT77), .A3(new_n518), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n502), .A2(new_n520), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n502), .A2(new_n520), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n501), .A2(G179), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n328), .B2(new_n501), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT80), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n513), .B2(new_n519), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n526), .A2(KEYINPUT80), .A3(new_n518), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n529), .A2(new_n531), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n493), .A2(new_n286), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n539), .A2(G270), .B1(new_n410), .B2(new_n493), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(new_n357), .C1(new_n260), .C2(new_n261), .ZN(new_n541));
  OAI211_X1 g0341(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n542));
  INV_X1    g0342(.A(G303), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n315), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n286), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n328), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n275), .A2(G116), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n517), .B2(G116), .ZN(new_n548));
  INV_X1    g0348(.A(G116), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n247), .A2(new_n212), .B1(G20), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n473), .A2(new_n475), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n445), .A2(G97), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n316), .A2(new_n318), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT20), .B(new_n550), .C1(new_n551), .C2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n476), .A2(new_n211), .A3(new_n552), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT20), .B1(new_n556), .B2(new_n550), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n548), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n546), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n540), .A2(new_n545), .A3(G179), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n559), .A2(new_n560), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n546), .A2(new_n558), .A3(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n540), .A2(new_n545), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n279), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n565), .A2(new_n300), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n567), .A2(new_n558), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n315), .A2(G257), .A3(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n315), .A2(G250), .A3(new_n357), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G294), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n286), .B1(G264), .B2(new_n539), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n325), .A3(new_n494), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n494), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n328), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n316), .B(new_n318), .C1(new_n260), .C2(new_n261), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT22), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n315), .A2(new_n211), .A3(new_n582), .A4(G87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT23), .B1(new_n204), .B2(G107), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G116), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(G20), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(KEYINPUT23), .A2(G107), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n319), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT24), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT24), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n584), .A2(new_n592), .A3(new_n589), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n249), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G13), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(G1), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(G20), .A3(new_n509), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT25), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n516), .A2(new_n509), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n576), .B(new_n578), .C1(new_n594), .C2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G250), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n491), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n203), .A2(new_n408), .A3(G45), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n292), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n219), .A2(new_n357), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n221), .A2(G1698), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n260), .C2(new_n261), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(new_n586), .ZN(new_n610));
  OAI211_X1 g0410(.A(G179), .B(new_n606), .C1(new_n610), .C2(new_n292), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n292), .B1(new_n609), .B2(new_n586), .ZN(new_n612));
  INV_X1    g0412(.A(new_n606), .ZN(new_n613));
  OAI21_X1  g0413(.A(G169), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n316), .A2(new_n318), .A3(G33), .A4(G97), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n315), .A2(new_n211), .A3(G68), .ZN(new_n619));
  NAND3_X1  g0419(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n316), .A2(new_n318), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n507), .A2(new_n580), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n618), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n248), .B1(new_n276), .B2(new_n392), .ZN(new_n625));
  INV_X1    g0425(.A(new_n392), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n517), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n615), .A2(KEYINPUT81), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT81), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n611), .A2(new_n614), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n612), .A2(new_n613), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT82), .B1(new_n631), .B2(G190), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT82), .ZN(new_n633));
  NOR4_X1   g0433(.A1(new_n612), .A2(new_n613), .A3(new_n633), .A4(new_n300), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n624), .A2(new_n248), .ZN(new_n636));
  OAI21_X1  g0436(.A(G200), .B1(new_n612), .B2(new_n613), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n392), .A2(new_n276), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n517), .A2(G87), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n628), .A2(new_n630), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n593), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n592), .B1(new_n584), .B2(new_n589), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n248), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n577), .A2(G200), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n575), .A2(G190), .A3(new_n494), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n600), .A4(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n602), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n471), .A2(new_n538), .A3(new_n570), .A4(new_n649), .ZN(G372));
  NAND2_X1  g0450(.A1(new_n305), .A2(new_n308), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n415), .A2(new_n385), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n382), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT85), .B1(new_n307), .B2(new_n336), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT85), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n324), .A2(new_n655), .A3(new_n330), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n654), .A2(KEYINPUT18), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT18), .B1(new_n654), .B2(new_n656), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n466), .B(new_n463), .C1(new_n653), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n469), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n625), .A2(new_n627), .B1(new_n611), .B2(new_n614), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT83), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n640), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n631), .A2(G190), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n625), .A2(KEYINPUT83), .A3(new_n637), .A4(new_n639), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n663), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT84), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT84), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(new_n671), .A3(new_n663), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n591), .A2(new_n593), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n601), .B1(new_n674), .B2(new_n248), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n578), .A2(new_n576), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n562), .B(new_n563), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n673), .A2(new_n538), .A3(new_n648), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n520), .A2(new_n527), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n533), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT26), .B1(new_n673), .B2(new_n681), .ZN(new_n682));
  AND4_X1   g0482(.A1(KEYINPUT26), .A2(new_n642), .A3(new_n533), .A4(new_n537), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n663), .B(new_n678), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n661), .B1(new_n471), .B2(new_n684), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT86), .Z(G369));
  NAND2_X1  g0486(.A1(new_n211), .A2(new_n596), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  OAI21_X1  g0488(.A(G213), .B1(new_n687), .B2(KEYINPUT27), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G343), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n692), .A2(new_n558), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n564), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n695));
  INV_X1    g0495(.A(new_n570), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n693), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n694), .A2(KEYINPUT87), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n602), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n692), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n602), .B(new_n648), .C1(new_n675), .C2(new_n691), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n699), .A2(G330), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n564), .A2(new_n602), .A3(new_n648), .A4(new_n691), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n691), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n709), .ZN(G399));
  NOR2_X1   g0510(.A1(new_n208), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n622), .A2(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n214), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT89), .B1(new_n684), .B2(new_n691), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n529), .A2(new_n531), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n537), .A2(new_n533), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n677), .A3(new_n720), .A4(new_n648), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n640), .A2(new_n664), .B1(G190), .B2(new_n631), .ZN(new_n722));
  AOI211_X1 g0522(.A(KEYINPUT84), .B(new_n662), .C1(new_n722), .C2(new_n667), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n671), .B1(new_n668), .B2(new_n663), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n663), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n681), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT26), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n683), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI211_X1 g0529(.A(KEYINPUT89), .B(new_n691), .C1(new_n726), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n717), .B1(new_n718), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n642), .A2(new_n728), .A3(new_n533), .A4(new_n537), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n678), .A2(new_n663), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n728), .B1(new_n673), .B2(new_n681), .ZN(new_n735));
  OAI211_X1 g0535(.A(KEYINPUT29), .B(new_n691), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n575), .A2(new_n631), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n484), .A2(new_n495), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n325), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n738), .A2(new_n740), .A3(KEYINPUT30), .A4(new_n566), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n501), .A2(G179), .A3(new_n631), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n565), .A3(new_n577), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n575), .A2(new_n545), .A3(new_n540), .A4(new_n631), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(new_n532), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT88), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n649), .A2(new_n538), .A3(new_n570), .A4(new_n691), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n747), .B2(new_n692), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n748), .A2(KEYINPUT88), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n749), .A2(new_n750), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G330), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n737), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n716), .B1(new_n756), .B2(G1), .ZN(G364));
  NOR2_X1   g0557(.A1(new_n319), .A2(new_n595), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n203), .B1(new_n758), .B2(G45), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n712), .A2(KEYINPUT90), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT90), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(new_n711), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n699), .B2(G330), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G330), .B2(new_n699), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT91), .Z(new_n768));
  AOI21_X1  g0568(.A(new_n212), .B1(G20), .B2(new_n328), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n204), .A2(new_n300), .A3(new_n279), .A4(G179), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G87), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n319), .A2(new_n325), .A3(new_n300), .A4(G200), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n315), .C1(new_n509), .C2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n319), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G159), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n300), .A2(G200), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n211), .B1(new_n325), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n774), .B(new_n779), .C1(G97), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n211), .A2(new_n325), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(new_n300), .A3(new_n279), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(KEYINPUT94), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n784), .A2(new_n780), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT93), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n789), .A2(G77), .B1(G58), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n784), .A2(new_n300), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G50), .A2(new_n794), .B1(new_n796), .B2(G68), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n783), .A2(new_n792), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  INV_X1    g0599(.A(new_n771), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n262), .B1(new_n773), .B2(new_n799), .C1(new_n543), .C2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G329), .B2(new_n777), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n785), .A2(new_n803), .B1(new_n790), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G294), .B2(new_n782), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n796), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n794), .A2(G326), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n802), .A2(new_n806), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n770), .B1(new_n798), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n242), .A2(G45), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n208), .A2(new_n315), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G45), .C2(new_n214), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n208), .A2(new_n262), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G355), .B1(new_n549), .B2(new_n208), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT92), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n822), .B(new_n769), .C1(new_n818), .C2(KEYINPUT92), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n764), .B(new_n811), .C1(new_n819), .C2(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT95), .Z(new_n825));
  NOR2_X1   g0625(.A1(new_n697), .A2(new_n698), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n822), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n768), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  AND2_X1   g0630(.A1(new_n421), .A2(new_n691), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n726), .B2(new_n729), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n718), .A2(new_n731), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n415), .A2(new_n691), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n691), .B1(new_n399), .B2(new_n401), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n416), .B2(new_n420), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n834), .B1(new_n836), .B2(new_n415), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT98), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n832), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n765), .B1(new_n839), .B2(new_n755), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n755), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n769), .A2(new_n820), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n791), .A2(G143), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G137), .A2(new_n794), .B1(new_n796), .B2(G150), .ZN(new_n845));
  INV_X1    g0645(.A(new_n789), .ZN(new_n846));
  INV_X1    g0646(.A(G159), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n849));
  OR2_X1    g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  INV_X1    g0651(.A(new_n773), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(G68), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n777), .A2(G132), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n262), .B1(new_n771), .B2(G50), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G58), .B2(new_n782), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n850), .A2(new_n851), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n789), .A2(G116), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n773), .A2(new_n580), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n262), .B1(new_n800), .B2(new_n509), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n860), .B(new_n861), .C1(G311), .C2(new_n777), .ZN(new_n862));
  INV_X1    g0662(.A(new_n790), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n863), .A2(G294), .B1(new_n782), .B2(G97), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G283), .A2(new_n796), .B1(new_n794), .B2(G303), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n859), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n765), .B1(G77), .B2(new_n843), .C1(new_n867), .C2(new_n770), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT97), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  INV_X1    g0671(.A(new_n837), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n870), .B(new_n871), .C1(new_n821), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n841), .A2(new_n873), .ZN(G384));
  OR2_X1    g0674(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(new_n876), .A3(G116), .A4(new_n213), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT36), .Z(new_n878));
  OAI211_X1 g0678(.A(new_n215), .B(G77), .C1(new_n448), .C2(new_n218), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n442), .A2(G68), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n203), .B(G13), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n267), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n306), .B1(new_n266), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n690), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n338), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n302), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n324), .A2(new_n889), .B1(new_n885), .B2(new_n886), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n885), .A2(new_n336), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n307), .A2(new_n302), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n324), .A2(new_n330), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n324), .A2(new_n690), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n888), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n888), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(KEYINPUT100), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT100), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n899), .A2(new_n905), .A3(new_n900), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n355), .A2(new_n692), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n382), .A2(new_n385), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n373), .A2(KEYINPUT14), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n380), .A3(new_n376), .ZN(new_n912));
  INV_X1    g0712(.A(new_n385), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n355), .B(new_n692), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT99), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n832), .A2(new_n916), .A3(new_n834), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n832), .B2(new_n834), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n908), .B(new_n915), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n912), .A2(new_n355), .A3(new_n691), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n903), .A2(KEYINPUT101), .A3(KEYINPUT39), .A4(new_n906), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n305), .A2(new_n308), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n657), .B2(new_n658), .ZN(new_n926));
  INV_X1    g0726(.A(new_n895), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n307), .A2(KEYINPUT85), .A3(new_n336), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n655), .B1(new_n324), .B2(new_n330), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n893), .A2(new_n895), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT37), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n926), .A2(new_n927), .B1(new_n932), .B2(new_n897), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n924), .B(new_n902), .C1(new_n933), .C2(KEYINPUT38), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT101), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n921), .B(new_n922), .C1(new_n923), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n659), .A2(new_n886), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n919), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n736), .A2(new_n471), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n661), .B1(new_n941), .B2(new_n732), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n939), .B(new_n942), .Z(new_n943));
  INV_X1    g0743(.A(G330), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n837), .B1(new_n910), .B2(new_n914), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n748), .A2(new_n751), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n750), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n948), .A2(new_n949), .A3(new_n906), .A4(new_n903), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n888), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n654), .A2(new_n656), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT18), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n654), .A2(KEYINPUT18), .A3(new_n656), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n651), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n897), .ZN(new_n957));
  INV_X1    g0757(.A(new_n931), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n896), .B1(new_n958), .B2(new_n952), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n956), .A2(new_n895), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n951), .B1(new_n960), .B2(new_n900), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n945), .A2(new_n947), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT40), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n950), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n471), .A2(new_n947), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n944), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n965), .B2(new_n964), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n943), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n203), .B2(new_n758), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n943), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n882), .B1(new_n969), .B2(new_n970), .ZN(G367));
  NOR2_X1   g0771(.A1(new_n822), .A2(new_n769), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n207), .B2(new_n392), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n813), .B2(new_n238), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT106), .Z(new_n975));
  AOI22_X1  g0775(.A1(new_n789), .A2(G283), .B1(G303), .B2(new_n791), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n852), .A2(G97), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n978), .B2(new_n776), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n800), .A2(new_n549), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n262), .B1(new_n509), .B2(new_n781), .C1(new_n980), .C2(KEYINPUT46), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n979), .B(new_n981), .C1(KEYINPUT46), .C2(new_n980), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G294), .A2(new_n796), .B1(new_n794), .B2(G311), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n976), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n789), .A2(G50), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G143), .A2(new_n794), .B1(new_n796), .B2(G159), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n852), .A2(G77), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n315), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT107), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n777), .A2(G137), .B1(G58), .B2(new_n771), .ZN(new_n990));
  INV_X1    g0790(.A(G150), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n990), .B1(new_n991), .B2(new_n790), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G68), .B2(new_n782), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n985), .A2(new_n986), .A3(new_n989), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n984), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n764), .B(new_n975), .C1(new_n996), .C2(new_n769), .ZN(new_n997));
  INV_X1    g0797(.A(new_n822), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n625), .A2(new_n639), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n692), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n673), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n662), .A2(new_n999), .A3(new_n692), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n997), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n706), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n564), .A2(new_n691), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(new_n703), .B2(new_n1006), .ZN(new_n1007));
  OR4_X1    g0807(.A1(KEYINPUT105), .A2(new_n826), .A3(new_n1007), .A4(new_n944), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT105), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n699), .A2(new_n1009), .A3(G330), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT105), .B1(new_n826), .B2(new_n944), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1011), .A3(new_n1007), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n737), .A2(new_n755), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n679), .A2(new_n692), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n538), .A2(new_n1015), .B1(new_n681), .B2(new_n692), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(new_n709), .A3(KEYINPUT45), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1016), .B2(new_n708), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT104), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1022), .B(KEYINPUT44), .C1(new_n1017), .C2(new_n709), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT44), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1022), .A2(KEYINPUT44), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1016), .A2(new_n708), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1021), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n705), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n705), .A2(new_n1021), .A3(new_n1023), .A4(new_n1026), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n756), .B1(new_n1014), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n711), .B(KEYINPUT41), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n762), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n705), .A2(new_n1016), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1016), .A2(new_n706), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT42), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n720), .B1(new_n1016), .B2(new_n602), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n691), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1003), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT43), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n1042), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT103), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1045), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1048), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(KEYINPUT103), .B1(new_n1054), .B2(new_n1044), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1037), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1050), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(KEYINPUT103), .A3(new_n1044), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n1036), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1004), .B1(new_n1035), .B2(new_n1060), .ZN(G387));
  INV_X1    g0861(.A(new_n713), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n815), .A2(new_n1062), .B1(new_n509), .B2(new_n208), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n388), .A2(new_n390), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n442), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT50), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n289), .B1(new_n218), .B2(new_n220), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1066), .A2(new_n1062), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n813), .B1(new_n235), .B2(new_n289), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1063), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n764), .B1(new_n1070), .B2(new_n972), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n704), .B2(new_n998), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n977), .B(new_n315), .C1(new_n220), .C2(new_n800), .ZN(new_n1073));
  XOR2_X1   g0873(.A(KEYINPUT108), .B(G150), .Z(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n777), .B2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n785), .A2(new_n218), .B1(new_n790), .B2(new_n442), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n781), .A2(new_n392), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n796), .A2(new_n387), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n794), .A2(G159), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1075), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n782), .A2(G283), .B1(new_n771), .B2(G294), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT109), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n789), .A2(G303), .B1(G317), .B2(new_n791), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n803), .A2(new_n795), .B1(new_n793), .B2(new_n804), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT110), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(KEYINPUT110), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT48), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1089), .B2(new_n1088), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT49), .Z(new_n1092));
  AOI21_X1  g0892(.A(new_n315), .B1(new_n777), .B2(G326), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n549), .B2(new_n773), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1081), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1072), .B1(new_n1095), .B2(new_n769), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n762), .B2(new_n1013), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n756), .A2(new_n1013), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1014), .A2(new_n711), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  INV_X1    g0900(.A(new_n1031), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n762), .ZN(new_n1102));
  INV_X1    g0902(.A(G97), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n813), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n972), .B1(new_n1103), .B2(new_n207), .C1(new_n1104), .C2(new_n245), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n765), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n789), .A2(new_n1064), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n796), .A2(G50), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n315), .B1(new_n800), .B2(new_n218), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n860), .B(new_n1109), .C1(G143), .C2(new_n777), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n782), .A2(G77), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n793), .A2(new_n991), .B1(new_n790), .B2(new_n847), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT51), .Z(new_n1114));
  OAI221_X1 g0914(.A(new_n262), .B1(new_n773), .B2(new_n509), .C1(new_n799), .C2(new_n800), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G322), .B2(new_n777), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n786), .A2(G294), .B1(G116), .B2(new_n782), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n543), .C2(new_n795), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n793), .A2(new_n978), .B1(new_n790), .B2(new_n803), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1112), .A2(new_n1114), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1106), .B1(new_n1122), .B2(new_n769), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1017), .B2(new_n998), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1102), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1014), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n712), .B1(new_n1126), .B2(new_n1101), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1014), .A2(new_n1031), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(G390));
  AOI21_X1  g0930(.A(new_n944), .B1(new_n946), .B2(new_n750), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n945), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(new_n935), .A3(new_n934), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1134), .A2(new_n920), .B1(new_n1136), .B2(new_n922), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n836), .A2(new_n415), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n691), .B(new_n1138), .C1(new_n734), .C2(new_n735), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n834), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n921), .B(new_n961), .C1(new_n1140), .C2(new_n915), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n922), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n915), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n832), .A2(new_n834), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT99), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n832), .A2(new_n916), .A3(new_n834), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1144), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1143), .B1(new_n1148), .B2(new_n921), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n902), .B1(new_n933), .B2(KEYINPUT38), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1140), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n920), .B(new_n1150), .C1(new_n1151), .C2(new_n1144), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n754), .A2(G330), .A3(new_n945), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1149), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1142), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n471), .A2(new_n1131), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n942), .A2(KEYINPUT112), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n661), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n691), .B1(new_n726), .B2(new_n729), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT89), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT29), .B1(new_n1161), .B2(new_n730), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1158), .B(new_n1156), .C1(new_n1162), .C2(new_n940), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT112), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n754), .A2(G330), .A3(new_n872), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1166), .A2(new_n1144), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1167), .A2(new_n1133), .B1(new_n917), .B2(new_n918), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n838), .A2(new_n1131), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1144), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1151), .A2(new_n1170), .A3(new_n1153), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1157), .A2(new_n1165), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n712), .B1(new_n1155), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1165), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1177), .A2(new_n1154), .A3(new_n1142), .A4(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1143), .A2(new_n820), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n765), .B1(new_n387), .B2(new_n843), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n793), .A2(new_n799), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n853), .A2(new_n262), .A3(new_n772), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(G294), .C2(new_n777), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n509), .B2(new_n795), .C1(new_n846), .C2(new_n1103), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1111), .B1(new_n549), .B2(new_n790), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT113), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n771), .A2(new_n1074), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT53), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G132), .B2(new_n863), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT54), .B(G143), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1190), .B1(new_n847), .B2(new_n781), .C1(new_n846), .C2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n773), .A2(new_n442), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n262), .B(new_n1193), .C1(G125), .C2(new_n777), .ZN(new_n1194));
  INV_X1    g0994(.A(G128), .ZN(new_n1195));
  INV_X1    g0995(.A(G137), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n793), .C1(new_n1196), .C2(new_n795), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n1185), .A2(new_n1187), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1181), .B1(new_n1198), .B2(new_n769), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1180), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1155), .B2(new_n759), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1179), .A2(new_n1202), .ZN(G378));
  AND2_X1   g1003(.A1(new_n937), .A2(new_n938), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n904), .A2(new_n1205), .A3(new_n907), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n949), .B1(new_n948), .B2(new_n1150), .ZN(new_n1207));
  OAI21_X1  g1007(.A(G330), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n467), .A2(new_n886), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n470), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT116), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1211), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n463), .A2(new_n466), .A3(new_n469), .A4(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1213), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1210), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT116), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1209), .A3(new_n1216), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1208), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n964), .A2(new_n1223), .A3(G330), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1204), .A2(new_n1225), .A3(new_n919), .A4(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n964), .A2(new_n1223), .A3(G330), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1223), .B1(new_n964), .B2(G330), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n939), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1230), .A3(new_n762), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n262), .A2(new_n288), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G77), .B2(new_n771), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n448), .B2(new_n773), .C1(new_n799), .C2(new_n776), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT114), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n786), .A2(new_n626), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n863), .A2(G107), .B1(new_n782), .B2(G68), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G97), .A2(new_n796), .B1(new_n794), .B2(G116), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G50), .B1(new_n445), .B2(new_n288), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1239), .A2(new_n1240), .B1(new_n1232), .B2(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(G33), .B(G41), .C1(new_n777), .C2(G124), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n794), .A2(G125), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1191), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n782), .A2(G150), .B1(new_n771), .B2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1244), .B(new_n1246), .C1(new_n1195), .C2(new_n790), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G132), .A2(new_n796), .B1(new_n786), .B2(G137), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(KEYINPUT115), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(KEYINPUT115), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1247), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT59), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1243), .B1(new_n847), .B2(new_n773), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1242), .B1(new_n1240), .B2(new_n1239), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n769), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n765), .C1(G50), .C2(new_n843), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1223), .B2(new_n820), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT117), .Z(new_n1259));
  NAND2_X1  g1059(.A1(new_n1231), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT118), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT118), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1231), .A2(new_n1262), .A3(new_n1259), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1157), .A2(new_n1165), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1153), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1137), .A2(new_n1141), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1132), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1265), .B1(new_n1269), .B2(new_n1172), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1227), .A2(new_n1230), .A3(KEYINPUT57), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n711), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1177), .B1(new_n1155), .B2(new_n1173), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT57), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1264), .B1(new_n1272), .B2(new_n1275), .ZN(G375));
  INV_X1    g1076(.A(new_n1172), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1034), .A3(new_n1173), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1144), .A2(new_n820), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT119), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n843), .A2(G68), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n315), .B1(new_n771), .B2(G97), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n987), .B(new_n1283), .C1(new_n543), .C2(new_n776), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1077), .B(new_n1284), .C1(G283), .C2(new_n863), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G116), .A2(new_n796), .B1(new_n794), .B2(G294), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1285), .B(new_n1286), .C1(new_n509), .C2(new_n846), .ZN(new_n1287));
  XOR2_X1   g1087(.A(new_n1287), .B(KEYINPUT120), .Z(new_n1288));
  AOI22_X1  g1088(.A1(G132), .A2(new_n794), .B1(new_n796), .B2(new_n1245), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n791), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(new_n1196), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(KEYINPUT121), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(KEYINPUT121), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n785), .A2(new_n991), .B1(new_n781), .B2(new_n442), .ZN(new_n1294));
  XOR2_X1   g1094(.A(new_n1294), .B(KEYINPUT122), .Z(new_n1295));
  OAI221_X1 g1095(.A(new_n315), .B1(new_n773), .B2(new_n448), .C1(new_n847), .C2(new_n800), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G128), .B2(new_n777), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1293), .A2(new_n1295), .A3(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1288), .B1(new_n1292), .B2(new_n1298), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n764), .B(new_n1282), .C1(new_n1299), .C2(new_n769), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1172), .A2(new_n762), .B1(new_n1281), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1279), .A2(new_n1301), .ZN(G381));
  OAI211_X1 g1102(.A(new_n829), .B(new_n1097), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(G381), .A2(G384), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1201), .B1(new_n1178), .B2(new_n1174), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1129), .B(new_n1004), .C1(new_n1035), .C2(new_n1060), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1308), .A2(G375), .ZN(G407));
  INV_X1    g1109(.A(G213), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(G343), .ZN(new_n1311));
  XOR2_X1   g1111(.A(new_n1311), .B(KEYINPUT123), .Z(new_n1312));
  NAND2_X1  g1112(.A1(new_n1305), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G407), .B(G213), .C1(G375), .C2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(KEYINPUT124), .ZN(G409));
  NAND2_X1  g1115(.A1(G387), .A2(G390), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1306), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G393), .A2(G396), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1303), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT61), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1316), .A2(new_n1306), .A3(new_n1319), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(G378), .B(new_n1264), .C1(new_n1272), .C2(new_n1275), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1273), .A2(new_n1034), .A3(new_n1274), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1305), .B1(new_n1326), .B2(new_n1260), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1312), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(G384), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1173), .A2(new_n711), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1278), .A2(KEYINPUT60), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT60), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1265), .A2(new_n1332), .A3(new_n1277), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1330), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1301), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1329), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1330), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1332), .B1(new_n1265), .B2(new_n1277), .ZN(new_n1338));
  AOI211_X1 g1138(.A(KEYINPUT60), .B(new_n1172), .C1(new_n1157), .C2(new_n1165), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1337), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(G384), .A3(new_n1301), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1336), .A2(new_n1341), .A3(KEYINPUT63), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1324), .B1(new_n1328), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1311), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1334), .A2(new_n1329), .A3(new_n1335), .ZN(new_n1346));
  AOI21_X1  g1146(.A(G384), .B1(new_n1340), .B2(new_n1301), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1344), .A2(new_n1345), .A3(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT63), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1312), .ZN(new_n1352));
  INV_X1    g1152(.A(G2897), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(new_n1336), .B2(new_n1341), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1345), .A2(new_n1353), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1355), .B1(new_n1348), .B2(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1311), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT125), .ZN(new_n1359));
  NOR3_X1   g1159(.A1(new_n1357), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1336), .A2(new_n1341), .A3(new_n1356), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1362), .B1(new_n1348), .B2(new_n1354), .ZN(new_n1363));
  AOI21_X1  g1163(.A(KEYINPUT125), .B1(new_n1361), .B2(new_n1363), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1343), .B(new_n1351), .C1(new_n1360), .C2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT126), .ZN(new_n1366));
  AND3_X1   g1166(.A1(new_n1316), .A2(new_n1306), .A3(new_n1319), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1319), .B1(new_n1316), .B2(new_n1306), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1366), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1321), .A2(KEYINPUT126), .A3(new_n1323), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT62), .ZN(new_n1372));
  NOR3_X1   g1172(.A1(new_n1346), .A2(new_n1347), .A3(new_n1372), .ZN(new_n1373));
  AOI22_X1  g1173(.A1(new_n1349), .A2(new_n1372), .B1(new_n1328), .B2(new_n1373), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1322), .B1(new_n1357), .B2(new_n1328), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1371), .B1(new_n1374), .B2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1365), .A2(new_n1376), .ZN(G405));
  XNOR2_X1  g1177(.A(G375), .B(G378), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1348), .A2(KEYINPUT127), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT127), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1381), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1382));
  AND3_X1   g1182(.A1(new_n1369), .A2(new_n1370), .A3(new_n1382), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1382), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1384));
  NOR3_X1   g1184(.A1(new_n1380), .A2(new_n1383), .A3(new_n1384), .ZN(new_n1385));
  INV_X1    g1185(.A(new_n1382), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1371), .A2(new_n1386), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1369), .A2(new_n1370), .A3(new_n1382), .ZN(new_n1388));
  AOI22_X1  g1188(.A1(new_n1387), .A2(new_n1388), .B1(new_n1379), .B2(new_n1378), .ZN(new_n1389));
  NOR2_X1   g1189(.A1(new_n1385), .A2(new_n1389), .ZN(G402));
endmodule


