

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n360) );
  XNOR2_X1 U324 ( .A(n361), .B(n360), .ZN(n391) );
  XNOR2_X1 U325 ( .A(n431), .B(n295), .ZN(n296) );
  XNOR2_X1 U326 ( .A(n375), .B(n296), .ZN(n297) );
  XNOR2_X1 U327 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U328 ( .A(n307), .B(n306), .ZN(n546) );
  INV_X1 U329 ( .A(G190GAT), .ZN(n447) );
  NOR2_X1 U330 ( .A1(n519), .A2(n446), .ZN(n551) );
  XNOR2_X1 U331 ( .A(n447), .B(KEYINPUT58), .ZN(n448) );
  XNOR2_X1 U332 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT64), .B(KEYINPUT74), .Z(n292) );
  XNOR2_X1 U334 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n298) );
  XOR2_X1 U336 ( .A(G29GAT), .B(G43GAT), .Z(n294) );
  XNOR2_X1 U337 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n375) );
  XOR2_X1 U339 ( .A(G50GAT), .B(G162GAT), .Z(n431) );
  AND2_X1 U340 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U341 ( .A(n298), .B(n297), .Z(n307) );
  XOR2_X1 U342 ( .A(G92GAT), .B(G85GAT), .Z(n300) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G106GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n367) );
  XNOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n301), .B(G218GAT), .ZN(n328) );
  XNOR2_X1 U347 ( .A(n367), .B(n328), .ZN(n305) );
  XOR2_X1 U348 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n303) );
  XNOR2_X1 U349 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U351 ( .A(KEYINPUT75), .B(n546), .ZN(n529) );
  XOR2_X1 U352 ( .A(KEYINPUT81), .B(G71GAT), .Z(n309) );
  XNOR2_X1 U353 ( .A(G176GAT), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n321) );
  XOR2_X1 U355 ( .A(G190GAT), .B(G99GAT), .Z(n313) );
  XOR2_X1 U356 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n311) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n336) );
  XNOR2_X1 U359 ( .A(G15GAT), .B(n336), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U361 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n315) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U364 ( .A(n317), .B(n316), .Z(n319) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U367 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U368 ( .A(G127GAT), .B(G134GAT), .Z(n323) );
  XNOR2_X1 U369 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U371 ( .A(G113GAT), .B(n324), .Z(n409) );
  XOR2_X2 U372 ( .A(n325), .B(n409), .Z(n519) );
  XOR2_X1 U373 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n445) );
  XOR2_X1 U374 ( .A(KEYINPUT71), .B(G64GAT), .Z(n327) );
  XNOR2_X1 U375 ( .A(G176GAT), .B(G204GAT), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n364) );
  XOR2_X1 U377 ( .A(n328), .B(KEYINPUT94), .Z(n330) );
  NAND2_X1 U378 ( .A1(G226GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n333) );
  XOR2_X1 U380 ( .A(G8GAT), .B(G183GAT), .Z(n349) );
  XNOR2_X1 U381 ( .A(G92GAT), .B(n349), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n331), .B(KEYINPUT93), .ZN(n332) );
  XOR2_X1 U383 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U384 ( .A(G211GAT), .B(KEYINPUT21), .Z(n335) );
  XNOR2_X1 U385 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n430) );
  XNOR2_X1 U387 ( .A(n336), .B(n430), .ZN(n337) );
  XNOR2_X1 U388 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U389 ( .A(n364), .B(n339), .ZN(n505) );
  XOR2_X1 U390 ( .A(KEYINPUT36), .B(KEYINPUT102), .Z(n340) );
  XNOR2_X1 U391 ( .A(n529), .B(n340), .ZN(n578) );
  XOR2_X1 U392 ( .A(KEYINPUT79), .B(KEYINPUT76), .Z(n342) );
  XNOR2_X1 U393 ( .A(KEYINPUT14), .B(KEYINPUT80), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U395 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n344) );
  XNOR2_X1 U396 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n359) );
  XOR2_X1 U399 ( .A(G64GAT), .B(G78GAT), .Z(n348) );
  XNOR2_X1 U400 ( .A(G127GAT), .B(G211GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n350) );
  XOR2_X1 U402 ( .A(n350), .B(n349), .Z(n357) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G1GAT), .Z(n376) );
  XOR2_X1 U404 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n352) );
  XNOR2_X1 U405 ( .A(G71GAT), .B(G57GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n366) );
  XOR2_X1 U407 ( .A(G22GAT), .B(G155GAT), .Z(n425) );
  XOR2_X1 U408 ( .A(n366), .B(n425), .Z(n354) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n376), .B(n355), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n359), .B(n358), .Z(n543) );
  INV_X1 U414 ( .A(n543), .ZN(n575) );
  NAND2_X1 U415 ( .A1(n578), .A2(n575), .ZN(n361) );
  XOR2_X1 U416 ( .A(G148GAT), .B(G78GAT), .Z(n428) );
  XOR2_X1 U417 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n363) );
  XNOR2_X1 U418 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U420 ( .A(n365), .B(n364), .Z(n369) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U423 ( .A(n428), .B(n370), .Z(n372) );
  NAND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n571) );
  XOR2_X1 U426 ( .A(G22GAT), .B(G197GAT), .Z(n374) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(G113GAT), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n389) );
  XOR2_X1 U429 ( .A(n376), .B(n375), .Z(n378) );
  XNOR2_X1 U430 ( .A(G50GAT), .B(G36GAT), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U432 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n380) );
  NAND2_X1 U433 ( .A1(G229GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U435 ( .A(n382), .B(n381), .Z(n387) );
  XOR2_X1 U436 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n384) );
  XNOR2_X1 U437 ( .A(G141GAT), .B(G8GAT), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n385), .B(KEYINPUT29), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n568) );
  NOR2_X1 U442 ( .A1(n571), .A2(n568), .ZN(n390) );
  AND2_X1 U443 ( .A1(n391), .A2(n390), .ZN(n393) );
  INV_X1 U444 ( .A(KEYINPUT109), .ZN(n392) );
  XNOR2_X1 U445 ( .A(n393), .B(n392), .ZN(n399) );
  XNOR2_X1 U446 ( .A(KEYINPUT41), .B(n571), .ZN(n536) );
  INV_X1 U447 ( .A(n536), .ZN(n550) );
  NAND2_X1 U448 ( .A1(n550), .A2(n568), .ZN(n394) );
  XNOR2_X1 U449 ( .A(KEYINPUT46), .B(n394), .ZN(n395) );
  XOR2_X1 U450 ( .A(KEYINPUT108), .B(n575), .Z(n557) );
  NAND2_X1 U451 ( .A1(n395), .A2(n557), .ZN(n396) );
  NOR2_X1 U452 ( .A1(n546), .A2(n396), .ZN(n397) );
  XOR2_X1 U453 ( .A(KEYINPUT47), .B(n397), .Z(n398) );
  NOR2_X1 U454 ( .A1(n399), .A2(n398), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n400), .B(KEYINPUT48), .ZN(n514) );
  NOR2_X1 U456 ( .A1(n505), .A2(n514), .ZN(n401) );
  XNOR2_X1 U457 ( .A(KEYINPUT54), .B(n401), .ZN(n565) );
  NAND2_X1 U458 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XOR2_X1 U459 ( .A(G155GAT), .B(G148GAT), .Z(n403) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(G1GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U462 ( .A(G162GAT), .B(G85GAT), .Z(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n421) );
  XOR2_X1 U466 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n411) );
  XNOR2_X1 U467 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n413) );
  XNOR2_X1 U470 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U473 ( .A(KEYINPUT88), .B(KEYINPUT2), .Z(n417) );
  XNOR2_X1 U474 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U476 ( .A(G141GAT), .B(n418), .Z(n438) );
  XOR2_X1 U477 ( .A(n419), .B(n438), .Z(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n564) );
  XOR2_X1 U479 ( .A(KEYINPUT23), .B(KEYINPUT85), .Z(n423) );
  XNOR2_X1 U480 ( .A(G204GAT), .B(KEYINPUT84), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U482 ( .A(n424), .B(G106GAT), .Z(n427) );
  XNOR2_X1 U483 ( .A(n425), .B(G218GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U485 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U488 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n435) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U491 ( .A(n437), .B(n436), .Z(n441) );
  INV_X1 U492 ( .A(n438), .ZN(n439) );
  XOR2_X1 U493 ( .A(n439), .B(KEYINPUT86), .Z(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n459) );
  INV_X1 U495 ( .A(n459), .ZN(n442) );
  AND2_X1 U496 ( .A1(n564), .A2(n442), .ZN(n443) );
  AND2_X1 U497 ( .A1(n565), .A2(n443), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U499 ( .A(n551), .ZN(n556) );
  NOR2_X1 U500 ( .A1(n529), .A2(n556), .ZN(n449) );
  INV_X1 U501 ( .A(n568), .ZN(n534) );
  NOR2_X1 U502 ( .A1(n534), .A2(n571), .ZN(n482) );
  XNOR2_X1 U503 ( .A(KEYINPUT27), .B(n505), .ZN(n456) );
  NOR2_X1 U504 ( .A1(n564), .A2(n456), .ZN(n512) );
  XOR2_X1 U505 ( .A(n459), .B(KEYINPUT66), .Z(n450) );
  XNOR2_X1 U506 ( .A(KEYINPUT28), .B(n450), .ZN(n517) );
  NAND2_X1 U507 ( .A1(n512), .A2(n517), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n451), .B(KEYINPUT95), .ZN(n452) );
  NAND2_X1 U509 ( .A1(n452), .A2(n519), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(KEYINPUT96), .ZN(n465) );
  XOR2_X1 U511 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n455) );
  NAND2_X1 U512 ( .A1(n459), .A2(n519), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(n567) );
  NOR2_X1 U514 ( .A1(n567), .A2(n456), .ZN(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT98), .B(n457), .Z(n462) );
  NOR2_X1 U516 ( .A1(n519), .A2(n505), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U518 ( .A(KEYINPUT25), .B(n460), .ZN(n461) );
  NAND2_X1 U519 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n564), .A2(n463), .ZN(n464) );
  NAND2_X1 U521 ( .A1(n465), .A2(n464), .ZN(n478) );
  NAND2_X1 U522 ( .A1(n575), .A2(n529), .ZN(n466) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(n466), .Z(n467) );
  AND2_X1 U524 ( .A1(n478), .A2(n467), .ZN(n493) );
  NAND2_X1 U525 ( .A1(n482), .A2(n493), .ZN(n476) );
  NOR2_X1 U526 ( .A1(n564), .A2(n476), .ZN(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n470), .ZN(G1324GAT) );
  NOR2_X1 U530 ( .A1(n505), .A2(n476), .ZN(n471) );
  XOR2_X1 U531 ( .A(G8GAT), .B(n471), .Z(G1325GAT) );
  NOR2_X1 U532 ( .A1(n476), .A2(n519), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n473) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT101), .ZN(n472) );
  XNOR2_X1 U535 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NOR2_X1 U537 ( .A1(n517), .A2(n476), .ZN(n477) );
  XOR2_X1 U538 ( .A(G22GAT), .B(n477), .Z(G1327GAT) );
  NAND2_X1 U539 ( .A1(n543), .A2(n478), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT103), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n480), .A2(n578), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(n481), .ZN(n503) );
  NAND2_X1 U543 ( .A1(n503), .A2(n482), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n491) );
  NOR2_X1 U546 ( .A1(n564), .A2(n491), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NOR2_X1 U549 ( .A1(n505), .A2(n491), .ZN(n487) );
  XOR2_X1 U550 ( .A(G36GAT), .B(n487), .Z(G1329GAT) );
  NOR2_X1 U551 ( .A1(n519), .A2(n491), .ZN(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  NOR2_X1 U555 ( .A1(n517), .A2(n491), .ZN(n492) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n492), .Z(G1331GAT) );
  NOR2_X1 U557 ( .A1(n568), .A2(n536), .ZN(n502) );
  NAND2_X1 U558 ( .A1(n502), .A2(n493), .ZN(n499) );
  NOR2_X1 U559 ( .A1(n564), .A2(n499), .ZN(n494) );
  XOR2_X1 U560 ( .A(G57GAT), .B(n494), .Z(n495) );
  XNOR2_X1 U561 ( .A(KEYINPUT42), .B(n495), .ZN(G1332GAT) );
  NOR2_X1 U562 ( .A1(n505), .A2(n499), .ZN(n496) );
  XOR2_X1 U563 ( .A(G64GAT), .B(n496), .Z(G1333GAT) );
  NOR2_X1 U564 ( .A1(n519), .A2(n499), .ZN(n497) );
  XOR2_X1 U565 ( .A(KEYINPUT106), .B(n497), .Z(n498) );
  XNOR2_X1 U566 ( .A(G71GAT), .B(n498), .ZN(G1334GAT) );
  NOR2_X1 U567 ( .A1(n517), .A2(n499), .ZN(n501) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n501), .B(n500), .ZN(G1335GAT) );
  NAND2_X1 U570 ( .A1(n503), .A2(n502), .ZN(n509) );
  NOR2_X1 U571 ( .A1(n564), .A2(n509), .ZN(n504) );
  XOR2_X1 U572 ( .A(G85GAT), .B(n504), .Z(G1336GAT) );
  NOR2_X1 U573 ( .A1(n505), .A2(n509), .ZN(n507) );
  XNOR2_X1 U574 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(G1337GAT) );
  NOR2_X1 U576 ( .A1(n519), .A2(n509), .ZN(n508) );
  XOR2_X1 U577 ( .A(G99GAT), .B(n508), .Z(G1338GAT) );
  NOR2_X1 U578 ( .A1(n517), .A2(n509), .ZN(n510) );
  XOR2_X1 U579 ( .A(KEYINPUT44), .B(n510), .Z(n511) );
  XNOR2_X1 U580 ( .A(G106GAT), .B(n511), .ZN(G1339GAT) );
  INV_X1 U581 ( .A(n512), .ZN(n513) );
  OR2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U583 ( .A(KEYINPUT110), .B(n515), .ZN(n533) );
  INV_X1 U584 ( .A(n533), .ZN(n516) );
  NAND2_X1 U585 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n523) );
  NAND2_X1 U587 ( .A1(n523), .A2(n568), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(n520), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT49), .Z(n522) );
  NAND2_X1 U590 ( .A1(n523), .A2(n550), .ZN(n521) );
  XNOR2_X1 U591 ( .A(n522), .B(n521), .ZN(G1341GAT) );
  INV_X1 U592 ( .A(n523), .ZN(n528) );
  NOR2_X1 U593 ( .A1(n557), .A2(n528), .ZN(n524) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(n524), .Z(n525) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n525), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n527) );
  XNOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n526) );
  XNOR2_X1 U598 ( .A(n527), .B(n526), .ZN(n531) );
  NOR2_X1 U599 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U600 ( .A(n531), .B(n530), .Z(n532) );
  XNOR2_X1 U601 ( .A(KEYINPUT111), .B(n532), .ZN(G1343GAT) );
  NOR2_X1 U602 ( .A1(n567), .A2(n533), .ZN(n545) );
  INV_X1 U603 ( .A(n545), .ZN(n542) );
  NOR2_X1 U604 ( .A1(n534), .A2(n542), .ZN(n535) );
  XOR2_X1 U605 ( .A(G141GAT), .B(n535), .Z(G1344GAT) );
  NOR2_X1 U606 ( .A1(n536), .A2(n542), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n538) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n537) );
  XNOR2_X1 U609 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U610 ( .A(KEYINPUT114), .B(n539), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U613 ( .A(G155GAT), .B(n544), .Z(G1346GAT) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT116), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n548), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n568), .A2(n551), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n549), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT118), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n553) );
  NAND2_X1 U621 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G183GAT), .B(n558), .Z(G1350GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT119), .B(KEYINPUT121), .Z(n560) );
  XNOR2_X1 U627 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U629 ( .A(n561), .B(KEYINPUT122), .Z(n563) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT120), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n568), .A2(n579), .ZN(n569) );
  XOR2_X1 U635 ( .A(n570), .B(n569), .Z(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n573) );
  NAND2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NAND2_X1 U640 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT124), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1355GAT) );
endmodule

