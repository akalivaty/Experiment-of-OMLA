//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND4_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT74), .A4(KEYINPUT16), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n188), .B2(KEYINPUT16), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G128), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(new_n201), .C1(G119), .C2(new_n200), .ZN(new_n202));
  XNOR2_X1  g016(.A(G119), .B(G128), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  OAI22_X1  g018(.A1(new_n202), .A2(G110), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n188), .A2(new_n190), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n196), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n211), .B(KEYINPUT75), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT22), .B(G137), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n202), .A2(G110), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n204), .A2(new_n203), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n206), .B(new_n191), .C1(new_n192), .C2(new_n194), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n196), .B2(new_n219), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n209), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n220), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n214), .B1(new_n222), .B2(new_n208), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT78), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n208), .A3(new_n214), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n215), .B1(new_n209), .B2(new_n220), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G217), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT72), .B(G902), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G234), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G902), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n233), .B(KEYINPUT73), .Z(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  INV_X1    g052(.A(new_n232), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n227), .B2(new_n226), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT77), .B(new_n238), .C1(new_n240), .C2(KEYINPUT76), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n232), .B1(new_n221), .B2(new_n223), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT25), .B1(new_n240), .B2(KEYINPUT77), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n237), .B(new_n241), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n235), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(G237), .A2(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(KEYINPUT27), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(G134), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n260), .A3(KEYINPUT66), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n258), .A3(G134), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n262), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT69), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT66), .B1(new_n256), .B2(G137), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n258), .A2(G134), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n261), .A2(new_n262), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n206), .A2(G143), .ZN(new_n277));
  INV_X1    g091(.A(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT1), .B1(new_n278), .B2(G146), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(G128), .A3(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n277), .B(new_n279), .C1(KEYINPUT1), .C2(new_n200), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n269), .A2(new_n276), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(KEYINPUT65), .A2(G131), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n261), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n257), .A2(new_n259), .A3(new_n286), .A4(new_n260), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT0), .A4(G128), .ZN(new_n293));
  XNOR2_X1  g107(.A(G143), .B(G146), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G128), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n288), .A2(KEYINPUT68), .A3(new_n289), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n292), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(G116), .B(G119), .Z(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT2), .B(G113), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n285), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n285), .A2(new_n299), .A3(KEYINPUT70), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n273), .A2(new_n275), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n284), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n297), .A2(new_n290), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n309), .B1(new_n308), .B2(new_n284), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n302), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n306), .A2(new_n307), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT28), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n304), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n312), .B2(new_n313), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n285), .A2(new_n299), .A3(KEYINPUT30), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n302), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(new_n306), .A3(new_n307), .A4(new_n253), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n306), .A2(new_n307), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n327), .A2(KEYINPUT31), .A3(new_n253), .A4(new_n323), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n254), .A2(new_n319), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G472), .A2(G902), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT32), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n319), .A2(new_n254), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(new_n328), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT32), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n330), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n306), .A2(KEYINPUT71), .A3(new_n307), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n285), .A2(new_n299), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n302), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT71), .B1(new_n306), .B2(new_n307), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT28), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND4_X1   g158(.A1(KEYINPUT29), .A2(new_n344), .A3(new_n318), .A4(new_n253), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n316), .A2(new_n318), .A3(new_n253), .ZN(new_n346));
  INV_X1    g160(.A(new_n323), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n306), .A2(new_n307), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n254), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n232), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G472), .B1(new_n345), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n248), .B1(new_n338), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G902), .ZN(new_n355));
  OR2_X1    g169(.A1(KEYINPUT83), .A2(G143), .ZN(new_n356));
  NAND2_X1  g170(.A1(KEYINPUT83), .A2(G143), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n356), .A2(new_n357), .B1(new_n249), .B2(G214), .ZN(new_n358));
  INV_X1    g172(.A(G237), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n210), .A3(G214), .ZN(new_n360));
  NOR2_X1   g174(.A1(KEYINPUT83), .A2(G143), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT18), .A2(G131), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n188), .A2(new_n190), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G146), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n363), .A2(new_n364), .B1(new_n207), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n357), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n360), .B1(new_n368), .B2(new_n361), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n356), .A2(G214), .A3(new_n249), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n364), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT84), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n374), .B(new_n364), .C1(new_n369), .C2(new_n370), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n367), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT85), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n367), .B(new_n378), .C1(new_n373), .C2(new_n375), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n262), .B1(new_n369), .B2(new_n370), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT17), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n196), .A2(new_n382), .A3(new_n219), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n371), .A2(G131), .ZN(new_n386));
  OR3_X1    g200(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n381), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n196), .A2(new_n382), .A3(KEYINPUT88), .A4(new_n219), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G113), .B(G122), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT87), .B(G104), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n390), .B(new_n391), .Z(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n380), .B2(new_n389), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n355), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G475), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT86), .B1(new_n386), .B2(new_n381), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n363), .A2(new_n262), .ZN(new_n399));
  INV_X1    g213(.A(new_n381), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT86), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  XOR2_X1   g216(.A(new_n365), .B(KEYINPUT19), .Z(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n206), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n398), .A2(new_n402), .A3(new_n404), .A4(new_n196), .ZN(new_n405));
  INV_X1    g219(.A(new_n379), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n372), .B1(new_n358), .B2(new_n362), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n374), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n371), .A2(KEYINPUT84), .A3(new_n372), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n378), .B1(new_n410), .B2(new_n367), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n405), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n392), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n393), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT89), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n417));
  NOR2_X1   g231(.A1(G475), .A2(G902), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n416), .A2(new_n417), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(new_n420), .A3(new_n417), .A4(new_n418), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n397), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G214), .B1(G237), .B2(G902), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n210), .A2(G952), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(G234), .B2(G237), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n210), .B1(G234), .B2(G237), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n239), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT93), .Z(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(G898), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G104), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT3), .B1(new_n433), .B2(G107), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT3), .ZN(new_n435));
  INV_X1    g249(.A(G107), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(G104), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(G107), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(G101), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n439), .A2(G101), .ZN(new_n442));
  INV_X1    g256(.A(G101), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n434), .A2(new_n437), .A3(new_n443), .A4(new_n438), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT4), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n302), .B(new_n441), .C1(new_n442), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT5), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n198), .A3(G116), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT79), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G116), .B(G119), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(new_n449), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n450), .A2(new_n452), .A3(G113), .A4(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n300), .A2(new_n301), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n433), .A2(G107), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n436), .A2(G104), .ZN(new_n457));
  OAI21_X1  g271(.A(G101), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n454), .A2(new_n455), .A3(new_n444), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n446), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n446), .A2(new_n461), .A3(new_n459), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n463), .A2(KEYINPUT80), .A3(new_n464), .A4(KEYINPUT6), .ZN(new_n465));
  NAND2_X1  g279(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n460), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n297), .A2(G125), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n282), .A2(new_n283), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n468), .B1(G125), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n210), .A2(G224), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n465), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(KEYINPUT82), .A2(KEYINPUT7), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n471), .A2(KEYINPUT7), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n454), .A2(new_n455), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n444), .A2(new_n458), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(KEYINPUT81), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n482), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n461), .B(KEYINPUT8), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n470), .A2(KEYINPUT7), .A3(new_n471), .A4(new_n476), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n479), .A2(new_n464), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n355), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n473), .A2(new_n475), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n488), .A2(new_n355), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n465), .A2(new_n467), .A3(new_n472), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n474), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n424), .B(new_n432), .C1(new_n490), .C2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT9), .B(G234), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n495), .A2(new_n231), .A3(G953), .ZN(new_n496));
  INV_X1    g310(.A(G116), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G122), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT91), .B1(new_n498), .B2(KEYINPUT14), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G122), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G116), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n498), .B2(KEYINPUT14), .ZN(new_n505));
  OAI21_X1  g319(.A(G107), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n498), .A3(new_n436), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n278), .A2(G128), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n200), .A2(G143), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n256), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n510), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G134), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n504), .A2(new_n498), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G107), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n200), .B2(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n510), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n509), .A2(new_n518), .ZN(new_n521));
  OAI21_X1  g335(.A(G134), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n522), .A3(new_n511), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n506), .A2(new_n514), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n517), .A2(new_n522), .A3(KEYINPUT90), .A4(new_n511), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n496), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n498), .A2(KEYINPUT14), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n505), .B1(new_n531), .B2(new_n499), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n514), .B1(new_n436), .B2(new_n532), .ZN(new_n533));
  AND4_X1   g347(.A1(new_n526), .A2(new_n528), .A3(new_n533), .A4(new_n496), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n232), .B1(new_n527), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G478), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  OAI211_X1 g353(.A(KEYINPUT92), .B(new_n232), .C1(new_n527), .C2(new_n534), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n535), .A2(new_n539), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n423), .A2(new_n494), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G221), .B1(new_n495), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G469), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n292), .A2(new_n298), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n469), .A2(new_n481), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT10), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n297), .B(new_n441), .C1(new_n442), .C2(new_n445), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n469), .B2(new_n481), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n548), .A2(new_n550), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n292), .A2(new_n298), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n469), .B(new_n481), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G140), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n210), .A2(G227), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n283), .A2(new_n282), .B1(new_n444), .B2(new_n458), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n290), .B1(new_n549), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT12), .ZN(new_n565));
  AND4_X1   g379(.A1(new_n554), .A2(new_n558), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n555), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n562), .B1(new_n568), .B2(new_n554), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n547), .B(new_n232), .C1(new_n566), .C2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n547), .A2(new_n355), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n558), .A2(new_n554), .A3(new_n565), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n561), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n554), .A3(new_n562), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(G469), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n546), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n354), .A2(new_n544), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(G101), .ZN(G3));
  OAI21_X1  g394(.A(G472), .B1(new_n329), .B2(new_n239), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n335), .A2(new_n330), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n248), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n578), .ZN(new_n585));
  OR3_X1    g399(.A1(new_n583), .A2(new_n585), .A3(KEYINPUT94), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT94), .B1(new_n583), .B2(new_n585), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT95), .Z(new_n589));
  AND2_X1   g403(.A1(new_n537), .A2(new_n540), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n525), .A2(new_n526), .A3(new_n496), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n528), .A2(new_n533), .A3(new_n526), .ZN(new_n592));
  INV_X1    g406(.A(new_n496), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n595), .B(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n239), .A2(new_n538), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n590), .A2(new_n538), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n423), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n494), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n589), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT34), .B(G104), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  AOI21_X1  g421(.A(new_n417), .B1(new_n415), .B2(new_n418), .ZN(new_n608));
  INV_X1    g422(.A(new_n418), .ZN(new_n609));
  AOI211_X1 g423(.A(KEYINPUT20), .B(new_n609), .C1(new_n414), .C2(new_n393), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n543), .B(new_n397), .C1(new_n608), .C2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n494), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n589), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT97), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NAND2_X1  g430(.A1(new_n222), .A2(new_n208), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n214), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n234), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n247), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n578), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n544), .A2(new_n582), .A3(new_n623), .A4(new_n581), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT98), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT37), .B(G110), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  AOI21_X1  g441(.A(new_n622), .B1(new_n338), .B2(new_n353), .ZN(new_n628));
  INV_X1    g442(.A(new_n611), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n630));
  INV_X1    g444(.A(new_n424), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n475), .B1(new_n473), .B2(new_n489), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n491), .A2(new_n474), .A3(new_n492), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n426), .B(KEYINPUT99), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n429), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n629), .A2(new_n630), .A3(new_n634), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n415), .A2(new_n418), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT20), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n644), .A2(new_n397), .A3(new_n543), .A4(new_n639), .ZN(new_n645));
  INV_X1    g459(.A(new_n634), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT100), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n628), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND2_X1  g463(.A1(new_n327), .A2(new_n323), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n253), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n355), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n342), .A2(new_n343), .A3(new_n253), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n338), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT101), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n638), .B(KEYINPUT39), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n578), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n490), .A2(new_n493), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT38), .Z(new_n662));
  AOI21_X1  g476(.A(new_n420), .B1(new_n414), .B2(new_n393), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n641), .B1(KEYINPUT20), .B2(new_n663), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n664), .A2(new_n421), .B1(G475), .B2(new_n396), .ZN(new_n665));
  INV_X1    g479(.A(new_n543), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n621), .A2(new_n631), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n660), .A2(new_n662), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n656), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n278), .ZN(G45));
  NAND3_X1  g485(.A1(new_n423), .A2(new_n602), .A3(new_n639), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n646), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n628), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  OAI21_X1  g489(.A(new_n232), .B1(new_n566), .B2(new_n569), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G469), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n678), .A3(new_n570), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n676), .A2(KEYINPUT102), .A3(G469), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n546), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n354), .A2(new_n604), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT103), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n682), .B(new_n684), .ZN(G15));
  NAND2_X1  g499(.A1(new_n338), .A2(new_n353), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n584), .A3(new_n612), .A4(new_n681), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  NAND4_X1  g502(.A1(new_n665), .A2(new_n432), .A3(new_n621), .A4(new_n666), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n679), .A2(new_n680), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n634), .A3(new_n545), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n686), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  XOR2_X1   g508(.A(new_n330), .B(KEYINPUT104), .Z(new_n695));
  AOI21_X1  g509(.A(new_n253), .B1(new_n344), .B2(new_n318), .ZN(new_n696));
  INV_X1    g510(.A(new_n334), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n581), .A2(new_n698), .A3(new_n584), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n494), .A2(new_n665), .A3(new_n666), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n681), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  NOR2_X1   g516(.A1(new_n672), .A2(new_n691), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n581), .A2(new_n698), .A3(new_n621), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT105), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n664), .A2(new_n421), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n601), .B1(new_n707), .B2(new_n397), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n634), .A3(new_n639), .A4(new_n681), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n581), .A2(new_n698), .A3(new_n621), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n706), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  NOR3_X1   g527(.A1(new_n490), .A2(new_n493), .A3(new_n631), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n575), .A2(KEYINPUT106), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n574), .A2(new_n716), .A3(new_n561), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(G469), .A3(new_n576), .A4(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n546), .B1(new_n573), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n672), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n354), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n354), .A2(KEYINPUT42), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  NOR2_X1   g541(.A1(new_n720), .A2(new_n645), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n354), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n575), .B2(new_n576), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n547), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n715), .A2(KEYINPUT45), .A3(new_n576), .A4(new_n717), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n735));
  OR3_X1    g549(.A1(new_n734), .A2(new_n735), .A3(new_n571), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n735), .B1(new_n734), .B2(new_n571), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n570), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n545), .A3(new_n657), .A4(new_n714), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n423), .A2(KEYINPUT43), .A3(new_n601), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n665), .B2(new_n602), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n583), .B2(new_n621), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n247), .A2(new_n620), .ZN(new_n746));
  AOI211_X1 g560(.A(KEYINPUT107), .B(new_n746), .C1(new_n581), .C2(new_n582), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n743), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n739), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(KEYINPUT44), .B(new_n743), .C1(new_n745), .C2(new_n747), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G137), .ZN(G39));
  NAND2_X1  g567(.A1(new_n738), .A2(new_n545), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n738), .A2(KEYINPUT47), .A3(new_n545), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n714), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n686), .A2(new_n584), .A3(new_n672), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G140), .ZN(G42));
  NAND2_X1  g576(.A1(new_n681), .A2(new_n714), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT115), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n764), .A2(new_n636), .A3(new_n743), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(new_n354), .ZN(new_n766));
  NOR2_X1   g580(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n767));
  AND2_X1   g581(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n656), .A2(new_n584), .A3(new_n426), .A4(new_n764), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n603), .ZN(new_n772));
  INV_X1    g586(.A(new_n691), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n743), .A2(new_n636), .A3(new_n699), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n425), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n662), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(new_n631), .A3(new_n776), .A4(new_n681), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n771), .A2(new_n423), .A3(new_n602), .ZN(new_n782));
  INV_X1    g596(.A(new_n690), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n545), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n714), .B(new_n774), .C1(new_n758), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n765), .A2(new_n704), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n770), .B(new_n775), .C1(new_n781), .C2(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n782), .A2(new_n785), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n788), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n682), .A2(new_n687), .A3(new_n693), .A4(new_n701), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT110), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n700), .A2(new_n681), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n797), .A2(new_n699), .B1(new_n692), .B2(new_n686), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n682), .A4(new_n687), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n644), .A2(new_n397), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n543), .A3(new_n638), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n628), .A2(new_n714), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n721), .A2(new_n704), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n729), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n724), .B2(new_n725), .ZN(new_n807));
  INV_X1    g621(.A(new_n494), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n423), .A2(KEYINPUT111), .A3(new_n666), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT111), .B1(new_n423), .B2(new_n666), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n603), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n586), .A2(new_n808), .A3(new_n811), .A4(new_n587), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n579), .A3(new_n624), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n801), .A2(new_n807), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n796), .B2(new_n800), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT112), .A3(new_n807), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n746), .A2(new_n719), .A3(new_n639), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n655), .A2(new_n634), .A3(new_n667), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n712), .A2(new_n821), .A3(new_n648), .A4(new_n674), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT52), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n817), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n647), .A2(new_n640), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n705), .A2(new_n711), .B1(new_n826), .B2(new_n628), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n823), .B1(new_n815), .B2(new_n816), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n834), .B2(new_n819), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT54), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n825), .A2(new_n830), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n813), .A2(new_n830), .ZN(new_n839));
  INV_X1    g653(.A(new_n795), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n807), .A3(new_n829), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n823), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n837), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n794), .A2(new_n836), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(G952), .B2(G953), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n776), .A2(new_n665), .A3(new_n602), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(KEYINPUT49), .B2(new_n783), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n783), .A2(KEYINPUT49), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT109), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n584), .A2(new_n424), .A3(new_n545), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT108), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n848), .A2(new_n656), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n846), .A2(new_n853), .ZN(G75));
  NOR2_X1   g668(.A1(new_n210), .A2(G952), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT117), .Z(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n837), .A2(new_n843), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n239), .A3(new_n475), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n465), .A2(new_n467), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(new_n472), .Z(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT55), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n860), .A3(new_n864), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n857), .B1(new_n866), .B2(new_n867), .ZN(G51));
  XNOR2_X1  g682(.A(new_n571), .B(KEYINPUT57), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n838), .B1(new_n837), .B2(new_n843), .ZN(new_n870));
  AOI211_X1 g684(.A(KEYINPUT54), .B(new_n842), .C1(new_n825), .C2(new_n830), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n566), .A2(new_n569), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n858), .A2(new_n239), .A3(new_n734), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n855), .B1(new_n874), .B2(new_n875), .ZN(G54));
  NAND2_X1  g690(.A1(KEYINPUT58), .A2(G475), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n858), .A2(new_n239), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n393), .A3(new_n414), .ZN(new_n880));
  INV_X1    g694(.A(new_n855), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n858), .A2(new_n239), .A3(new_n415), .A4(new_n878), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G60));
  NAND2_X1  g697(.A1(G478), .A2(G902), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT59), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n599), .B(new_n885), .C1(new_n870), .C2(new_n871), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n856), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n836), .A2(new_n844), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n599), .B1(new_n888), .B2(new_n885), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n889), .ZN(G63));
  XNOR2_X1  g704(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n231), .A2(new_n355), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n837), .B2(new_n843), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(new_n230), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n619), .B(KEYINPUT119), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n893), .B(new_n897), .C1(new_n835), .C2(new_n842), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(KEYINPUT61), .A3(new_n856), .A4(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n898), .B(new_n856), .C1(new_n895), .C2(new_n230), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(G66));
  INV_X1    g717(.A(new_n818), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n210), .ZN(new_n905));
  INV_X1    g719(.A(G224), .ZN(new_n906));
  OAI21_X1  g720(.A(G953), .B1(new_n430), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(KEYINPUT120), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(KEYINPUT120), .B2(new_n905), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n862), .B1(G898), .B2(new_n210), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n909), .B(new_n910), .Z(G69));
  NAND2_X1  g725(.A1(new_n321), .A2(new_n322), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT121), .Z(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n403), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n658), .A2(new_n759), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n811), .A2(new_n354), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n752), .A2(new_n761), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n670), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n712), .A2(KEYINPUT122), .A3(new_n648), .A4(new_n674), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT122), .B1(new_n827), .B2(new_n674), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n917), .B1(new_n922), .B2(KEYINPUT62), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT105), .B1(new_n703), .B2(new_n704), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n709), .A2(new_n710), .A3(new_n706), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n648), .B(new_n674), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n919), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n930));
  AND4_X1   g744(.A1(KEYINPUT123), .A2(new_n929), .A3(new_n930), .A4(new_n918), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n670), .B1(new_n928), .B2(new_n919), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT123), .B1(new_n932), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n923), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n914), .B1(new_n934), .B2(new_n210), .ZN(new_n935));
  INV_X1    g749(.A(new_n657), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n667), .A2(new_n634), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n754), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n354), .B1(new_n938), .B2(new_n728), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n761), .A3(new_n726), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n942));
  AOI221_X4 g756(.A(new_n942), .B1(new_n750), .B2(new_n751), .C1(new_n928), .C2(new_n919), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT124), .B1(new_n929), .B2(new_n752), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(KEYINPUT125), .B(new_n941), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n210), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n914), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(G900), .B2(G953), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n935), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n210), .B1(G227), .B2(G900), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n952), .A2(KEYINPUT126), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n952), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n954), .A2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n934), .B2(new_n904), .ZN(new_n961));
  INV_X1    g775(.A(new_n651), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n855), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n349), .ZN(new_n964));
  INV_X1    g778(.A(new_n324), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n834), .A2(new_n819), .A3(new_n831), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n837), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI211_X1 g784(.A(KEYINPUT127), .B(new_n966), .C1(new_n837), .C2(new_n967), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n947), .A2(new_n818), .A3(new_n948), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n253), .B(new_n650), .C1(new_n973), .C2(new_n960), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(G57));
endmodule


