//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT66), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT69), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT67), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT70), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  INV_X1    g054(.A(new_n466), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n463), .B1(new_n480), .B2(new_n464), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n480), .B2(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n463), .A2(G138), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n469), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n490), .B(KEYINPUT4), .C1(new_n465), .C2(new_n466), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n489), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n499), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n501), .A2(KEYINPUT71), .A3(new_n493), .A4(new_n494), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT72), .B1(new_n505), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT73), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(new_n505), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n510), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT74), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n510), .A2(new_n514), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n515), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(G651), .B1(G50), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n522), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  AND3_X1   g106(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT75), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT75), .B1(new_n510), .B2(new_n514), .ZN(new_n533));
  OAI211_X1 g108(.A(G63), .B(G651), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n518), .A2(G89), .A3(new_n519), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G51), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n534), .A2(new_n535), .A3(new_n539), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  INV_X1    g118(.A(G651), .ZN(new_n544));
  OAI21_X1  g119(.A(G64), .B1(new_n532), .B2(new_n533), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT77), .B(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n518), .A2(new_n519), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n537), .A2(G52), .A3(new_n538), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n547), .A2(new_n551), .ZN(G171));
  OAI21_X1  g127(.A(G56), .B1(new_n532), .B2(new_n533), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n544), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n518), .A2(G81), .A3(new_n519), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n537), .A2(G43), .A3(new_n538), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n524), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT79), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(G65), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n544), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n518), .A2(G91), .A3(new_n519), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  AOI22_X1  g154(.A1(new_n521), .A2(G87), .B1(G49), .B2(new_n528), .ZN(new_n580));
  AND2_X1   g155(.A1(G74), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n524), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT75), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n581), .B1(new_n585), .B2(G651), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(KEYINPUT80), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  AOI211_X1 g163(.A(new_n588), .B(new_n581), .C1(new_n585), .C2(G651), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n580), .B1(new_n587), .B2(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n524), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n528), .A2(G48), .ZN(new_n597));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n520), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  AND2_X1   g176(.A1(new_n585), .A2(G60), .ZN(new_n602));
  AND2_X1   g177(.A1(G72), .A2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n537), .A2(new_n538), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n521), .A2(G85), .B1(new_n605), .B2(G47), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n520), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n518), .A2(KEYINPUT10), .A3(G92), .A4(new_n519), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n605), .A2(G54), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n567), .A2(G66), .A3(new_n568), .ZN(new_n615));
  AND2_X1   g190(.A1(G79), .A2(G543), .ZN(new_n616));
  OAI21_X1  g191(.A(G651), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n608), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n608), .B1(new_n619), .B2(G868), .ZN(G321));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(G299), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(G168), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n622), .B2(G168), .ZN(G280));
  INV_X1    g200(.A(G860), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n618), .B1(G559), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT82), .Z(G148));
  OR2_X1    g203(.A1(new_n618), .A2(G559), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT83), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n476), .A2(new_n469), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n481), .A2(G123), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n483), .A2(G135), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n640), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n637), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT85), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2451), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2435), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2438), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n648), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G14), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  AOI21_X1  g240(.A(KEYINPUT18), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n673), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  AOI22_X1  g254(.A1(new_n677), .A2(KEYINPUT20), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n681), .A2(new_n673), .A3(new_n676), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n680), .B(new_n682), .C1(KEYINPUT20), .C2(new_n677), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT87), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(G229));
  NAND2_X1  g266(.A1(new_n481), .A2(G119), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  OR2_X1    g268(.A1(G95), .A2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n694), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT90), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n483), .A2(G131), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g273(.A1(KEYINPUT88), .A2(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(KEYINPUT88), .A2(G29), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n698), .S(new_n701), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G1986), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G24), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G290), .B2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n705), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(G6), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n600), .B2(new_n707), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n707), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n707), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G1971), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n715), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n707), .A2(G23), .ZN(new_n721));
  INV_X1    g296(.A(G288), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n707), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT33), .B(G1976), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT91), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n720), .B(new_n726), .C1(G1971), .C2(new_n718), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n710), .B1(new_n727), .B2(KEYINPUT34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n709), .A2(new_n706), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n728), .B(new_n729), .C1(KEYINPUT34), .C2(new_n727), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT36), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n701), .A2(G27), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G164), .B2(new_n701), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT97), .B(G2078), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n707), .A2(G4), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n619), .B2(new_n707), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT93), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT92), .B(G1348), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n739), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G5), .A2(G16), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G171), .B2(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G1961), .ZN(new_n745));
  NOR2_X1   g320(.A1(G16), .A2(G19), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n559), .B2(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G1341), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT23), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n707), .A2(G20), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n749), .B(new_n750), .C1(G299), .C2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n749), .B2(new_n750), .ZN(new_n752));
  INV_X1    g327(.A(G1956), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n742), .A2(new_n745), .A3(new_n748), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n701), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G34), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G34), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G29), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n478), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT94), .Z(new_n765));
  NOR2_X1   g340(.A1(new_n755), .A2(new_n765), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(new_n463), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G139), .B2(new_n483), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n475), .A2(G103), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT25), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G29), .ZN(new_n775));
  OR2_X1    g350(.A1(G29), .A2(G33), .ZN(new_n776));
  AOI21_X1  g351(.A(G2072), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G29), .A2(G32), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n476), .A2(G105), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT26), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n483), .A2(G141), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n481), .A2(G129), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n779), .A2(new_n781), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT27), .B(G1996), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n775), .A2(G2072), .A3(new_n776), .ZN(new_n789));
  INV_X1    g364(.A(G28), .ZN(new_n790));
  AOI21_X1  g365(.A(G29), .B1(new_n790), .B2(KEYINPUT30), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n790), .A2(KEYINPUT30), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n789), .B(new_n794), .C1(new_n642), .C2(new_n756), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n777), .A2(new_n788), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT31), .B(G11), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n756), .A2(KEYINPUT28), .A3(G26), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n481), .A2(G128), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n483), .A2(G140), .ZN(new_n800));
  OR2_X1    g375(.A1(G104), .A2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n801), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(new_n761), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT28), .B1(new_n756), .B2(G26), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2067), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n756), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n756), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT29), .B(G2090), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n796), .A2(new_n797), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n762), .A2(new_n763), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n744), .B2(G1961), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n786), .B2(new_n787), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT96), .ZN(new_n817));
  NAND2_X1  g392(.A1(G168), .A2(G16), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G16), .B2(G21), .ZN(new_n819));
  INV_X1    g394(.A(G1966), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n821), .B(new_n822), .C1(new_n747), .C2(G1341), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n813), .A2(new_n817), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n766), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n731), .A2(new_n736), .A3(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  NAND2_X1  g402(.A1(new_n619), .A2(G559), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n518), .A2(G93), .A3(new_n519), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n537), .A2(G55), .A3(new_n538), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n583), .B2(new_n584), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(G651), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n831), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(G67), .B1(new_n532), .B2(new_n533), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n544), .B1(new_n841), .B2(new_n837), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n832), .A2(new_n833), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT98), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n840), .A2(new_n844), .B1(new_n555), .B2(new_n558), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n559), .B1(new_n842), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n830), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n626), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT99), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n840), .A2(new_n844), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G860), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT100), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT100), .B1(new_n493), .B2(new_n494), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n501), .B(new_n803), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n495), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n856), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n803), .B1(new_n863), .B2(new_n501), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n784), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n501), .B1(new_n857), .B2(new_n858), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n804), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n785), .A3(new_n859), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n774), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(KEYINPUT101), .A3(new_n774), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n865), .A2(new_n773), .A3(new_n868), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT102), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n865), .A2(new_n868), .A3(new_n876), .A4(new_n773), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n872), .A2(new_n873), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n698), .B(new_n635), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n481), .A2(G130), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n483), .A2(G142), .ZN(new_n881));
  NOR2_X1   g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n880), .B(new_n881), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n879), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT103), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n886), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n478), .B(new_n487), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n642), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n874), .A2(KEYINPUT102), .ZN(new_n892));
  INV_X1    g467(.A(new_n877), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT101), .B1(new_n869), .B2(new_n774), .ZN(new_n894));
  AOI211_X1 g469(.A(new_n871), .B(new_n773), .C1(new_n865), .C2(new_n868), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n892), .A2(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n885), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n887), .A2(new_n888), .A3(new_n891), .A4(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n896), .A2(new_n885), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n872), .A2(new_n873), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n875), .A2(new_n877), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n886), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n890), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n900), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n899), .A2(KEYINPUT104), .A3(new_n905), .A4(new_n900), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n855), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT105), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT40), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(G395));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n573), .B2(new_n577), .ZN(new_n921));
  NOR4_X1   g496(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT106), .A4(new_n576), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n921), .A2(new_n618), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n618), .A2(G299), .A3(KEYINPUT106), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G299), .A2(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(new_n922), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n619), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n618), .A2(G299), .A3(KEYINPUT106), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(KEYINPUT41), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n834), .A2(new_n839), .A3(new_n831), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT98), .B1(new_n842), .B2(new_n843), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n559), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI211_X1 g509(.A(new_n558), .B(new_n555), .C1(new_n839), .C2(new_n834), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(new_n629), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n937), .B1(new_n924), .B2(new_n923), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(G290), .A2(G166), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n604), .A2(G303), .A3(new_n606), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n942), .A2(G288), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(G288), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g520(.A(G305), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n943), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n722), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n942), .A2(G288), .A3(new_n943), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n600), .A3(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n946), .A2(new_n950), .A3(KEYINPUT107), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n941), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(new_n940), .ZN(new_n957));
  OAI21_X1  g532(.A(G868), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n851), .A2(new_n622), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(G295));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n961), .A3(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n940), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n941), .A2(new_n953), .A3(new_n954), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n622), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n959), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n962), .A2(new_n967), .ZN(G331));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n946), .A2(new_n950), .ZN(new_n970));
  INV_X1    g545(.A(G64), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n583), .B2(new_n584), .ZN(new_n972));
  INV_X1    g547(.A(new_n546), .ZN(new_n973));
  OAI21_X1  g548(.A(G651), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n974), .A2(KEYINPUT110), .A3(new_n550), .A4(new_n549), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n547), .B2(new_n551), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n977), .A3(G168), .ZN(new_n978));
  OAI211_X1 g553(.A(G286), .B(new_n976), .C1(new_n547), .C2(new_n551), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n847), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n923), .A2(new_n924), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n979), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n846), .A3(new_n845), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(KEYINPUT111), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n936), .A2(new_n987), .A3(new_n983), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n847), .A2(new_n980), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT112), .B1(new_n936), .B2(new_n983), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n986), .A2(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n925), .A2(new_n930), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n970), .B(new_n985), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n900), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n989), .B1(new_n847), .B2(new_n980), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n936), .A2(new_n983), .A3(KEYINPUT112), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n936), .A2(new_n987), .A3(new_n983), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n987), .B1(new_n936), .B2(new_n983), .ZN(new_n999));
  OAI22_X1  g574(.A1(new_n996), .A2(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n931), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n970), .B1(new_n1001), .B2(new_n985), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n969), .B1(new_n995), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n986), .A2(new_n988), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n990), .A2(new_n991), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n982), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n981), .A2(new_n984), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n931), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n970), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n969), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1012), .A2(new_n900), .A3(new_n994), .A4(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1003), .A2(new_n1004), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n970), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT43), .B1(new_n995), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n993), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1018));
  INV_X1    g593(.A(new_n985), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1011), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1020), .A2(new_n900), .A3(new_n994), .A4(new_n1013), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1004), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1015), .A2(new_n1022), .A3(KEYINPUT113), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1019), .B1(new_n1000), .B2(new_n931), .ZN(new_n1026));
  AOI21_X1  g601(.A(G37), .B1(new_n1026), .B2(new_n970), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n1027), .B2(new_n1012), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1021), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT44), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1003), .A2(new_n1004), .A3(new_n1014), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1024), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1023), .A2(new_n1032), .ZN(G397));
  XOR2_X1   g608(.A(KEYINPUT114), .B(G1384), .Z(new_n1034));
  NAND2_X1  g609(.A1(new_n866), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G40), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n478), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(G1996), .A3(new_n784), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1044));
  INV_X1    g619(.A(G2067), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n803), .A2(G2067), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G1996), .B2(new_n784), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n1043), .B(new_n1044), .C1(new_n1041), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1041), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n698), .B(new_n704), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n604), .A2(new_n706), .A3(new_n606), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G290), .A2(G1986), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n499), .B1(new_n862), .B2(new_n856), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G1384), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1060), .B2(new_n1039), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n599), .ZN(new_n1063));
  INV_X1    g638(.A(G1981), .ZN(new_n1064));
  INV_X1    g639(.A(new_n594), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n595), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n594), .A2(KEYINPUT81), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1063), .B(new_n1064), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G1981), .B1(new_n599), .B2(new_n1065), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1068), .A2(KEYINPUT49), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT49), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1062), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1976), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n722), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1068), .B(KEYINPUT118), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1062), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1384), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n500), .A2(new_n502), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT50), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n866), .A2(new_n1081), .A3(new_n1078), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1082), .A3(new_n1039), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2090), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1079), .A2(new_n1036), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n866), .A2(KEYINPUT45), .A3(new_n1034), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1039), .ZN(new_n1088));
  INV_X1    g663(.A(G1971), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1084), .A2(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G303), .A2(G8), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1090), .A2(new_n1058), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n1096));
  NAND2_X1  g671(.A1(G288), .A2(new_n1074), .ZN(new_n1097));
  OAI211_X1 g672(.A(G1976), .B(new_n580), .C1(new_n587), .C2(new_n589), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1061), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1061), .B2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1095), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n866), .A2(new_n1078), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT50), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n503), .A2(new_n1081), .A3(new_n1078), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1103), .A2(new_n1039), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1105), .A2(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1093), .B1(new_n1106), .B2(new_n1058), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1097), .A2(new_n1096), .A3(new_n1061), .A4(new_n1098), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT117), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1101), .A2(new_n1107), .A3(new_n1109), .A4(new_n1073), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1094), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1093), .B1(new_n1090), .B2(new_n1058), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1101), .A2(new_n1109), .A3(new_n1073), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT120), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1061), .A2(new_n1098), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1108), .B1(new_n1096), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1072), .B1(new_n1117), .B2(new_n1095), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1109), .A4(new_n1113), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n503), .A2(new_n1121), .A3(KEYINPUT45), .A4(new_n1078), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1102), .A2(new_n1036), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT119), .B1(new_n1079), .B2(new_n1036), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .A4(new_n1039), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1125), .A2(new_n820), .B1(new_n1084), .B2(new_n763), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1126), .A2(new_n1058), .A3(G286), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1115), .A2(new_n1120), .A3(new_n1127), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1077), .B(new_n1112), .C1(new_n1128), .C2(KEYINPUT63), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1127), .A2(new_n1111), .ZN(new_n1130));
  NAND2_X1  g705(.A1(G286), .A2(G8), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1125), .A2(new_n820), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1084), .A2(new_n763), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(KEYINPUT51), .B(G8), .C1(new_n1135), .C2(G286), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1137), .B(new_n1131), .C1(new_n1126), .C2(new_n1058), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1132), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT62), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1084), .A2(G1961), .ZN(new_n1141));
  INV_X1    g716(.A(G2078), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1086), .A2(new_n1087), .A3(new_n1142), .A4(new_n1039), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT124), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(new_n1147), .A3(new_n1144), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1040), .B1(new_n1036), .B2(new_n1102), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1144), .A2(G2078), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1124), .A3(new_n1122), .A4(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1141), .A2(new_n1146), .A3(new_n1148), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1130), .B1(new_n1140), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1129), .B1(new_n1155), .B2(new_n1110), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G299), .B(KEYINPUT57), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1103), .A2(new_n1104), .A3(new_n1039), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n753), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1087), .A2(new_n1039), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT56), .B(G2072), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n1086), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1163), .A2(KEYINPUT121), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1157), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT57), .ZN(new_n1168));
  XNOR2_X1  g743(.A(G299), .B(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1169), .A2(new_n1162), .A3(new_n1159), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1167), .A2(KEYINPUT61), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1163), .A2(new_n1157), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1170), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1060), .A2(new_n1045), .A3(new_n1039), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n1084), .B2(new_n740), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n618), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1173), .A2(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(KEYINPUT58), .B(G1341), .Z(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n1040), .B2(new_n1102), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n1088), .B2(G1996), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1182), .B(KEYINPUT122), .C1(new_n1088), .C2(G1996), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1185), .A2(new_n559), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT59), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1185), .A2(new_n1189), .A3(new_n559), .A4(new_n1186), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1178), .A2(new_n619), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1171), .A2(new_n1180), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1170), .A2(new_n619), .A3(new_n1176), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1167), .A2(new_n1194), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1193), .A2(KEYINPUT123), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT123), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1160), .A2(KEYINPUT53), .A3(new_n1142), .A4(new_n1037), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1141), .A2(new_n1146), .A3(new_n1148), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(G171), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1152), .A2(G171), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1199), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1202), .A2(new_n1203), .A3(KEYINPUT54), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1139), .A2(new_n1110), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT54), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1199), .A2(G171), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1207), .B1(new_n1154), .B2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1205), .A2(new_n1206), .A3(new_n1209), .A4(new_n1094), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1196), .A2(new_n1197), .A3(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1057), .B1(new_n1156), .B2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT48), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1053), .A2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n698), .A2(new_n703), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1050), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1051), .B1(new_n1217), .B2(new_n1046), .ZN(new_n1218));
  XNOR2_X1  g793(.A(KEYINPUT126), .B(KEYINPUT46), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1219), .B1(new_n1051), .B2(G1996), .ZN(new_n1220));
  INV_X1    g795(.A(G1996), .ZN(new_n1221));
  OAI211_X1 g796(.A(new_n1041), .B(new_n1221), .C1(KEYINPUT126), .C2(KEYINPUT46), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1048), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1041), .B1(new_n784), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1220), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  XOR2_X1   g800(.A(new_n1225), .B(KEYINPUT47), .Z(new_n1226));
  NOR3_X1   g801(.A1(new_n1215), .A2(new_n1218), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1212), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g803(.A(G401), .B1(new_n908), .B2(new_n910), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n1014), .ZN(new_n1231));
  NOR3_X1   g805(.A1(G229), .A2(new_n461), .A3(G227), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(G225));
  INV_X1    g807(.A(G225), .ZN(G308));
endmodule


