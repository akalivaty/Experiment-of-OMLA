

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770;

  NOR2_X1 U373 ( .A1(n562), .A2(n552), .ZN(n739) );
  XNOR2_X2 U374 ( .A(n411), .B(n354), .ZN(n629) );
  INV_X2 U375 ( .A(G953), .ZN(n761) );
  AND2_X1 U376 ( .A1(n404), .A2(n406), .ZN(n402) );
  NAND2_X1 U377 ( .A1(n731), .A2(n745), .ZN(n612) );
  INV_X1 U378 ( .A(n609), .ZN(n692) );
  INV_X1 U379 ( .A(n614), .ZN(n695) );
  NAND2_X1 U380 ( .A1(n361), .A2(n358), .ZN(n458) );
  AND2_X2 U381 ( .A1(n401), .A2(n400), .ZN(n678) );
  NAND2_X1 U382 ( .A1(n402), .A2(n403), .ZN(n401) );
  NAND2_X1 U383 ( .A1(n382), .A2(n630), .ZN(n689) );
  NAND2_X1 U384 ( .A1(n576), .A2(n458), .ZN(n604) );
  AND2_X1 U385 ( .A1(n480), .A2(n417), .ZN(n416) );
  AND2_X2 U386 ( .A1(n527), .A2(n589), .ZN(n576) );
  AND2_X1 U387 ( .A1(n363), .A2(n362), .ZN(n361) );
  INV_X1 U388 ( .A(n573), .ZN(n351) );
  OR2_X1 U389 ( .A1(n653), .A2(G902), .ZN(n453) );
  NAND2_X1 U390 ( .A1(n425), .A2(n424), .ZN(n516) );
  XNOR2_X1 U391 ( .A(G110), .B(KEYINPUT67), .ZN(n487) );
  XNOR2_X1 U392 ( .A(G119), .B(G110), .ZN(n436) );
  XNOR2_X1 U393 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n434) );
  XNOR2_X2 U394 ( .A(n388), .B(KEYINPUT81), .ZN(n627) );
  NAND2_X1 U395 ( .A1(n419), .A2(n495), .ZN(n410) );
  XNOR2_X1 U396 ( .A(G146), .B(G125), .ZN(n488) );
  INV_X1 U397 ( .A(KEYINPUT73), .ZN(n394) );
  XNOR2_X1 U398 ( .A(n533), .B(KEYINPUT1), .ZN(n609) );
  INV_X1 U399 ( .A(n604), .ZN(n376) );
  NAND2_X1 U400 ( .A1(n433), .A2(n360), .ZN(n359) );
  XNOR2_X1 U401 ( .A(n380), .B(n379), .ZN(n378) );
  XNOR2_X1 U402 ( .A(G143), .B(G131), .ZN(n380) );
  XNOR2_X1 U403 ( .A(KEYINPUT94), .B(KEYINPUT12), .ZN(n379) );
  XNOR2_X1 U404 ( .A(n507), .B(n508), .ZN(n381) );
  XNOR2_X1 U405 ( .A(G140), .B(G113), .ZN(n507) );
  XNOR2_X1 U406 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n508) );
  INV_X1 U407 ( .A(KEYINPUT10), .ZN(n439) );
  INV_X1 U408 ( .A(G122), .ZN(n482) );
  INV_X1 U409 ( .A(KEYINPUT11), .ZN(n505) );
  XOR2_X1 U410 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n504) );
  INV_X1 U411 ( .A(KEYINPUT64), .ZN(n409) );
  INV_X1 U412 ( .A(G214), .ZN(n475) );
  NAND2_X1 U413 ( .A1(n372), .A2(n368), .ZN(n399) );
  NAND2_X1 U414 ( .A1(n604), .A2(n369), .ZN(n368) );
  NAND2_X1 U415 ( .A1(n376), .A2(n373), .ZN(n372) );
  NAND2_X1 U416 ( .A1(n371), .A2(n370), .ZN(n369) );
  INV_X1 U417 ( .A(n458), .ZN(n533) );
  XNOR2_X1 U418 ( .A(n493), .B(n492), .ZN(n494) );
  AND2_X1 U419 ( .A1(n753), .A2(n355), .ZN(n383) );
  INV_X1 U420 ( .A(n396), .ZN(n393) );
  XNOR2_X1 U421 ( .A(n415), .B(n414), .ZN(n721) );
  XNOR2_X1 U422 ( .A(KEYINPUT101), .B(KEYINPUT33), .ZN(n414) );
  AND2_X1 U423 ( .A1(n578), .A2(n692), .ZN(n415) );
  NAND2_X1 U424 ( .A1(n351), .A2(n478), .ZN(n385) );
  INV_X1 U425 ( .A(n689), .ZN(n400) );
  NOR2_X1 U426 ( .A1(G953), .A2(G237), .ZN(n502) );
  INV_X1 U427 ( .A(n528), .ZN(n465) );
  NAND2_X1 U428 ( .A1(n352), .A2(n459), .ZN(n371) );
  NAND2_X1 U429 ( .A1(KEYINPUT104), .A2(KEYINPUT75), .ZN(n370) );
  NAND2_X1 U430 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U431 ( .A1(n459), .A2(KEYINPUT75), .ZN(n374) );
  NAND2_X1 U432 ( .A1(n352), .A2(KEYINPUT104), .ZN(n375) );
  XNOR2_X1 U433 ( .A(G128), .B(KEYINPUT23), .ZN(n435) );
  INV_X1 U434 ( .A(G128), .ZN(n423) );
  INV_X1 U435 ( .A(KEYINPUT8), .ZN(n441) );
  XNOR2_X1 U436 ( .A(G140), .B(G137), .ZN(n443) );
  XNOR2_X1 U437 ( .A(G131), .B(G134), .ZN(n426) );
  NOR2_X1 U438 ( .A1(G902), .A2(G237), .ZN(n474) );
  OR2_X1 U439 ( .A1(n465), .A2(KEYINPUT75), .ZN(n417) );
  NAND2_X1 U440 ( .A1(G469), .A2(G902), .ZN(n362) );
  XNOR2_X1 U441 ( .A(G116), .B(G107), .ZN(n517) );
  XNOR2_X1 U442 ( .A(G134), .B(G122), .ZN(n514) );
  XNOR2_X1 U443 ( .A(n513), .B(n512), .ZN(n631) );
  XNOR2_X1 U444 ( .A(n510), .B(n509), .ZN(n513) );
  XNOR2_X1 U445 ( .A(n381), .B(n378), .ZN(n509) );
  AND2_X1 U446 ( .A1(n409), .A2(n420), .ZN(n405) );
  XOR2_X1 U447 ( .A(G104), .B(G107), .Z(n428) );
  XNOR2_X1 U448 ( .A(G146), .B(G101), .ZN(n427) );
  OR2_X1 U449 ( .A1(n384), .A2(n692), .ZN(n570) );
  OR2_X1 U450 ( .A1(n548), .A2(n706), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n390), .B(n501), .ZN(n575) );
  INV_X1 U452 ( .A(KEYINPUT6), .ZN(n377) );
  XNOR2_X1 U453 ( .A(n398), .B(n556), .ZN(n582) );
  NAND2_X1 U454 ( .A1(n351), .A2(n478), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n562) );
  XNOR2_X1 U456 ( .A(G475), .B(KEYINPUT13), .ZN(n386) );
  OR2_X1 U457 ( .A1(n631), .A2(G902), .ZN(n387) );
  BUF_X1 U458 ( .A(n544), .Z(n698) );
  BUF_X1 U459 ( .A(n527), .Z(n614) );
  INV_X1 U460 ( .A(n646), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n631), .B(KEYINPUT59), .ZN(n632) );
  XNOR2_X1 U462 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U463 ( .A1(n634), .A2(G953), .ZN(n683) );
  NAND2_X1 U464 ( .A1(n383), .A2(n393), .ZN(n382) );
  XNOR2_X1 U465 ( .A(n418), .B(KEYINPUT40), .ZN(n541) );
  NAND2_X1 U466 ( .A1(n575), .A2(n739), .ZN(n418) );
  OR2_X1 U467 ( .A1(n548), .A2(n385), .ZN(n550) );
  INV_X1 U468 ( .A(n653), .ZN(n654) );
  NAND2_X1 U469 ( .A1(n465), .A2(KEYINPUT75), .ZN(n352) );
  AND2_X1 U470 ( .A1(n621), .A2(n620), .ZN(n353) );
  INV_X1 U471 ( .A(G902), .ZN(n360) );
  XOR2_X1 U472 ( .A(KEYINPUT80), .B(KEYINPUT45), .Z(n354) );
  XNOR2_X1 U473 ( .A(n470), .B(n443), .ZN(n643) );
  AND2_X1 U474 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n355) );
  INV_X1 U475 ( .A(KEYINPUT2), .ZN(n420) );
  XNOR2_X2 U476 ( .A(n357), .B(n356), .ZN(n483) );
  XNOR2_X2 U477 ( .A(G119), .B(KEYINPUT3), .ZN(n356) );
  XNOR2_X2 U478 ( .A(G113), .B(G101), .ZN(n357) );
  XNOR2_X1 U479 ( .A(n453), .B(n452), .ZN(n527) );
  OR2_X1 U480 ( .A1(n671), .A2(n359), .ZN(n358) );
  NAND2_X1 U481 ( .A1(n671), .A2(G469), .ZN(n363) );
  XNOR2_X1 U482 ( .A(n470), .B(n364), .ZN(n661) );
  XNOR2_X1 U483 ( .A(n365), .B(n468), .ZN(n364) );
  XNOR2_X1 U484 ( .A(n483), .B(n366), .ZN(n365) );
  XNOR2_X1 U485 ( .A(n469), .B(n367), .ZN(n366) );
  INV_X1 U486 ( .A(G116), .ZN(n367) );
  XNOR2_X2 U487 ( .A(n392), .B(n426), .ZN(n470) );
  XNOR2_X2 U488 ( .A(n516), .B(KEYINPUT4), .ZN(n392) );
  XNOR2_X1 U489 ( .A(n544), .B(n377), .ZN(n597) );
  XNOR2_X2 U490 ( .A(n473), .B(n472), .ZN(n544) );
  XNOR2_X1 U491 ( .A(n643), .B(n432), .ZN(n671) );
  NAND2_X2 U492 ( .A1(n627), .A2(n642), .ZN(n396) );
  NAND2_X1 U493 ( .A1(n389), .A2(n641), .ZN(n388) );
  XNOR2_X1 U494 ( .A(n569), .B(n568), .ZN(n389) );
  NAND2_X1 U495 ( .A1(n564), .A2(n500), .ZN(n390) );
  XNOR2_X1 U496 ( .A(n391), .B(n481), .ZN(n564) );
  NAND2_X1 U497 ( .A1(n399), .A2(n416), .ZN(n391) );
  XNOR2_X1 U498 ( .A(n392), .B(n486), .ZN(n493) );
  NAND2_X1 U499 ( .A1(n753), .A2(n393), .ZN(n687) );
  XNOR2_X2 U500 ( .A(n396), .B(n394), .ZN(n622) );
  XNOR2_X1 U501 ( .A(n396), .B(n395), .ZN(n645) );
  XNOR2_X2 U502 ( .A(n397), .B(n583), .ZN(n607) );
  NAND2_X1 U503 ( .A1(n582), .A2(n581), .ZN(n397) );
  NAND2_X1 U504 ( .A1(n408), .A2(n407), .ZN(n403) );
  NAND2_X1 U505 ( .A1(n622), .A2(n405), .ZN(n404) );
  NAND2_X1 U506 ( .A1(n410), .A2(n409), .ZN(n406) );
  NAND2_X1 U507 ( .A1(n622), .A2(n420), .ZN(n407) );
  NOR2_X1 U508 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X1 U509 ( .A1(n412), .A2(n353), .ZN(n411) );
  XNOR2_X1 U510 ( .A(n413), .B(n603), .ZN(n412) );
  AND2_X1 U511 ( .A1(n602), .A2(n770), .ZN(n413) );
  NAND2_X1 U512 ( .A1(n607), .A2(n721), .ZN(n585) );
  INV_X1 U513 ( .A(n541), .ZN(n658) );
  NAND2_X1 U514 ( .A1(n629), .A2(n420), .ZN(n419) );
  NOR2_X1 U515 ( .A1(n707), .A2(n706), .ZN(n421) );
  INV_X1 U516 ( .A(KEYINPUT104), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n506), .B(n505), .ZN(n510) );
  XNOR2_X1 U518 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U519 ( .A(KEYINPUT34), .ZN(n584) );
  XNOR2_X1 U520 ( .A(n585), .B(n584), .ZN(n587) );
  INV_X1 U521 ( .A(KEYINPUT74), .ZN(n481) );
  INV_X1 U522 ( .A(KEYINPUT60), .ZN(n636) );
  INV_X1 U523 ( .A(G143), .ZN(n422) );
  NAND2_X1 U524 ( .A1(G128), .A2(n422), .ZN(n425) );
  NAND2_X1 U525 ( .A1(n423), .A2(G143), .ZN(n424) );
  XNOR2_X1 U526 ( .A(n428), .B(n427), .ZN(n431) );
  NAND2_X1 U527 ( .A1(n761), .A2(G227), .ZN(n429) );
  XNOR2_X1 U528 ( .A(n487), .B(n429), .ZN(n430) );
  XNOR2_X1 U529 ( .A(n431), .B(n430), .ZN(n432) );
  INV_X1 U530 ( .A(G469), .ZN(n433) );
  XNOR2_X1 U531 ( .A(n435), .B(n434), .ZN(n438) );
  XNOR2_X1 U532 ( .A(n436), .B(KEYINPUT87), .ZN(n437) );
  XNOR2_X1 U533 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U534 ( .A(n488), .B(n439), .ZN(n644) );
  XNOR2_X1 U535 ( .A(n440), .B(n644), .ZN(n446) );
  NAND2_X1 U536 ( .A1(n761), .A2(G234), .ZN(n442) );
  XNOR2_X1 U537 ( .A(n442), .B(n441), .ZN(n520) );
  NAND2_X1 U538 ( .A1(n520), .A2(G221), .ZN(n444) );
  XNOR2_X1 U539 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U540 ( .A(n446), .B(n445), .ZN(n653) );
  INV_X1 U541 ( .A(KEYINPUT15), .ZN(n447) );
  XNOR2_X1 U542 ( .A(n447), .B(G902), .ZN(n495) );
  INV_X1 U543 ( .A(n495), .ZN(n623) );
  NAND2_X1 U544 ( .A1(n623), .A2(G234), .ZN(n449) );
  INV_X1 U545 ( .A(KEYINPUT20), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n449), .B(n448), .ZN(n455) );
  INV_X1 U547 ( .A(n455), .ZN(n450) );
  AND2_X1 U548 ( .A1(n450), .A2(G217), .ZN(n451) );
  XNOR2_X1 U549 ( .A(n451), .B(KEYINPUT25), .ZN(n452) );
  INV_X1 U550 ( .A(G221), .ZN(n454) );
  OR2_X1 U551 ( .A1(n455), .A2(n454), .ZN(n457) );
  INV_X1 U552 ( .A(KEYINPUT21), .ZN(n456) );
  XNOR2_X1 U553 ( .A(n457), .B(n456), .ZN(n589) );
  NAND2_X1 U554 ( .A1(G237), .A2(G234), .ZN(n460) );
  XNOR2_X1 U555 ( .A(n460), .B(KEYINPUT14), .ZN(n691) );
  NAND2_X1 U556 ( .A1(n761), .A2(G952), .ZN(n462) );
  NAND2_X1 U557 ( .A1(G953), .A2(G902), .ZN(n461) );
  NAND2_X1 U558 ( .A1(n462), .A2(n461), .ZN(n463) );
  AND2_X1 U559 ( .A1(n691), .A2(n463), .ZN(n580) );
  NAND2_X1 U560 ( .A1(G953), .A2(G900), .ZN(n464) );
  NAND2_X1 U561 ( .A1(n580), .A2(n464), .ZN(n528) );
  NAND2_X1 U562 ( .A1(n502), .A2(G210), .ZN(n467) );
  XOR2_X1 U563 ( .A(G137), .B(KEYINPUT72), .Z(n466) );
  XNOR2_X1 U564 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U565 ( .A(G146), .B(KEYINPUT5), .ZN(n469) );
  NAND2_X1 U566 ( .A1(n661), .A2(n360), .ZN(n473) );
  INV_X1 U567 ( .A(KEYINPUT69), .ZN(n471) );
  XNOR2_X1 U568 ( .A(n471), .B(G472), .ZN(n472) );
  XNOR2_X1 U569 ( .A(n474), .B(KEYINPUT71), .ZN(n496) );
  INV_X1 U570 ( .A(n496), .ZN(n476) );
  OR2_X1 U571 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U572 ( .A(n477), .B(KEYINPUT85), .ZN(n706) );
  INV_X1 U573 ( .A(n706), .ZN(n478) );
  AND2_X1 U574 ( .A1(n544), .A2(n478), .ZN(n479) );
  XNOR2_X1 U575 ( .A(n479), .B(KEYINPUT30), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n482), .B(G104), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n483), .B(n511), .ZN(n485) );
  XNOR2_X1 U578 ( .A(n517), .B(KEYINPUT16), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n485), .B(n484), .ZN(n760) );
  XNOR2_X1 U580 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n486) );
  XNOR2_X1 U581 ( .A(n488), .B(n487), .ZN(n491) );
  NAND2_X1 U582 ( .A1(n761), .A2(G224), .ZN(n489) );
  XNOR2_X1 U583 ( .A(n489), .B(KEYINPUT77), .ZN(n490) );
  XNOR2_X1 U584 ( .A(n760), .B(n494), .ZN(n680) );
  OR2_X1 U585 ( .A1(n680), .A2(n495), .ZN(n498) );
  NAND2_X1 U586 ( .A1(n496), .A2(G210), .ZN(n497) );
  XNOR2_X2 U587 ( .A(n498), .B(n497), .ZN(n573) );
  INV_X1 U588 ( .A(KEYINPUT38), .ZN(n499) );
  XNOR2_X1 U589 ( .A(n573), .B(n499), .ZN(n707) );
  INV_X1 U590 ( .A(n707), .ZN(n500) );
  XNOR2_X1 U591 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n501) );
  NAND2_X1 U592 ( .A1(n502), .A2(G214), .ZN(n503) );
  XNOR2_X1 U593 ( .A(n504), .B(n503), .ZN(n506) );
  XOR2_X1 U594 ( .A(n511), .B(n644), .Z(n512) );
  XOR2_X1 U595 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n515) );
  XNOR2_X1 U596 ( .A(n515), .B(n514), .ZN(n519) );
  XNOR2_X1 U597 ( .A(n516), .B(n517), .ZN(n518) );
  XNOR2_X1 U598 ( .A(n519), .B(n518), .ZN(n524) );
  AND2_X1 U599 ( .A1(n520), .A2(G217), .ZN(n522) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n521) );
  XNOR2_X1 U601 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U602 ( .A(n524), .B(n523), .ZN(n669) );
  NAND2_X1 U603 ( .A1(n669), .A2(n360), .ZN(n526) );
  INV_X1 U604 ( .A(G478), .ZN(n525) );
  XNOR2_X1 U605 ( .A(n526), .B(n525), .ZN(n561) );
  INV_X1 U606 ( .A(n561), .ZN(n552) );
  INV_X1 U607 ( .A(n589), .ZN(n694) );
  NOR2_X1 U608 ( .A1(n694), .A2(n528), .ZN(n529) );
  NAND2_X1 U609 ( .A1(n695), .A2(n529), .ZN(n530) );
  XNOR2_X1 U610 ( .A(n530), .B(KEYINPUT66), .ZN(n546) );
  INV_X1 U611 ( .A(n698), .ZN(n595) );
  NOR2_X1 U612 ( .A1(n546), .A2(n595), .ZN(n532) );
  XNOR2_X1 U613 ( .A(KEYINPUT28), .B(KEYINPUT105), .ZN(n531) );
  XNOR2_X1 U614 ( .A(n532), .B(n531), .ZN(n534) );
  NOR2_X1 U615 ( .A1(n534), .A2(n533), .ZN(n557) );
  AND2_X1 U616 ( .A1(n562), .A2(n561), .ZN(n708) );
  NAND2_X1 U617 ( .A1(n421), .A2(n708), .ZN(n535) );
  XNOR2_X1 U618 ( .A(n535), .B(KEYINPUT41), .ZN(n720) );
  NAND2_X1 U619 ( .A1(n557), .A2(n720), .ZN(n539) );
  XOR2_X1 U620 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n537) );
  INV_X1 U621 ( .A(KEYINPUT106), .ZN(n536) );
  XNOR2_X1 U622 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U623 ( .A(n539), .B(n538), .ZN(n767) );
  INV_X1 U624 ( .A(n767), .ZN(n540) );
  NAND2_X1 U625 ( .A1(n541), .A2(n540), .ZN(n543) );
  INV_X1 U626 ( .A(KEYINPUT46), .ZN(n542) );
  XNOR2_X1 U627 ( .A(n543), .B(n542), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n739), .A2(n597), .ZN(n545) );
  NOR2_X1 U629 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U630 ( .A(KEYINPUT102), .B(n547), .Z(n548) );
  XOR2_X1 U631 ( .A(KEYINPUT36), .B(KEYINPUT108), .Z(n549) );
  XNOR2_X1 U632 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U633 ( .A1(n551), .A2(n692), .ZN(n750) );
  NAND2_X1 U634 ( .A1(n562), .A2(n552), .ZN(n554) );
  INV_X1 U635 ( .A(KEYINPUT97), .ZN(n553) );
  XNOR2_X1 U636 ( .A(n554), .B(n553), .ZN(n746) );
  INV_X1 U637 ( .A(n739), .ZN(n742) );
  NAND2_X1 U638 ( .A1(n746), .A2(n742), .ZN(n555) );
  XNOR2_X1 U639 ( .A(n555), .B(KEYINPUT98), .ZN(n710) );
  XNOR2_X1 U640 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n556) );
  AND2_X1 U641 ( .A1(n557), .A2(n582), .ZN(n740) );
  NAND2_X1 U642 ( .A1(n710), .A2(n740), .ZN(n559) );
  INV_X1 U643 ( .A(KEYINPUT47), .ZN(n558) );
  XNOR2_X1 U644 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U645 ( .A1(n750), .A2(n560), .ZN(n565) );
  NOR2_X1 U646 ( .A1(n562), .A2(n561), .ZN(n586) );
  AND2_X1 U647 ( .A1(n586), .A2(n351), .ZN(n563) );
  AND2_X1 U648 ( .A1(n564), .A2(n563), .ZN(n638) );
  NOR2_X1 U649 ( .A1(n565), .A2(n638), .ZN(n566) );
  NAND2_X1 U650 ( .A1(n567), .A2(n566), .ZN(n569) );
  XNOR2_X1 U651 ( .A(KEYINPUT65), .B(KEYINPUT48), .ZN(n568) );
  XNOR2_X1 U652 ( .A(n570), .B(KEYINPUT103), .ZN(n572) );
  INV_X1 U653 ( .A(KEYINPUT43), .ZN(n571) );
  XNOR2_X1 U654 ( .A(n572), .B(n571), .ZN(n574) );
  NAND2_X1 U655 ( .A1(n574), .A2(n573), .ZN(n641) );
  INV_X1 U656 ( .A(n746), .ZN(n736) );
  NAND2_X1 U657 ( .A1(n575), .A2(n736), .ZN(n642) );
  INV_X1 U658 ( .A(n597), .ZN(n615) );
  INV_X1 U659 ( .A(n576), .ZN(n577) );
  NOR2_X1 U660 ( .A1(n615), .A2(n577), .ZN(n578) );
  XNOR2_X1 U661 ( .A(KEYINPUT86), .B(G898), .ZN(n762) );
  NAND2_X1 U662 ( .A1(n762), .A2(G953), .ZN(n579) );
  AND2_X1 U663 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U664 ( .A(KEYINPUT0), .ZN(n583) );
  NAND2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U666 ( .A(n588), .B(KEYINPUT35), .ZN(n768) );
  NAND2_X1 U667 ( .A1(n708), .A2(n589), .ZN(n591) );
  INV_X1 U668 ( .A(KEYINPUT100), .ZN(n590) );
  XNOR2_X1 U669 ( .A(n591), .B(n590), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n607), .A2(n592), .ZN(n594) );
  XNOR2_X1 U671 ( .A(KEYINPUT70), .B(KEYINPUT22), .ZN(n593) );
  XNOR2_X1 U672 ( .A(n594), .B(n593), .ZN(n600) );
  OR2_X1 U673 ( .A1(n600), .A2(n692), .ZN(n617) );
  NAND2_X1 U674 ( .A1(n595), .A2(n695), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n617), .A2(n596), .ZN(n639) );
  NOR2_X1 U676 ( .A1(n768), .A2(n639), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n597), .A2(n614), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n598), .A2(n692), .ZN(n599) );
  NOR2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U680 ( .A(KEYINPUT32), .B(n601), .Z(n770) );
  INV_X1 U681 ( .A(KEYINPUT44), .ZN(n618) );
  NAND2_X1 U682 ( .A1(n618), .A2(KEYINPUT68), .ZN(n603) );
  NOR2_X1 U683 ( .A1(n604), .A2(n698), .ZN(n605) );
  AND2_X1 U684 ( .A1(n607), .A2(n605), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n606), .B(KEYINPUT89), .ZN(n731) );
  INV_X1 U686 ( .A(n607), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n698), .A2(n576), .ZN(n608) );
  OR2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n702) );
  NOR2_X1 U689 ( .A1(n610), .A2(n702), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n611), .B(KEYINPUT31), .ZN(n745) );
  NAND2_X1 U691 ( .A1(n612), .A2(n710), .ZN(n613) );
  XOR2_X1 U692 ( .A(KEYINPUT99), .B(n613), .Z(n621) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n640) );
  NOR2_X1 U695 ( .A1(n618), .A2(KEYINPUT68), .ZN(n619) );
  NOR2_X1 U696 ( .A1(n640), .A2(n619), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n642), .A2(KEYINPUT2), .ZN(n625) );
  INV_X1 U698 ( .A(KEYINPUT78), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n629), .A2(n626), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n630) );
  INV_X1 U702 ( .A(n629), .ZN(n753) );
  NAND2_X1 U703 ( .A1(n678), .A2(G475), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n633), .B(n632), .ZN(n635) );
  INV_X1 U705 ( .A(G952), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n635), .A2(n683), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(G60) );
  XOR2_X1 U708 ( .A(G143), .B(n638), .Z(G45) );
  XOR2_X1 U709 ( .A(G110), .B(n639), .Z(G12) );
  XOR2_X1 U710 ( .A(G101), .B(n640), .Z(G3) );
  XNOR2_X1 U711 ( .A(n641), .B(G140), .ZN(G42) );
  XNOR2_X1 U712 ( .A(n642), .B(G134), .ZN(G36) );
  XNOR2_X1 U713 ( .A(n643), .B(n644), .ZN(n646) );
  NAND2_X1 U714 ( .A1(n645), .A2(n761), .ZN(n652) );
  XOR2_X1 U715 ( .A(G227), .B(n646), .Z(n647) );
  XNOR2_X1 U716 ( .A(n647), .B(KEYINPUT124), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n648), .A2(G900), .ZN(n649) );
  NAND2_X1 U718 ( .A1(G953), .A2(n649), .ZN(n650) );
  XOR2_X1 U719 ( .A(KEYINPUT125), .B(n650), .Z(n651) );
  NAND2_X1 U720 ( .A1(n652), .A2(n651), .ZN(G72) );
  NAND2_X1 U721 ( .A1(n678), .A2(G217), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U723 ( .A1(n656), .A2(n683), .ZN(n657) );
  XNOR2_X1 U724 ( .A(n657), .B(KEYINPUT121), .ZN(G66) );
  XNOR2_X1 U725 ( .A(G131), .B(KEYINPUT127), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n658), .B(n659), .ZN(G33) );
  NAND2_X1 U727 ( .A1(n678), .A2(G472), .ZN(n663) );
  XOR2_X1 U728 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n664), .A2(n683), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT84), .B(KEYINPUT63), .Z(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT83), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(G57) );
  NAND2_X1 U735 ( .A1(n678), .A2(G478), .ZN(n668) );
  XOR2_X1 U736 ( .A(n669), .B(n668), .Z(n670) );
  INV_X1 U737 ( .A(n683), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n670), .A2(n676), .ZN(G63) );
  NAND2_X1 U739 ( .A1(n678), .A2(G469), .ZN(n675) );
  XOR2_X1 U740 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n672) );
  XNOR2_X1 U741 ( .A(n672), .B(KEYINPUT58), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n671), .B(n673), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n675), .B(n674), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(G54) );
  NAND2_X1 U745 ( .A1(n678), .A2(G210), .ZN(n682) );
  XNOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n682), .B(n681), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n686) );
  XNOR2_X1 U749 ( .A(KEYINPUT119), .B(KEYINPUT56), .ZN(n685) );
  XNOR2_X1 U750 ( .A(n686), .B(n685), .ZN(G51) );
  NAND2_X1 U751 ( .A1(n687), .A2(n420), .ZN(n688) );
  XNOR2_X1 U752 ( .A(n688), .B(KEYINPUT79), .ZN(n690) );
  OR2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n727) );
  NAND2_X1 U754 ( .A1(G952), .A2(n691), .ZN(n719) );
  NOR2_X1 U755 ( .A1(n692), .A2(n576), .ZN(n693) );
  XOR2_X1 U756 ( .A(KEYINPUT50), .B(n693), .Z(n700) );
  NAND2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U758 ( .A(n696), .B(KEYINPUT49), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U761 ( .A(n701), .B(KEYINPUT116), .ZN(n703) );
  NAND2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U763 ( .A(KEYINPUT51), .B(n704), .Z(n705) );
  NAND2_X1 U764 ( .A1(n720), .A2(n705), .ZN(n715) );
  NAND2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U767 ( .A1(n421), .A2(n710), .ZN(n711) );
  NAND2_X1 U768 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U769 ( .A1(n721), .A2(n713), .ZN(n714) );
  NAND2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U771 ( .A(KEYINPUT117), .B(n716), .ZN(n717) );
  XNOR2_X1 U772 ( .A(KEYINPUT52), .B(n717), .ZN(n718) );
  NOR2_X1 U773 ( .A1(n719), .A2(n718), .ZN(n723) );
  AND2_X1 U774 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U775 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U776 ( .A(KEYINPUT118), .B(n724), .Z(n725) );
  NOR2_X1 U777 ( .A1(n725), .A2(G953), .ZN(n726) );
  NAND2_X1 U778 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U779 ( .A(KEYINPUT53), .B(n728), .Z(G75) );
  NOR2_X1 U780 ( .A1(n742), .A2(n731), .ZN(n729) );
  XOR2_X1 U781 ( .A(KEYINPUT110), .B(n729), .Z(n730) );
  XNOR2_X1 U782 ( .A(G104), .B(n730), .ZN(G6) );
  NOR2_X1 U783 ( .A1(n731), .A2(n746), .ZN(n735) );
  XOR2_X1 U784 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n733) );
  XNOR2_X1 U785 ( .A(G107), .B(KEYINPUT111), .ZN(n732) );
  XNOR2_X1 U786 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n735), .B(n734), .ZN(G9) );
  XOR2_X1 U788 ( .A(G128), .B(KEYINPUT29), .Z(n738) );
  NAND2_X1 U789 ( .A1(n740), .A2(n736), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n738), .B(n737), .ZN(G30) );
  NAND2_X1 U791 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n741), .B(G146), .ZN(G48) );
  NOR2_X1 U793 ( .A1(n742), .A2(n745), .ZN(n743) );
  XOR2_X1 U794 ( .A(KEYINPUT112), .B(n743), .Z(n744) );
  XNOR2_X1 U795 ( .A(G113), .B(n744), .ZN(G15) );
  NOR2_X1 U796 ( .A1(n746), .A2(n745), .ZN(n748) );
  XNOR2_X1 U797 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U799 ( .A(G116), .B(n749), .ZN(G18) );
  XNOR2_X1 U800 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n751) );
  XNOR2_X1 U801 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U802 ( .A(G125), .B(n752), .ZN(G27) );
  NAND2_X1 U803 ( .A1(n753), .A2(n761), .ZN(n758) );
  NAND2_X1 U804 ( .A1(G224), .A2(G953), .ZN(n754) );
  XNOR2_X1 U805 ( .A(n754), .B(KEYINPUT61), .ZN(n755) );
  XNOR2_X1 U806 ( .A(n755), .B(KEYINPUT122), .ZN(n756) );
  NAND2_X1 U807 ( .A1(n756), .A2(n762), .ZN(n757) );
  NAND2_X1 U808 ( .A1(n758), .A2(n757), .ZN(n766) );
  XNOR2_X1 U809 ( .A(G110), .B(KEYINPUT123), .ZN(n759) );
  XNOR2_X1 U810 ( .A(n760), .B(n759), .ZN(n764) );
  NOR2_X1 U811 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U812 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U813 ( .A(n766), .B(n765), .ZN(G69) );
  XOR2_X1 U814 ( .A(n767), .B(G137), .Z(G39) );
  XOR2_X1 U815 ( .A(n768), .B(G122), .Z(n769) );
  XNOR2_X1 U816 ( .A(KEYINPUT126), .B(n769), .ZN(G24) );
  XNOR2_X1 U817 ( .A(G119), .B(n770), .ZN(G21) );
endmodule

