//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1178, new_n1179, new_n1181, new_n1182, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n213), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G97), .A2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n223), .B1(new_n202), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  AND2_X1   g0028(.A1(KEYINPUT67), .A2(G77), .ZN(new_n229));
  NOR2_X1   g0029(.A1(KEYINPUT67), .A2(G77), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT68), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n210), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OR2_X1    g0035(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n237));
  AND3_X1   g0037(.A1(new_n222), .A2(new_n236), .A3(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n256), .A2(new_n208), .A3(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n214), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n207), .A2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G50), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n257), .ZN(new_n263));
  XOR2_X1   g0063(.A(KEYINPUT8), .B(G58), .Z(new_n264));
  NAND2_X1  g0064(.A1(new_n208), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n264), .A2(new_n266), .B1(G150), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(G20), .B1(new_n218), .B2(G50), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n259), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n262), .B1(G50), .B2(new_n263), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  XOR2_X1   g0072(.A(new_n272), .B(KEYINPUT9), .Z(new_n273));
  AOI21_X1  g0073(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n277), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n224), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n231), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n289), .A2(G223), .B1(new_n290), .B2(new_n287), .ZN(new_n291));
  INV_X1    g0091(.A(G222), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT3), .B(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n288), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n282), .B1(new_n295), .B2(new_n274), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(G190), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n273), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n300), .B(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n272), .B1(new_n296), .B2(G169), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G68), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n203), .B2(new_n265), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n311), .A2(new_n259), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n312), .A2(KEYINPUT11), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n257), .A2(new_n309), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT12), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(KEYINPUT11), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n260), .A2(G68), .A3(new_n261), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n313), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n274), .A2(new_n278), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(G238), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT71), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT71), .B1(G33), .B2(G97), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n294), .B2(new_n224), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n289), .A2(G232), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n322), .B1(new_n332), .B2(new_n280), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n322), .C1(new_n332), .C2(new_n280), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n319), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT14), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n336), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n304), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n337), .A2(new_n338), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n318), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n334), .A2(G190), .A3(new_n336), .ZN(new_n345));
  INV_X1    g0145(.A(new_n318), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n298), .B1(new_n334), .B2(new_n336), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n348), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n350), .A2(KEYINPUT72), .A3(new_n345), .A4(new_n346), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n260), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n264), .A2(new_n261), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n354), .A2(new_n355), .B1(new_n263), .B2(new_n264), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT7), .B1(new_n287), .B2(new_n208), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT7), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n359), .B(G20), .C1(new_n284), .C2(new_n286), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(G58), .A2(G68), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n362), .B2(new_n201), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n267), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n271), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n285), .A2(G33), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT73), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n208), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n360), .B1(new_n375), .B2(new_n359), .ZN(new_n376));
  OAI211_X1 g0176(.A(KEYINPUT16), .B(new_n366), .C1(new_n376), .C2(new_n309), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT74), .B1(new_n369), .B2(new_n377), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n357), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n279), .B1(new_n240), .B2(new_n281), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n279), .B(KEYINPUT75), .C1(new_n240), .C2(new_n281), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n293), .A2(G223), .A3(new_n288), .ZN(new_n386));
  INV_X1    g0186(.A(G87), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n293), .A2(G1698), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n386), .B1(new_n283), .B2(new_n387), .C1(new_n388), .C2(new_n224), .ZN(new_n389));
  AOI21_X1  g0189(.A(G179), .B1(new_n389), .B2(new_n274), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n381), .B1(new_n274), .B2(new_n389), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n385), .A2(new_n390), .B1(new_n392), .B2(new_n319), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n380), .A2(KEYINPUT18), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT76), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n380), .A2(new_n396), .A3(KEYINPUT18), .A4(new_n393), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT74), .ZN(new_n399));
  INV_X1    g0199(.A(new_n377), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n359), .B1(new_n293), .B2(G20), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n365), .B1(new_n403), .B2(G68), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n259), .B1(new_n404), .B2(KEYINPUT16), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n399), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n377), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n356), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n385), .A2(new_n390), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(G169), .B2(new_n391), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n398), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n395), .A2(new_n397), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n383), .A2(new_n384), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n389), .A2(new_n274), .ZN(new_n414));
  INV_X1    g0214(.A(G190), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n413), .A2(new_n416), .B1(new_n391), .B2(G200), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n357), .B(new_n417), .C1(new_n378), .C2(new_n379), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n412), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n279), .B1(new_n228), .B2(new_n281), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n289), .A2(G238), .B1(G107), .B2(new_n287), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n240), .B2(new_n294), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(new_n274), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n304), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(G20), .A2(new_n290), .B1(new_n430), .B2(new_n266), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n264), .A2(new_n267), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n271), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n260), .A2(G77), .A3(new_n261), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n290), .B2(new_n263), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n428), .B1(G169), .B2(new_n427), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n427), .A2(G190), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n433), .A2(new_n435), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(new_n438), .C1(new_n298), .C2(new_n427), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n308), .A2(new_n353), .A3(new_n423), .A4(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n293), .A2(G257), .A3(new_n288), .ZN(new_n442));
  INV_X1    g0242(.A(G303), .ZN(new_n443));
  INV_X1    g0243(.A(G264), .ZN(new_n444));
  OAI221_X1 g0244(.A(new_n442), .B1(new_n443), .B2(new_n293), .C1(new_n388), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n274), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT5), .B(G41), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(new_n274), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(G270), .B1(new_n276), .B2(new_n450), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n263), .A2(G116), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n260), .B1(G1), .B2(new_n283), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n208), .C1(G33), .C2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n259), .C1(new_n208), .C2(G116), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n461), .A2(new_n462), .ZN(new_n464));
  OAI221_X1 g0264(.A(new_n455), .B1(new_n456), .B2(new_n457), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n453), .A2(G179), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n446), .A2(new_n452), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n467), .A2(new_n465), .A3(KEYINPUT21), .A4(G169), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n465), .A3(G169), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT21), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n465), .B1(new_n467), .B2(G200), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n415), .B2(new_n467), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT19), .B1(new_n325), .B2(new_n326), .ZN(new_n477));
  NOR2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n477), .A2(new_n208), .B1(new_n387), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n293), .A2(new_n208), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n265), .A2(new_n459), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n480), .A2(new_n309), .B1(KEYINPUT19), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n259), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n429), .A2(new_n257), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n483), .A2(KEYINPUT77), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT77), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n485), .A2(new_n486), .B1(new_n429), .B2(new_n456), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G116), .ZN(new_n488));
  INV_X1    g0288(.A(G238), .ZN(new_n489));
  OAI221_X1 g0289(.A(new_n488), .B1(new_n388), .B2(new_n228), .C1(new_n489), .C2(new_n294), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n274), .ZN(new_n491));
  INV_X1    g0291(.A(G250), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n274), .A2(new_n492), .A3(new_n449), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n276), .B2(new_n449), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n304), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n487), .B(new_n497), .C1(G169), .C2(new_n496), .ZN(new_n498));
  INV_X1    g0298(.A(new_n456), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G87), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n485), .B2(new_n486), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n298), .B1(new_n491), .B2(new_n494), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n496), .B2(G190), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n480), .B2(new_n387), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n293), .A2(new_n208), .A3(G87), .A4(new_n506), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n208), .B2(G107), .ZN(new_n512));
  INV_X1    g0312(.A(G107), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(KEYINPUT23), .A3(G20), .ZN(new_n514));
  INV_X1    g0314(.A(new_n488), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n512), .A2(new_n514), .B1(new_n515), .B2(new_n208), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(KEYINPUT24), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT24), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n510), .B2(new_n516), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n259), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT25), .B1(new_n257), .B2(new_n513), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n513), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n456), .A2(new_n513), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n293), .A2(G257), .A3(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G294), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n294), .C2(new_n492), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n274), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n450), .A2(new_n276), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n447), .A2(new_n449), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n280), .A3(G264), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G169), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n533), .A2(new_n280), .A3(KEYINPUT79), .A4(G264), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n538), .A2(new_n539), .B1(new_n530), .B2(new_n274), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n532), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n536), .B1(new_n541), .B2(new_n304), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n527), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n498), .A2(new_n505), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n293), .A2(G250), .A3(G1698), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n293), .A2(G244), .A3(new_n288), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n458), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n274), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n451), .A2(G257), .B1(new_n276), .B2(new_n450), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n267), .A2(G77), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT6), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n459), .A2(new_n513), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n478), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n513), .A2(KEYINPUT6), .A3(G97), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n555), .B1(new_n561), .B2(new_n208), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n513), .B1(new_n401), .B2(new_n402), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n259), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n263), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n499), .B2(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n552), .A2(G200), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n554), .A2(new_n564), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n553), .A2(new_n304), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n552), .A2(new_n319), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n535), .A2(G190), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n541), .B2(new_n298), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n527), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n476), .A2(new_n544), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n441), .A2(new_n578), .ZN(G372));
  NAND2_X1  g0379(.A1(new_n411), .A2(new_n394), .ZN(new_n580));
  INV_X1    g0380(.A(new_n343), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n436), .B(KEYINPUT82), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n352), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n422), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n306), .B1(new_n585), .B2(new_n302), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n501), .A2(KEYINPUT81), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT81), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n500), .C1(new_n485), .C2(new_n486), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n504), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n543), .A2(new_n472), .A3(new_n469), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n577), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT80), .B1(new_n496), .B2(G169), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT80), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n495), .A2(new_n595), .A3(new_n319), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n594), .A2(new_n487), .A3(new_n497), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n572), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n498), .A2(new_n505), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT26), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n591), .A2(new_n597), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n602), .A2(KEYINPUT26), .A3(new_n572), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n441), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n586), .A2(new_n605), .ZN(G369));
  INV_X1    g0406(.A(new_n473), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT83), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT27), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(G213), .ZN(new_n613));
  INV_X1    g0413(.A(G343), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n615), .A2(new_n465), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n476), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n616), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  XOR2_X1   g0420(.A(KEYINPUT84), .B(G330), .Z(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT85), .ZN(new_n623));
  INV_X1    g0423(.A(new_n615), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n521), .B2(new_n526), .ZN(new_n625));
  OAI221_X1 g0425(.A(new_n543), .B1(new_n527), .B2(new_n575), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n625), .A2(new_n623), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n543), .B2(new_n624), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n473), .A2(new_n615), .ZN(new_n631));
  INV_X1    g0431(.A(new_n543), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(new_n624), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(G399));
  INV_X1    g0434(.A(new_n211), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(G41), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n478), .A2(new_n387), .A3(new_n457), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n636), .A2(new_n637), .A3(new_n207), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n220), .B2(new_n636), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT86), .ZN(new_n640));
  XOR2_X1   g0440(.A(new_n640), .B(KEYINPUT28), .Z(new_n641));
  NAND2_X1  g0441(.A1(new_n578), .A2(new_n624), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n496), .A2(new_n453), .A3(G179), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n541), .A3(new_n552), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n467), .A2(new_n304), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(new_n496), .A3(new_n540), .A4(new_n553), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT30), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n615), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT31), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n621), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n604), .A2(new_n624), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(KEYINPUT29), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(new_n602), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n598), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n498), .A2(new_n505), .A3(new_n598), .A4(new_n657), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n593), .A2(new_n597), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n624), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(KEYINPUT29), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n654), .A2(new_n656), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n641), .B1(new_n664), .B2(G1), .ZN(G364));
  NOR2_X1   g0465(.A1(new_n256), .A2(G20), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n207), .B1(new_n666), .B2(G45), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n636), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n622), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n621), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n619), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n214), .B1(G20), .B2(new_n319), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n208), .A2(new_n304), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(G190), .A3(new_n298), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(G190), .A2(G200), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n677), .A2(G58), .B1(new_n680), .B2(new_n290), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(KEYINPUT89), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(G200), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n415), .ZN(new_n685));
  AOI211_X1 g0485(.A(new_n287), .B(new_n683), .C1(G50), .C2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n684), .A2(G190), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n208), .A2(G179), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(G190), .A3(G200), .ZN(new_n690));
  OAI22_X1  g0490(.A1(new_n688), .A2(new_n309), .B1(new_n387), .B2(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n415), .A2(G179), .A3(G200), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n208), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n691), .B1(G97), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT32), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n689), .A2(new_n678), .ZN(new_n697));
  INV_X1    g0497(.A(G159), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n697), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT32), .A3(G159), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n682), .A2(KEYINPUT89), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n689), .A2(new_n415), .A3(G200), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT90), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G107), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n686), .A2(new_n695), .A3(new_n702), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(G283), .ZN(new_n711));
  INV_X1    g0511(.A(G322), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n676), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G311), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n287), .B1(new_n679), .B2(new_n714), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n713), .B(new_n715), .C1(G329), .C2(new_n700), .ZN(new_n716));
  XNOR2_X1  g0516(.A(KEYINPUT91), .B(G326), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(G294), .A2(new_n694), .B1(new_n685), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g0519(.A(KEYINPUT33), .B(G317), .ZN(new_n720));
  INV_X1    g0520(.A(new_n690), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n687), .A2(new_n720), .B1(new_n721), .B2(G303), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n711), .A2(new_n716), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n674), .B1(new_n710), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n673), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT73), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT73), .B1(new_n284), .B2(new_n286), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n211), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT88), .Z(new_n734));
  NAND2_X1  g0534(.A1(new_n254), .A2(G45), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n734), .B(new_n735), .C1(G45), .C2(new_n219), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n635), .A2(new_n287), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n737), .A2(G355), .B1(new_n457), .B2(new_n635), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n729), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n669), .B(KEYINPUT87), .Z(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n724), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n727), .B(KEYINPUT92), .Z(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n619), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n672), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(G396));
  NOR2_X1   g0546(.A1(new_n624), .A2(new_n438), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n582), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n440), .A2(new_n747), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT94), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n655), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n624), .B(new_n750), .C1(new_n601), .C2(new_n603), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n654), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n669), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n654), .A2(new_n752), .A3(new_n753), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n674), .A2(new_n726), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n740), .B1(G77), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G294), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n676), .A2(new_n760), .B1(new_n697), .B2(new_n714), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n293), .B(new_n761), .C1(G116), .C2(new_n680), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n708), .A2(G87), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n694), .A2(G97), .B1(new_n721), .B2(G107), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT93), .B(G283), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G303), .A2(new_n685), .B1(new_n687), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n677), .A2(G143), .B1(new_n680), .B2(G159), .ZN(new_n769));
  INV_X1    g0569(.A(new_n685), .ZN(new_n770));
  INV_X1    g0570(.A(G137), .ZN(new_n771));
  INV_X1    g0571(.A(G150), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n769), .B1(new_n770), .B2(new_n771), .C1(new_n772), .C2(new_n688), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT34), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n708), .A2(G68), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n732), .B1(G132), .B2(new_n700), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n694), .A2(G58), .B1(new_n721), .B2(G50), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n773), .A2(new_n774), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n768), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n759), .B1(new_n781), .B2(new_n673), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n750), .B2(new_n726), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n757), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G384));
  OR2_X1    g0585(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n786), .A2(G116), .A3(new_n217), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT36), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n219), .A2(new_n362), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n790), .A2(new_n231), .B1(G50), .B2(new_n309), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G1), .A3(new_n256), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT95), .Z(new_n794));
  NOR2_X1   g0594(.A1(new_n346), .A2(new_n624), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n353), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n343), .B(new_n352), .C1(new_n346), .C2(new_n624), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n436), .A2(new_n615), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n753), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT98), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n366), .B1(new_n376), .B2(new_n309), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n271), .B1(new_n804), .B2(new_n368), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT96), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n377), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(KEYINPUT96), .B(new_n271), .C1(new_n804), .C2(new_n368), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n357), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n613), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n809), .A2(new_n393), .B1(new_n408), .B2(new_n417), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT97), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(KEYINPUT7), .B1(new_n732), .B2(new_n208), .ZN(new_n815));
  OAI21_X1  g0615(.A(G68), .B1(new_n815), .B2(new_n360), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT16), .B1(new_n816), .B2(new_n366), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT96), .B1(new_n817), .B2(new_n271), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n805), .A2(new_n806), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n377), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n410), .B1(new_n820), .B2(new_n357), .ZN(new_n821));
  INV_X1    g0621(.A(new_n419), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n821), .A2(KEYINPUT97), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(KEYINPUT37), .B1(new_n814), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n380), .A2(new_n393), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n380), .A2(new_n810), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n419), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n811), .B1(new_n412), .B2(new_n422), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT38), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n828), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT97), .B1(new_n821), .B2(new_n822), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n809), .A2(new_n393), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(new_n813), .A3(new_n419), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(new_n836), .A3(new_n811), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n833), .B1(new_n837), .B2(KEYINPUT37), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n838), .A2(new_n839), .A3(new_n830), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n803), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n838), .B2(new_n830), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n829), .A2(KEYINPUT38), .A3(new_n831), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT98), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n802), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n580), .A2(new_n810), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT99), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n802), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT98), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT98), .B1(new_n842), .B2(new_n843), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT99), .ZN(new_n852));
  INV_X1    g0652(.A(new_n846), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n408), .A2(new_n398), .A3(new_n410), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT18), .B1(new_n380), .B2(new_n393), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n421), .B(new_n418), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n408), .A2(new_n613), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n419), .B1(new_n408), .B2(new_n410), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n859), .B2(new_n858), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n857), .A2(new_n858), .B1(new_n860), .B2(new_n828), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT100), .B1(new_n861), .B2(KEYINPUT38), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n860), .A2(new_n828), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n826), .B1(new_n422), .B2(new_n580), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n863), .B(new_n839), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n843), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n581), .A2(new_n624), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n847), .A2(new_n854), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n441), .B1(new_n656), .B2(new_n663), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n876), .A2(new_n586), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n875), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n642), .A2(new_n652), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n798), .A2(new_n879), .A3(new_n750), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n849), .B2(new_n850), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n880), .A2(new_n883), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT101), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n868), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n867), .A2(new_n843), .A3(KEYINPUT101), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n441), .A2(new_n879), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n621), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n207), .B2(new_n666), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n878), .A2(new_n893), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n794), .B1(new_n895), .B2(new_n896), .ZN(G367));
  NAND2_X1  g0697(.A1(new_n630), .A2(new_n631), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n570), .A2(new_n615), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n568), .A2(new_n572), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n598), .A2(new_n615), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT42), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n900), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT103), .Z(new_n905));
  AOI21_X1  g0705(.A(new_n598), .B1(new_n905), .B2(new_n632), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n903), .B1(new_n615), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n590), .A2(new_n624), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n597), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n658), .B2(new_n908), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT102), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n912));
  OR3_X1    g0712(.A1(new_n907), .A2(KEYINPUT104), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT104), .B1(new_n907), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n907), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n629), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(KEYINPUT105), .A3(new_n905), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n905), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n920), .B(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n636), .B(KEYINPUT41), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n633), .A2(new_n904), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT45), .Z(new_n928));
  NOR2_X1   g0728(.A1(new_n633), .A2(new_n904), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(new_n918), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT107), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT106), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n628), .B2(new_n631), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n898), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(KEYINPUT106), .B2(new_n898), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(new_n622), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n664), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n932), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n933), .B2(new_n939), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n926), .B1(new_n941), .B2(new_n664), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n925), .B1(new_n942), .B2(new_n668), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n728), .B1(new_n211), .B2(new_n429), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n734), .B2(new_n246), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n676), .A2(new_n772), .B1(new_n679), .B2(new_n202), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n287), .B(new_n946), .C1(G137), .C2(new_n700), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n708), .A2(new_n290), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G143), .A2(new_n685), .B1(new_n687), .B2(G159), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n694), .A2(G68), .B1(new_n721), .B2(G58), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n707), .A2(new_n459), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n700), .A2(G317), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n679), .B2(new_n765), .C1(new_n443), .C2(new_n676), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n688), .A2(new_n760), .B1(new_n513), .B2(new_n693), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n732), .B1(new_n770), .B2(new_n714), .ZN(new_n956));
  OR4_X1    g0756(.A1(new_n952), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT108), .B1(new_n690), .B2(new_n457), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n951), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT109), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n741), .B(new_n945), .C1(new_n962), .C2(new_n673), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n911), .B2(new_n743), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n943), .A2(new_n964), .ZN(G387));
  NAND2_X1  g0765(.A1(new_n938), .A2(new_n668), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT110), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n677), .A2(G317), .B1(new_n680), .B2(G303), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n770), .B2(new_n712), .C1(new_n714), .C2(new_n688), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT48), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n760), .B2(new_n690), .C1(new_n693), .C2(new_n765), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n969), .A2(new_n970), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT49), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT49), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n732), .B1(new_n697), .B2(new_n717), .C1(new_n707), .C2(new_n457), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT114), .Z(new_n978));
  NAND3_X1  g0778(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n687), .A2(new_n264), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n429), .B2(new_n693), .C1(new_n770), .C2(new_n698), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n676), .A2(new_n202), .B1(new_n679), .B2(new_n309), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n981), .A2(new_n732), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT113), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n690), .A2(new_n231), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT112), .B(G150), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n985), .B1(new_n700), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n952), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n983), .B(new_n988), .C1(new_n984), .C2(new_n987), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n674), .B1(new_n979), .B2(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n737), .A2(new_n637), .B1(new_n513), .B2(new_n635), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  AOI211_X1 g0792(.A(G45), .B(new_n637), .C1(G68), .C2(G77), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT50), .B1(new_n264), .B2(new_n202), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n264), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n734), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n243), .A2(new_n448), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n992), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n741), .B(new_n990), .C1(new_n728), .C2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n628), .B2(new_n743), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n967), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n636), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n664), .B2(new_n938), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n664), .B2(new_n938), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1002), .A2(new_n1005), .ZN(G393));
  AOI21_X1  g0806(.A(new_n1003), .B1(new_n932), .B2(new_n939), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n941), .A2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n932), .A2(new_n667), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n734), .A2(new_n251), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n729), .B1(G97), .B2(new_n635), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n741), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n293), .B1(new_n700), .B2(G322), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n709), .B(new_n1013), .C1(new_n690), .C2(new_n765), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT116), .Z(new_n1015));
  OAI22_X1  g0815(.A1(new_n693), .A2(new_n457), .B1(new_n679), .B2(new_n760), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G317), .A2(new_n685), .B1(new_n677), .B2(G311), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT52), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(G303), .C2(new_n687), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n732), .B1(G143), .B2(new_n700), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n763), .B(new_n1020), .C1(new_n309), .C2(new_n690), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G150), .A2(new_n685), .B1(new_n677), .B2(G159), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT51), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n694), .A2(G77), .B1(new_n680), .B2(new_n264), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n202), .B2(new_n688), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT115), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1015), .A2(new_n1019), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n727), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1012), .B1(new_n674), .B2(new_n1028), .C1(new_n905), .C2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1009), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1008), .A2(new_n1031), .ZN(G390));
  NAND2_X1  g0832(.A1(new_n870), .A2(new_n873), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n725), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n740), .B1(new_n264), .B2(new_n758), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n685), .A2(G128), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n698), .B2(new_n693), .C1(new_n688), .C2(new_n771), .ZN(new_n1037));
  INV_X1    g0837(.A(G132), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n293), .B1(new_n676), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT54), .B(G143), .ZN(new_n1040));
  INV_X1    g0840(.A(G125), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n679), .A2(new_n1040), .B1(new_n697), .B2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1037), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n721), .A2(new_n986), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT53), .Z(new_n1045));
  OAI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(new_n202), .C2(new_n707), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n685), .A2(G283), .B1(new_n680), .B2(G97), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n513), .B2(new_n688), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT118), .Z(new_n1049));
  OAI21_X1  g0849(.A(new_n287), .B1(new_n697), .B2(new_n760), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G116), .B2(new_n677), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n694), .A2(G77), .B1(new_n721), .B2(G87), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n776), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1046), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1035), .B1(new_n1054), .B2(new_n673), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1034), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n802), .A2(new_n871), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1033), .A2(new_n1057), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n879), .A2(new_n671), .A3(new_n750), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n798), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT117), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n867), .A2(KEYINPUT101), .A3(new_n843), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT101), .B1(new_n867), .B2(new_n843), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n624), .B(new_n750), .C1(new_n659), .C2(new_n661), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n800), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n872), .B1(new_n1066), .B2(new_n798), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1061), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  AND4_X1   g0868(.A1(new_n1061), .A2(new_n887), .A3(new_n888), .A4(new_n1067), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1058), .B(new_n1060), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1064), .A2(new_n1061), .A3(new_n1067), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n887), .A2(new_n888), .A3(new_n1067), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT117), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1071), .A2(new_n1073), .B1(new_n1033), .B2(new_n1057), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n879), .A2(G330), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n750), .A3(new_n798), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1070), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1056), .B1(new_n1078), .B2(new_n667), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1076), .A2(new_n441), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n876), .A2(new_n586), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1077), .B1(new_n798), .B2(new_n1059), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n801), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n797), .B(new_n796), .C1(new_n1075), .C2(new_n751), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1060), .A2(new_n1084), .A3(new_n800), .A4(new_n1065), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1081), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1003), .B1(new_n1078), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1070), .B(new_n1086), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1079), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G378));
  NAND2_X1  g0891(.A1(new_n889), .A2(G330), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n841), .A2(new_n844), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT40), .B1(new_n1093), .B2(new_n881), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n272), .A2(new_n810), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n308), .B(new_n1095), .Z(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1092), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(G330), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1064), .B2(new_n885), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1098), .B1(new_n1102), .B2(new_n884), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n875), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n847), .A2(new_n854), .A3(new_n874), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1099), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(new_n884), .A3(new_n1098), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1104), .A2(KEYINPUT119), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1105), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT119), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1081), .B(KEYINPUT120), .Z(new_n1113));
  NAND2_X1  g0913(.A1(new_n1089), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1109), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT57), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1003), .B1(new_n1118), .B2(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1109), .A2(new_n668), .A3(new_n1112), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1098), .A2(new_n725), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n669), .B1(new_n758), .B2(G50), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n688), .A2(new_n1038), .B1(new_n770), .B2(new_n1041), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n677), .A2(G128), .B1(new_n680), .B2(G137), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n690), .B2(new_n1040), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(G150), .C2(new_n694), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n708), .A2(G159), .ZN(new_n1131));
  AOI211_X1 g0931(.A(G33), .B(G41), .C1(new_n700), .C2(G124), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n676), .A2(new_n513), .B1(new_n679), .B2(new_n429), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n732), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(G41), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1134), .B(new_n1137), .C1(G283), .C2(new_n700), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n708), .A2(G58), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n985), .B1(G68), .B2(new_n694), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G97), .A2(new_n687), .B1(new_n685), .B2(G116), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT58), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1137), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1133), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1123), .B1(new_n1147), .B2(new_n673), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1122), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1121), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1120), .A2(new_n1150), .ZN(G375));
  AND2_X1   g0951(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1081), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n926), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n1154), .A3(new_n1087), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n740), .B1(G68), .B2(new_n758), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n679), .A2(new_n513), .B1(new_n697), .B2(new_n443), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n293), .B(new_n1157), .C1(G283), .C2(new_n677), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n708), .A2(G77), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n430), .A2(new_n694), .B1(new_n687), .B2(G116), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n685), .A2(G294), .B1(new_n721), .B2(G97), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT121), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n694), .A2(G50), .B1(new_n721), .B2(G159), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1038), .B2(new_n770), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1135), .B1(new_n688), .B2(new_n1040), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n700), .A2(G128), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n772), .B2(new_n679), .C1(new_n771), .C2(new_n676), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1162), .A2(new_n1163), .B1(new_n1169), .B2(new_n1139), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1163), .B2(new_n1162), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1156), .B1(new_n1171), .B2(new_n673), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT122), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n798), .B2(new_n726), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1152), .B2(new_n667), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1155), .A2(new_n1176), .ZN(G381));
  NAND3_X1  g0977(.A1(new_n1002), .A2(new_n745), .A3(new_n1005), .ZN(new_n1178));
  OR4_X1    g0978(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1178), .ZN(new_n1179));
  OR4_X1    g0979(.A1(G387), .A2(new_n1179), .A3(G375), .A4(G378), .ZN(G407));
  NAND2_X1  g0980(.A1(new_n614), .A2(G213), .ZN(new_n1181));
  OR3_X1    g0981(.A1(G375), .A2(G378), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(G407), .A2(G213), .A3(new_n1182), .ZN(G409));
  NAND2_X1  g0983(.A1(new_n1087), .A2(new_n636), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT125), .B1(new_n1152), .B2(new_n1081), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT60), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT60), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1184), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n784), .B1(new_n1188), .B2(new_n1175), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1185), .A2(KEYINPUT60), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1185), .A2(KEYINPUT60), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G384), .B(new_n1176), .C1(new_n1192), .C2(new_n1184), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1189), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1120), .A2(G378), .A3(new_n1150), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n667), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1149), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT123), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n668), .B1(new_n1200), .B2(new_n1110), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT123), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(new_n1149), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1109), .A2(new_n1114), .A3(new_n1154), .A4(new_n1112), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1199), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(KEYINPUT124), .A3(new_n1090), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1196), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT124), .B1(new_n1205), .B2(new_n1090), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1181), .B(new_n1195), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT62), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1181), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n614), .A2(G213), .A3(G2897), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1189), .A2(new_n1193), .A3(KEYINPUT126), .A4(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1189), .A2(new_n1193), .A3(KEYINPUT126), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1212), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT126), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1211), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT61), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1205), .A2(new_n1090), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT124), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n1206), .A3(new_n1196), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n1181), .A4(new_n1195), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1210), .A2(new_n1219), .A3(new_n1220), .A4(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n943), .A2(new_n964), .A3(G390), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G390), .B1(new_n943), .B2(new_n964), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1178), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n745), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1229), .A2(new_n1230), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1230), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1228), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1227), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT63), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1237), .B1(new_n1209), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT61), .B1(new_n1211), .B2(new_n1218), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n1239), .C2(new_n1209), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1238), .A2(new_n1242), .ZN(G405));
  NAND2_X1  g1043(.A1(G375), .A2(new_n1090), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1196), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1195), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1237), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT127), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1246), .A2(new_n1237), .A3(new_n1247), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1250), .A2(new_n1252), .ZN(G402));
endmodule


