//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n207), .A2(KEYINPUT76), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT76), .ZN(new_n209));
  XNOR2_X1  g008(.A(G197gat), .B(G204gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n203), .B1(new_n213), .B2(KEYINPUT29), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n216), .B(KEYINPUT80), .C1(KEYINPUT2), .C2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G141gat), .ZN(new_n221));
  INV_X1    g020(.A(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G148gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT2), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n219), .B1(new_n224), .B2(new_n215), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT81), .B(G141gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n221), .B1(new_n226), .B2(new_n220), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G155gat), .ZN(new_n229));
  INV_X1    g028(.A(G162gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT2), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT82), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n233), .B(KEYINPUT2), .C1(new_n229), .C2(new_n230), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n234), .A3(new_n215), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n218), .B(new_n225), .C1(new_n228), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n228), .A2(new_n235), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n218), .A2(new_n225), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(new_n203), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT29), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n213), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G228gat), .ZN(new_n245));
  INV_X1    g044(.A(G233gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n237), .A2(new_n243), .A3(G228gat), .A4(G233gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n202), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT90), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n202), .A3(new_n248), .ZN(new_n251));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G50gat), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(KEYINPUT90), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n251), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(new_n249), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n255), .B(KEYINPUT89), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n259), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G113gat), .ZN(new_n266));
  INV_X1    g065(.A(G113gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G120gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT1), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G127gat), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n270), .A2(KEYINPUT72), .A3(G134gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n269), .A2(KEYINPUT73), .A3(new_n273), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT73), .B1(new_n269), .B2(new_n273), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT4), .B1(new_n280), .B2(new_n236), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n269), .A2(new_n273), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n284), .A2(new_n277), .B1(new_n275), .B2(new_n272), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n285), .A2(new_n238), .A3(new_n239), .A4(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n281), .A2(new_n287), .A3(KEYINPUT85), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT85), .B1(new_n281), .B2(new_n287), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n277), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n236), .A2(KEYINPUT3), .B1(new_n291), .B2(new_n276), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n240), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n280), .B(new_n236), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(new_n296), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(KEYINPUT39), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G1gat), .B(G29gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT0), .ZN(new_n302));
  XNOR2_X1  g101(.A(G57gat), .B(G85gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(KEYINPUT39), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n294), .A2(new_n305), .A3(new_n296), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n300), .A2(KEYINPUT40), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT83), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n281), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n287), .A2(new_n308), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n295), .B(new_n293), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n298), .B2(new_n296), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n313), .ZN(new_n316));
  AOI211_X1 g115(.A(new_n296), .B(new_n316), .C1(new_n292), .C2(new_n240), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT86), .B1(new_n290), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n281), .A2(new_n287), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n281), .A2(new_n287), .A3(KEYINPUT85), .ZN(new_n322));
  AND4_X1   g121(.A1(KEYINPUT86), .A2(new_n317), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n315), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n304), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT40), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n300), .A2(new_n304), .A3(new_n306), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331));
  NOR3_X1   g130(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  AND2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  OAI22_X1  g137(.A1(new_n332), .A2(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G183gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT69), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n345));
  AOI21_X1  g144(.A(G190gat), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n338), .A2(KEYINPUT28), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n343), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT27), .B(G183gat), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n353), .A2(KEYINPUT70), .A3(KEYINPUT28), .A4(new_n338), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n339), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT71), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n347), .A2(new_n348), .B1(new_n352), .B2(new_n354), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT71), .B1(new_n359), .B2(new_n339), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT24), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n337), .A2(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n338), .A2(G183gat), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT65), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT65), .ZN(new_n370));
  XNOR2_X1  g169(.A(G183gat), .B(G190gat), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n370), .B(new_n367), .C1(new_n371), .C2(new_n363), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374));
  INV_X1    g173(.A(G169gat), .ZN(new_n375));
  INV_X1    g174(.A(G176gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n335), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT66), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT66), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n382), .A3(new_n335), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n362), .B1(new_n373), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT67), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n382), .B1(new_n379), .B2(new_n335), .ZN(new_n388));
  AOI211_X1 g187(.A(KEYINPUT66), .B(new_n334), .C1(new_n377), .C2(new_n378), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n369), .A2(new_n372), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(KEYINPUT67), .A3(new_n362), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n362), .B1(new_n335), .B2(KEYINPUT68), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n379), .B(new_n395), .C1(KEYINPUT68), .C2(new_n335), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n367), .B1(new_n371), .B2(new_n363), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n361), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT77), .B(new_n331), .C1(new_n400), .C2(KEYINPUT29), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT77), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT67), .B1(new_n392), .B2(new_n362), .ZN(new_n403));
  AOI211_X1 g202(.A(new_n386), .B(KEYINPUT25), .C1(new_n390), .C2(new_n391), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n358), .A2(new_n360), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n331), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n356), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT78), .B1(new_n411), .B2(new_n408), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n413), .B(new_n331), .C1(new_n405), .C2(new_n410), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n401), .B(new_n409), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n213), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n400), .B2(new_n331), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n398), .B1(new_n387), .B2(new_n393), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT79), .B(new_n408), .C1(new_n419), .C2(new_n361), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n213), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n411), .A2(new_n241), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n331), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n425), .A3(new_n429), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n416), .A2(new_n434), .A3(new_n425), .A4(new_n429), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n330), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n415), .A2(new_n422), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n213), .A3(new_n424), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT37), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT91), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n415), .A2(new_n422), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT37), .A4(new_n438), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n429), .B1(new_n416), .B2(new_n425), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n430), .A2(KEYINPUT37), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n440), .B(new_n443), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n444), .A2(new_n445), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n446), .A2(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n317), .A2(new_n321), .A3(new_n322), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n290), .A2(KEYINPUT86), .A3(new_n317), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n453), .A2(new_n454), .B1(new_n312), .B2(new_n314), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n304), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT92), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT6), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n324), .B2(new_n325), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(new_n456), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT92), .B1(new_n326), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n432), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n264), .B(new_n436), .C1(new_n450), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT64), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n285), .B1(new_n419), .B2(new_n361), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n405), .A2(new_n406), .A3(new_n280), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT34), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n468), .A2(new_n467), .A3(new_n469), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n476));
  XOR2_X1   g275(.A(KEYINPUT74), .B(KEYINPUT33), .Z(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G15gat), .B(G43gat), .Z(new_n479));
  XNOR2_X1  g278(.A(G71gat), .B(G99gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n476), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n481), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n475), .B(KEYINPUT32), .C1(new_n477), .C2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT75), .B(new_n474), .C1(new_n482), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT75), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n472), .B2(new_n473), .ZN(new_n488));
  INV_X1    g287(.A(new_n467), .ZN(new_n489));
  INV_X1    g288(.A(new_n469), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n280), .B1(new_n405), .B2(new_n406), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT34), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n470), .A2(new_n471), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT75), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n478), .A3(new_n481), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n488), .A2(new_n495), .A3(new_n484), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n486), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n486), .A2(KEYINPUT36), .A3(new_n497), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n460), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n456), .A2(KEYINPUT87), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n326), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n456), .A2(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n416), .A2(new_n425), .A3(new_n429), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n510), .A2(new_n444), .A3(new_n434), .ZN(new_n511));
  INV_X1    g310(.A(new_n435), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n264), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n264), .A2(new_n498), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT35), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n433), .A2(new_n435), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n264), .A4(new_n498), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n465), .A2(new_n515), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(G15gat), .A2(G22gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(G15gat), .A2(G22gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT16), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT94), .ZN(new_n527));
  INV_X1    g326(.A(G8gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n522), .A2(G1gat), .A3(new_n523), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n527), .A2(new_n528), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n539));
  AOI21_X1  g338(.A(G36gat), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n540), .A2(KEYINPUT15), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546));
  INV_X1    g345(.A(G43gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(G50gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n540), .B2(new_n542), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n543), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n550), .B(new_n544), .C1(new_n540), .C2(new_n542), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n535), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(KEYINPUT17), .A3(new_n553), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  INV_X1    g356(.A(G36gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n539), .ZN(new_n559));
  NOR2_X1   g358(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n549), .A3(new_n541), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n561), .A2(new_n541), .B1(new_n549), .B2(new_n548), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(new_n544), .ZN(new_n564));
  INV_X1    g363(.A(new_n553), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n557), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n556), .A2(new_n566), .B1(new_n533), .B2(new_n534), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n555), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n556), .A2(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n535), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT95), .ZN(new_n572));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n569), .A2(new_n572), .A3(KEYINPUT18), .A4(new_n573), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n535), .B(new_n554), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n573), .B(KEYINPUT13), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G197gat), .ZN(new_n583));
  XOR2_X1   g382(.A(KEYINPUT11), .B(G169gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT12), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n576), .A2(new_n586), .A3(new_n577), .A4(new_n580), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n521), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G64gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT96), .B1(new_n593), .B2(G57gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n595));
  INV_X1    g394(.A(G57gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(G64gat), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n594), .B(new_n597), .C1(new_n596), .C2(G64gat), .ZN(new_n598));
  OR2_X1    g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT97), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n598), .A2(new_n602), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G57gat), .B(G64gat), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n600), .B(new_n599), .C1(new_n608), .C2(new_n605), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n270), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n535), .B1(new_n611), .B2(new_n610), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT98), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n229), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n619), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n617), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT7), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT100), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G99gat), .ZN(new_n632));
  INV_X1    g431(.A(G106gat), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT8), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n631), .A2(KEYINPUT101), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT101), .B1(new_n631), .B2(new_n634), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n625), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G99gat), .B(G106gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n638), .B(new_n625), .C1(new_n635), .C2(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n570), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(KEYINPUT99), .Z(new_n648));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n643), .B(new_n651), .C1(new_n554), .C2(new_n642), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n644), .A2(new_n645), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n649), .ZN(new_n655));
  XOR2_X1   g454(.A(G134gat), .B(G162gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n654), .B2(new_n658), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(G120gat), .B(G148gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT104), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n631), .A2(new_n634), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n631), .A2(KEYINPUT101), .A3(new_n634), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n638), .B1(new_n671), .B2(new_n625), .ZN(new_n672));
  INV_X1    g471(.A(new_n641), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n610), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n675));
  INV_X1    g474(.A(new_n610), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n640), .A2(new_n676), .A3(new_n641), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n640), .A2(new_n676), .A3(KEYINPUT10), .A4(new_n641), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G230gat), .A2(G233gat), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT105), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683));
  INV_X1    g482(.A(new_n681), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n683), .B(new_n684), .C1(new_n678), .C2(new_n679), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n681), .B1(new_n674), .B2(new_n677), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n666), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n680), .A2(new_n681), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT103), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n680), .A2(new_n691), .A3(new_n681), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n687), .A2(new_n666), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n623), .A2(new_n662), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n509), .B(KEYINPUT106), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n592), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G1gat), .ZN(G1324gat));
  NOR4_X1   g500(.A1(new_n521), .A2(new_n519), .A3(new_n591), .A4(new_n697), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n528), .B2(new_n702), .ZN(new_n705));
  MUX2_X1   g504(.A(new_n704), .B(new_n705), .S(KEYINPUT42), .Z(G1325gat));
  NAND3_X1  g505(.A1(new_n592), .A2(new_n502), .A3(new_n698), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G15gat), .ZN(new_n708));
  INV_X1    g507(.A(new_n498), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G15gat), .A3(new_n697), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n592), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(G1326gat));
  NAND3_X1  g511(.A1(new_n592), .A2(new_n514), .A3(new_n698), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(G1327gat));
  INV_X1    g518(.A(new_n623), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n696), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n662), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n592), .A2(new_n537), .A3(new_n699), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n486), .A2(KEYINPUT36), .A3(new_n497), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT36), .B1(new_n486), .B2(new_n497), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n513), .A2(new_n514), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n440), .A2(new_n443), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n444), .A2(new_n445), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n447), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n448), .A2(new_n449), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n464), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n436), .A2(new_n264), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n727), .B(new_n728), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n517), .A2(new_n520), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT44), .B1(new_n737), .B2(new_n661), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n739), .B(new_n662), .C1(new_n735), .C2(new_n736), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n721), .A2(new_n591), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n741), .A2(new_n699), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n724), .B1(new_n537), .B2(new_n743), .ZN(G1328gat));
  INV_X1    g543(.A(new_n519), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n592), .A2(new_n558), .A3(new_n745), .A4(new_n722), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT46), .Z(new_n747));
  OAI21_X1  g546(.A(new_n739), .B1(new_n521), .B2(new_n662), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n433), .A2(new_n435), .B1(new_n508), .B2(new_n507), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n727), .B1(new_n749), .B2(new_n264), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n732), .ZN(new_n751));
  INV_X1    g550(.A(new_n464), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n734), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n745), .A2(new_n516), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n519), .A2(new_n509), .A3(new_n264), .A4(new_n498), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n756), .A2(new_n518), .B1(new_n757), .B2(KEYINPUT35), .ZN(new_n758));
  OAI211_X1 g557(.A(KEYINPUT44), .B(new_n661), .C1(new_n755), .C2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n748), .A2(new_n745), .A3(new_n759), .A4(new_n742), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n558), .B1(new_n760), .B2(KEYINPUT108), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(KEYINPUT108), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n762), .ZN(G1329gat));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n502), .A3(new_n759), .A4(new_n742), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G43gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n592), .A2(new_n547), .A3(new_n498), .A4(new_n722), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(KEYINPUT47), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1330gat));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n514), .A3(new_n759), .A4(new_n742), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G50gat), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT48), .B1(new_n773), .B2(KEYINPUT109), .ZN(new_n774));
  INV_X1    g573(.A(G50gat), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n592), .A2(new_n775), .A3(new_n514), .A4(new_n722), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n773), .B(new_n776), .C1(KEYINPUT109), .C2(KEYINPUT48), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1331gat));
  NOR4_X1   g579(.A1(new_n720), .A2(new_n590), .A3(new_n661), .A4(new_n696), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n737), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n737), .A2(KEYINPUT110), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n699), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(new_n596), .ZN(G1332gat));
  NAND3_X1  g588(.A1(new_n784), .A2(new_n745), .A3(new_n785), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT49), .B(G64gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n784), .A2(new_n745), .A3(new_n785), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1333gat));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n502), .A3(new_n785), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G71gat), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n709), .A2(G71gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n785), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(KEYINPUT50), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1334gat));
  NOR2_X1   g608(.A1(new_n786), .A2(new_n264), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g610(.A1(new_n623), .A2(new_n590), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n696), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n741), .A2(new_n699), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n627), .A2(new_n629), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI211_X1 g616(.A(new_n662), .B(new_n813), .C1(new_n735), .C2(new_n736), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT51), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n737), .A2(new_n661), .A3(new_n812), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n696), .A2(new_n816), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n699), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n817), .A2(new_n825), .ZN(G1336gat));
  OAI21_X1  g625(.A(new_n821), .B1(new_n818), .B2(KEYINPUT112), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n820), .A2(new_n828), .A3(KEYINPUT51), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n519), .A2(G92gat), .A3(new_n696), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n748), .A2(new_n745), .A3(new_n759), .A4(new_n814), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G92gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(new_n823), .B2(new_n830), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1337gat));
  NAND4_X1  g637(.A1(new_n823), .A2(new_n632), .A3(new_n498), .A4(new_n695), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n741), .A2(new_n502), .A3(new_n814), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n632), .ZN(G1338gat));
  NAND4_X1  g640(.A1(new_n748), .A2(new_n514), .A3(new_n759), .A4(new_n814), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n633), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n741), .A2(KEYINPUT113), .A3(new_n514), .A4(new_n814), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n264), .A2(G106gat), .A3(new_n696), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT53), .B1(new_n823), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n827), .A2(new_n829), .A3(new_n847), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n842), .A2(G106gat), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT53), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(G1339gat));
  NOR2_X1   g652(.A1(new_n697), .A2(new_n590), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n678), .A2(new_n679), .A3(new_n684), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT114), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n678), .A2(new_n679), .A3(new_n857), .A4(new_n684), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(new_n690), .A3(KEYINPUT54), .A4(new_n692), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n689), .A2(new_n683), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n680), .A2(KEYINPUT105), .A3(new_n681), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n860), .A2(KEYINPUT55), .A3(new_n666), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n590), .A2(new_n865), .A3(new_n694), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867));
  AND4_X1   g666(.A1(KEYINPUT54), .A2(new_n859), .A3(new_n690), .A4(new_n692), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n864), .A2(new_n666), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n666), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n686), .B2(new_n862), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT55), .B1(new_n874), .B2(new_n860), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n866), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n573), .B1(new_n569), .B2(new_n572), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n578), .A2(new_n579), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n585), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n589), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n695), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n662), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n865), .A2(new_n881), .A3(new_n661), .A4(new_n694), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n871), .B(KEYINPUT55), .C1(new_n874), .C2(new_n860), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n854), .B1(new_n890), .B2(new_n720), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n514), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n699), .A2(new_n519), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n709), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n267), .A3(new_n591), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n891), .A2(new_n787), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n756), .A3(new_n590), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n267), .B2(new_n898), .ZN(G1340gat));
  OAI21_X1  g698(.A(G120gat), .B1(new_n895), .B2(new_n696), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(KEYINPUT116), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(KEYINPUT116), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(new_n756), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n695), .A2(new_n265), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT117), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n901), .A2(new_n902), .B1(new_n903), .B2(new_n905), .ZN(G1341gat));
  OAI21_X1  g705(.A(G127gat), .B1(new_n895), .B2(new_n720), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n623), .A2(new_n270), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n903), .B2(new_n908), .ZN(G1342gat));
  OR3_X1    g708(.A1(new_n903), .A2(G134gat), .A3(new_n662), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n911));
  OAI21_X1  g710(.A(G134gat), .B1(new_n895), .B2(new_n662), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G1343gat));
  AOI21_X1  g713(.A(new_n623), .B1(new_n884), .B2(new_n889), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT118), .B(new_n699), .C1(new_n915), .C2(new_n854), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n502), .A2(new_n264), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n885), .B1(new_n872), .B2(new_n876), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n590), .A2(new_n865), .A3(new_n694), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n887), .B2(new_n888), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n882), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n922), .B2(new_n662), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n923), .A2(new_n623), .B1(new_n590), .B2(new_n697), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT118), .B1(new_n924), .B2(new_n699), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT119), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n891), .B2(new_n787), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n917), .A4(new_n916), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n591), .A2(G141gat), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n926), .A2(new_n930), .A3(new_n519), .A4(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n917), .A3(new_n916), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n745), .B1(new_n935), .B2(KEYINPUT119), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n936), .A2(KEYINPUT120), .A3(new_n931), .A4(new_n930), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n699), .A2(new_n519), .A3(new_n727), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT57), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(new_n891), .B2(new_n264), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n514), .A2(KEYINPUT57), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n882), .B1(new_n866), .B2(new_n875), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n662), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n623), .B1(new_n944), .B2(new_n889), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n945), .B2(new_n854), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n938), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n590), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT58), .B1(new_n948), .B2(new_n226), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n937), .A3(new_n949), .ZN(new_n950));
  NOR4_X1   g749(.A1(new_n935), .A2(G141gat), .A3(new_n745), .A4(new_n591), .ZN(new_n951));
  INV_X1    g750(.A(new_n226), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n952), .B1(new_n947), .B2(new_n590), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT58), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n950), .A2(new_n954), .ZN(G1344gat));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n696), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n514), .B1(new_n945), .B2(new_n854), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(new_n959), .A3(new_n939), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n942), .B1(new_n915), .B2(new_n854), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n959), .B1(new_n958), .B2(new_n939), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n956), .B(new_n957), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G148gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n958), .A2(new_n939), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT121), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n967), .A2(new_n961), .A3(new_n960), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n957), .B1(new_n968), .B2(new_n956), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT59), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n220), .A2(KEYINPUT59), .ZN(new_n971));
  INV_X1    g770(.A(new_n947), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(new_n696), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n936), .A2(new_n220), .A3(new_n695), .A4(new_n930), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1345gat));
  OAI21_X1  g775(.A(G155gat), .B1(new_n972), .B2(new_n720), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n936), .A2(new_n930), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n623), .A2(new_n229), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(G1346gat));
  NOR3_X1   g779(.A1(new_n972), .A2(new_n230), .A3(new_n662), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n936), .A2(new_n661), .A3(new_n930), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n230), .ZN(G1347gat));
  NAND2_X1  g782(.A1(new_n787), .A2(new_n745), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n984), .A2(new_n709), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n892), .A2(new_n985), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n986), .A2(new_n375), .A3(new_n591), .ZN(new_n987));
  NOR4_X1   g786(.A1(new_n891), .A2(new_n519), .A3(new_n516), .A4(new_n699), .ZN(new_n988));
  AOI21_X1  g787(.A(G169gat), .B1(new_n988), .B2(new_n590), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n987), .A2(new_n989), .ZN(G1348gat));
  OAI21_X1  g789(.A(G176gat), .B1(new_n986), .B2(new_n696), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n988), .A2(new_n376), .A3(new_n695), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT123), .ZN(G1349gat));
  OAI21_X1  g793(.A(G183gat), .B1(new_n986), .B2(new_n720), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n988), .A2(new_n353), .A3(new_n623), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g796(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n998));
  XNOR2_X1  g797(.A(new_n997), .B(new_n998), .ZN(G1350gat));
  NAND3_X1  g798(.A1(new_n988), .A2(new_n338), .A3(new_n661), .ZN(new_n1000));
  OAI21_X1  g799(.A(G190gat), .B1(new_n986), .B2(new_n662), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n1001), .A2(KEYINPUT61), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n1001), .A2(KEYINPUT61), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(G1351gat));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n984), .A2(new_n502), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n968), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1005), .B1(new_n1007), .B2(new_n591), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(G197gat), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n1007), .A2(new_n1005), .A3(new_n591), .ZN(new_n1010));
  NAND4_X1  g809(.A1(new_n924), .A2(new_n745), .A3(new_n787), .A4(new_n917), .ZN(new_n1011));
  OR2_X1    g810(.A1(new_n591), .A2(G197gat), .ZN(new_n1012));
  OAI22_X1  g811(.A1(new_n1009), .A2(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(G1352gat));
  NOR3_X1   g812(.A1(new_n1011), .A2(G204gat), .A3(new_n696), .ZN(new_n1014));
  XNOR2_X1  g813(.A(new_n1014), .B(KEYINPUT62), .ZN(new_n1015));
  OAI21_X1  g814(.A(G204gat), .B1(new_n1007), .B2(new_n696), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(G1353gat));
  NOR3_X1   g816(.A1(new_n1011), .A2(G211gat), .A3(new_n720), .ZN(new_n1018));
  OAI211_X1 g817(.A(new_n623), .B(new_n1006), .C1(new_n962), .C2(new_n963), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1019), .B2(G211gat), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1019), .A2(G211gat), .ZN(new_n1023));
  INV_X1    g822(.A(KEYINPUT63), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1025), .A2(KEYINPUT126), .ZN(new_n1026));
  NOR2_X1   g825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1022), .B1(new_n1026), .B2(new_n1027), .ZN(G1354gat));
  AND3_X1   g827(.A1(new_n968), .A2(KEYINPUT127), .A3(new_n1006), .ZN(new_n1029));
  AOI21_X1  g828(.A(KEYINPUT127), .B1(new_n968), .B2(new_n1006), .ZN(new_n1030));
  NOR3_X1   g829(.A1(new_n1029), .A2(new_n1030), .A3(new_n662), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n661), .A2(new_n206), .ZN(new_n1032));
  OAI22_X1  g831(.A1(new_n1031), .A2(new_n206), .B1(new_n1011), .B2(new_n1032), .ZN(G1355gat));
endmodule


