//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G137), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n469), .B1(new_n462), .B2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n468), .B1(new_n472), .B2(G101), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  AOI211_X1 g049(.A(KEYINPUT69), .B(new_n474), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT70), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G125), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(new_n467), .C1(new_n473), .C2(new_n475), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n477), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  NOR2_X1   g063(.A1(new_n481), .A2(new_n466), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n466), .A2(G112), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n481), .B2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n465), .A2(KEYINPUT71), .A3(new_n466), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G136), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n497), .A2(KEYINPUT72), .A3(G136), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n493), .B1(new_n500), .B2(new_n501), .ZN(G162));
  NAND2_X1  g077(.A1(KEYINPUT4), .A2(G138), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n463), .B2(new_n464), .ZN(new_n504));
  AND2_X1   g079(.A1(G102), .A2(G2104), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n466), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G126), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n507), .B1(new_n463), .B2(new_n464), .ZN(new_n508));
  AND2_X1   g083(.A1(G114), .A2(G2104), .ZN(new_n509));
  OAI21_X1  g084(.A(G2105), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(G138), .B(new_n466), .C1(new_n479), .C2(new_n480), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n506), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT73), .B1(new_n517), .B2(G50), .ZN(new_n518));
  AND4_X1   g093(.A1(KEYINPUT73), .A2(new_n516), .A3(G50), .A4(G543), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(new_n527), .A3(new_n516), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n523), .A2(new_n525), .B1(new_n522), .B2(G543), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n529), .A2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n517), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n528), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n535), .B(new_n536), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n532), .ZN(new_n546));
  INV_X1    g121(.A(new_n517), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT76), .B(G52), .Z(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n528), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n546), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n526), .A2(new_n527), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(KEYINPUT77), .A3(G651), .ZN(new_n560));
  INV_X1    g135(.A(new_n528), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G81), .B1(G43), .B2(new_n517), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g141(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n567));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND3_X1  g145(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n554), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n530), .A2(new_n581), .A3(new_n516), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(G91), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G299));
  INV_X1    g161(.A(G168), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  OR2_X1    g163(.A1(new_n530), .A2(G74), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G49), .B2(new_n517), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n580), .A2(G87), .A3(new_n582), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G288));
  NAND3_X1  g167(.A1(new_n526), .A2(G61), .A3(new_n527), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G48), .B2(new_n517), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n580), .A2(G86), .A3(new_n582), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n554), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(KEYINPUT80), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(KEYINPUT80), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n561), .A2(G85), .B1(G47), .B2(new_n517), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(G290));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(G301), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n554), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n615), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n580), .A2(G92), .A3(new_n582), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT82), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n580), .A2(new_n620), .A3(G92), .A4(new_n582), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n619), .B1(new_n618), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g201(.A(KEYINPUT83), .B(new_n616), .C1(new_n622), .C2(new_n623), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT84), .Z(new_n629));
  AOI21_X1  g204(.A(new_n612), .B1(new_n629), .B2(new_n611), .ZN(G284));
  AOI21_X1  g205(.A(new_n612), .B1(new_n629), .B2(new_n611), .ZN(G321));
  OAI21_X1  g206(.A(KEYINPUT85), .B1(new_n585), .B2(G868), .ZN(new_n632));
  NOR2_X1   g207(.A1(G168), .A2(new_n611), .ZN(new_n633));
  MUX2_X1   g208(.A(new_n632), .B(KEYINPUT85), .S(new_n633), .Z(G297));
  MUX2_X1   g209(.A(new_n632), .B(KEYINPUT85), .S(new_n633), .Z(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n629), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n629), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n472), .A2(new_n465), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT13), .Z(new_n644));
  INV_X1    g219(.A(G2100), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n497), .A2(G135), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(KEYINPUT86), .ZN(new_n650));
  INV_X1    g225(.A(G111), .ZN(new_n651));
  AOI22_X1  g226(.A1(new_n649), .A2(KEYINPUT86), .B1(new_n651), .B2(G2105), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n489), .A2(G123), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n646), .A2(new_n647), .A3(new_n655), .ZN(G156));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n660), .B(new_n666), .Z(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT87), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT17), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2084), .B(G2090), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n673), .B2(new_n675), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n674), .B2(new_n675), .ZN(new_n679));
  INV_X1    g254(.A(new_n675), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(new_n676), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT18), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1956), .B(G2474), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(new_n692), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT20), .Z(new_n696));
  AOI211_X1 g271(.A(new_n694), .B(new_n696), .C1(new_n689), .C2(new_n693), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT89), .ZN(new_n698));
  XOR2_X1   g273(.A(G1981), .B(G1986), .Z(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n698), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  XOR2_X1   g280(.A(KEYINPUT96), .B(KEYINPUT36), .Z(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G24), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G290), .B2(G16), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G1986), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G1986), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT90), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(KEYINPUT90), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT91), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n497), .A2(G131), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(G107), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G2105), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n489), .B2(G119), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n716), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n718), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n712), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G22), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n731), .A2(KEYINPUT95), .A3(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(KEYINPUT95), .B1(new_n731), .B2(G16), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n732), .B(new_n733), .C1(G166), .C2(new_n707), .ZN(new_n734));
  INV_X1    g309(.A(G1971), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G16), .A2(G23), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT94), .Z(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G288), .B2(new_n707), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT33), .B(G1976), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n736), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  MUX2_X1   g318(.A(G6), .B(G305), .S(G16), .Z(new_n744));
  XOR2_X1   g319(.A(KEYINPUT32), .B(G1981), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT93), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n744), .B(new_n746), .Z(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n743), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n743), .B2(new_n747), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n706), .B1(new_n730), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n728), .B1(new_n710), .B2(new_n711), .ZN(new_n754));
  INV_X1    g329(.A(new_n706), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n754), .A2(new_n755), .A3(new_n750), .A4(new_n751), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n713), .A2(G32), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n495), .A2(G141), .A3(new_n496), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT102), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n472), .A2(G105), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT103), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n489), .A2(G129), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n757), .B1(new_n769), .B2(new_n713), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT27), .ZN(new_n771));
  INV_X1    g346(.A(G1996), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n725), .A2(G35), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G162), .B2(new_n725), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT29), .Z(new_n776));
  INV_X1    g351(.A(G2090), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n707), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n707), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT104), .B(G1966), .Z(new_n781));
  XOR2_X1   g356(.A(new_n780), .B(new_n781), .Z(new_n782));
  NOR3_X1   g357(.A1(new_n773), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n716), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT28), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n489), .A2(G128), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n497), .A2(G140), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n788), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n785), .B1(new_n793), .B2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2067), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n497), .A2(G139), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT25), .Z(new_n798));
  NAND2_X1  g373(.A1(G115), .A2(G2104), .ZN(new_n799));
  INV_X1    g374(.A(G127), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n481), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G2105), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n796), .B(new_n798), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G33), .B(new_n805), .S(G29), .Z(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(G2072), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n795), .B1(new_n807), .B2(KEYINPUT100), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(KEYINPUT100), .B2(new_n807), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n707), .A2(G5), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G301), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT105), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT31), .B(G11), .Z(new_n815));
  NOR2_X1   g390(.A1(new_n654), .A2(new_n716), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT30), .B(G28), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n815), .B(new_n816), .C1(new_n713), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n811), .A2(new_n812), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n716), .A2(G27), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G164), .B2(new_n716), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(G2078), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(G2078), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n818), .A2(new_n819), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n814), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT24), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(G34), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(G34), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n716), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n487), .B2(new_n713), .ZN(new_n830));
  INV_X1    g405(.A(G2084), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n564), .A2(G16), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G16), .B2(G19), .ZN(new_n834));
  INV_X1    g409(.A(G1341), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n776), .A2(new_n777), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n809), .A2(new_n825), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n806), .A2(G2072), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT101), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n830), .A2(new_n831), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT106), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n707), .A2(G20), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT107), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT23), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G299), .B2(G16), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G1956), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n834), .A2(new_n835), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n840), .A2(new_n842), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n838), .A2(new_n849), .ZN(new_n850));
  AND4_X1   g425(.A1(new_n753), .A2(new_n756), .A3(new_n783), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(G4), .A2(G16), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n629), .B2(G16), .ZN(new_n853));
  INV_X1    g428(.A(G1348), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n851), .A2(new_n855), .ZN(G311));
  AND3_X1   g431(.A1(new_n851), .A2(KEYINPUT108), .A3(new_n855), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT108), .B1(new_n851), .B2(new_n855), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(G150));
  AOI22_X1  g434(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n532), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n517), .A2(G55), .ZN(new_n862));
  INV_X1    g437(.A(G93), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n528), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  INV_X1    g443(.A(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n563), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n563), .A2(new_n869), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n629), .A2(G559), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n629), .B2(G559), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n873), .A3(new_n877), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n866), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n868), .B1(new_n886), .B2(new_n887), .ZN(G145));
  NAND2_X1  g463(.A1(new_n497), .A2(G142), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n466), .A2(G118), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n890), .A2(KEYINPUT112), .ZN(new_n891));
  OAI21_X1  g466(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n890), .B2(KEYINPUT112), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n891), .A2(new_n893), .B1(new_n489), .B2(G130), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n643), .ZN(new_n896));
  INV_X1    g471(.A(new_n724), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n793), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n805), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n769), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n768), .A2(new_n901), .A3(new_n805), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n514), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n514), .A3(new_n904), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n900), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n909), .A2(new_n905), .A3(new_n793), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n899), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT113), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n793), .B1(new_n909), .B2(new_n905), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n906), .A2(new_n900), .A3(new_n907), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n898), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n487), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n654), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n487), .B(KEYINPUT110), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n654), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G162), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n898), .B1(new_n913), .B2(new_n914), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(KEYINPUT113), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n916), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n911), .A2(new_n925), .A3(new_n915), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT114), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT114), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n916), .A2(new_n927), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(KEYINPUT115), .B(KEYINPUT40), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n937), .B(new_n938), .ZN(G395));
  INV_X1    g514(.A(G290), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(G288), .ZN(new_n941));
  INV_X1    g516(.A(G288), .ZN(new_n942));
  NAND2_X1  g517(.A1(G290), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(G166), .B(G305), .Z(new_n944));
  AND3_X1   g519(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n941), .B2(new_n943), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n947), .B(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n624), .A2(new_n585), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n624), .A2(new_n585), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(KEYINPUT41), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(KEYINPUT116), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n624), .A2(KEYINPUT116), .A3(new_n585), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n953), .B1(KEYINPUT41), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n629), .A2(new_n636), .A3(new_n874), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n874), .B1(new_n629), .B2(new_n636), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n960), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n958), .A3(new_n956), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n949), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n949), .B1(new_n963), .B2(new_n961), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n869), .A2(new_n611), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n967), .ZN(G331));
  NOR3_X1   g544(.A1(new_n871), .A2(new_n872), .A3(G171), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(G171), .B1(new_n871), .B2(new_n872), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(G168), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n872), .ZN(new_n974));
  AOI21_X1  g549(.A(G301), .B1(new_n974), .B2(new_n870), .ZN(new_n975));
  OAI21_X1  g550(.A(G286), .B1(new_n975), .B2(new_n970), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(new_n954), .A3(new_n951), .A4(new_n955), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n957), .B2(new_n977), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n945), .A2(new_n946), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n973), .A2(KEYINPUT41), .A3(new_n976), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n952), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n947), .B(new_n983), .C1(new_n956), .C2(new_n982), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n981), .A2(KEYINPUT43), .A3(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n979), .A2(new_n980), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT43), .B1(new_n986), .B2(new_n981), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT44), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n986), .B2(new_n981), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n956), .A2(KEYINPUT41), .ZN(new_n992));
  INV_X1    g567(.A(new_n953), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n977), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n973), .A2(new_n976), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n956), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n980), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AND4_X1   g572(.A1(new_n990), .A2(new_n997), .A3(new_n930), .A4(new_n984), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n989), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n988), .A2(new_n999), .ZN(G397));
  INV_X1    g575(.A(G2067), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n793), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n768), .B(G1996), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n897), .A2(new_n727), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT127), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1005), .A2(new_n1007), .B1(new_n1001), .B2(new_n900), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n514), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n484), .A2(G40), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n477), .A2(new_n486), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1008), .A2(new_n1017), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n897), .A2(new_n727), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1005), .A2(new_n1006), .A3(new_n1019), .ZN(new_n1020));
  OR3_X1    g595(.A1(G290), .A2(new_n1017), .A3(G1986), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT48), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1020), .A2(new_n1016), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1022), .B2(new_n1021), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1016), .B1(new_n1003), .B2(new_n768), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n1017), .B2(G1996), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1016), .A2(KEYINPUT46), .A3(new_n772), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1024), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1018), .B(new_n1031), .C1(new_n1025), .C2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g607(.A(G8), .B1(new_n529), .B2(new_n533), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT55), .B(G8), .C1(new_n529), .C2(new_n533), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n514), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT45), .B1(new_n514), .B2(new_n1009), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n477), .A2(new_n486), .A3(new_n1014), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1971), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n514), .A2(new_n1043), .A3(new_n1009), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n514), .B2(new_n1009), .ZN(new_n1045));
  NOR4_X1   g620(.A1(new_n1015), .A2(new_n1044), .A3(new_n1045), .A4(G2090), .ZN(new_n1046));
  OAI211_X1 g621(.A(G8), .B(new_n1037), .C1(new_n1042), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1010), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n514), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n735), .B1(new_n1053), .B2(new_n1015), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(new_n1041), .A3(new_n777), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(KEYINPUT118), .A3(G8), .A4(new_n1037), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1049), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1010), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1062), .A2(new_n477), .A3(new_n486), .A4(new_n1014), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n590), .A2(new_n591), .A3(G1976), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1061), .A2(new_n1063), .A3(G8), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n1015), .B2(new_n1010), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G288), .A2(new_n1060), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT52), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n1069));
  INV_X1    g644(.A(G1981), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n596), .A2(new_n597), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n517), .A2(G48), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n530), .A2(G86), .A3(new_n516), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n530), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1072), .B(new_n1073), .C1(new_n1074), .C2(new_n532), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G1981), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  OAI211_X1 g653(.A(G8), .B(new_n1063), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1069), .B(KEYINPUT49), .C1(new_n1071), .C2(new_n1076), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1065), .B(new_n1068), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1037), .B1(new_n1057), .B2(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1059), .A2(new_n1083), .A3(KEYINPUT125), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT125), .B1(new_n1059), .B2(new_n1083), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1956), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n514), .A2(new_n1043), .A3(new_n1009), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(new_n1090), .B2(new_n1015), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1040), .A2(new_n1041), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n579), .B2(new_n584), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n583), .A2(new_n574), .A3(new_n578), .A4(KEYINPUT57), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1055), .A2(new_n1041), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n854), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n466), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT68), .B1(new_n466), .B2(G2104), .ZN(new_n1102));
  OAI21_X1  g677(.A(G101), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT69), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n472), .A2(new_n468), .A3(G101), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n485), .B1(new_n1106), .B2(new_n467), .ZN(new_n1107));
  INV_X1    g682(.A(new_n486), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1109), .A2(new_n1001), .A3(new_n1014), .A4(new_n1062), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1100), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n628), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1097), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1098), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1015), .A2(new_n1045), .A3(new_n1044), .ZN(new_n1115));
  OAI211_X1 g690(.A(KEYINPUT60), .B(new_n1110), .C1(new_n1115), .C2(G1348), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1100), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n1110), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n628), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n626), .A2(new_n1116), .A3(new_n1117), .A4(new_n627), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1111), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n563), .B1(new_n1126), .B2(KEYINPUT59), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1053), .A2(G1996), .A3(new_n1015), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT58), .B(G1341), .Z(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1041), .B2(new_n1062), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1127), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1126), .A2(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1133), .B(new_n1127), .C1(new_n1128), .C2(new_n1131), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1098), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n1113), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1113), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1114), .B1(new_n1125), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G2078), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1040), .A2(new_n1041), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1146), .A2(new_n1147), .B1(new_n1115), .B2(G1961), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1149), .A3(new_n1147), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1148), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G301), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1145), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n487), .A2(new_n1038), .A3(new_n1156), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n812), .A2(new_n1099), .B1(new_n1157), .B2(new_n1013), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT54), .B(new_n1154), .C1(new_n1159), .C2(G301), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n781), .B1(new_n1053), .B2(new_n1015), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1055), .A2(new_n1041), .A3(new_n831), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1161), .A2(G286), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(G286), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1164));
  OAI211_X1 g739(.A(KEYINPUT51), .B(G8), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT51), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1161), .A2(G168), .A3(new_n1162), .ZN(new_n1167));
  INV_X1    g742(.A(G8), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1152), .ZN(new_n1171));
  OAI211_X1 g746(.A(G301), .B(new_n1158), .C1(new_n1171), .C2(new_n1150), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1153), .B2(G301), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT54), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1086), .A2(new_n1144), .A3(new_n1160), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n942), .A2(new_n1060), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT119), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1066), .B1(new_n1179), .B2(KEYINPUT49), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1080), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1177), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1071), .B(KEYINPUT120), .ZN(new_n1183));
  OAI211_X1 g758(.A(G8), .B(new_n1063), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(new_n1059), .B2(new_n1081), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1184), .B(KEYINPUT121), .C1(new_n1059), .C2(new_n1081), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1164), .A2(G8), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1059), .A2(new_n1083), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1059), .A2(new_n1083), .A3(new_n1189), .A4(KEYINPUT63), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1187), .A2(new_n1188), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1176), .A2(KEYINPUT126), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT126), .B1(new_n1176), .B2(new_n1194), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1153), .A2(G301), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1170), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1165), .A2(new_n1169), .A3(KEYINPUT62), .ZN(new_n1200));
  AND4_X1   g775(.A1(new_n1197), .A2(new_n1086), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1195), .A2(new_n1196), .A3(new_n1201), .ZN(new_n1202));
  XOR2_X1   g777(.A(G290), .B(G1986), .Z(new_n1203));
  INV_X1    g778(.A(new_n1020), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1017), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1032), .B1(new_n1202), .B2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(G319), .ZN(new_n1208));
  NOR4_X1   g782(.A1(G229), .A2(new_n1208), .A3(G401), .A4(G227), .ZN(new_n1209));
  OAI211_X1 g783(.A(new_n937), .B(new_n1209), .C1(new_n991), .C2(new_n998), .ZN(G225));
  INV_X1    g784(.A(G225), .ZN(G308));
endmodule


