//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n549, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G219), .A2(G218), .A3(G220), .A4(G221), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT70), .B(G2104), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G101), .A3(new_n475), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n472), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  XNOR2_X1  g056(.A(new_n471), .B(KEYINPUT71), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n468), .B1(new_n477), .B2(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n475), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n483), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OR2_X1    g066(.A1(new_n475), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n484), .A2(new_n498), .A3(G138), .A4(new_n475), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n467), .A2(G138), .A3(new_n475), .A4(new_n469), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT72), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n473), .A2(new_n503), .A3(G138), .A4(new_n475), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n497), .B1(new_n502), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n507), .B(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n508), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n508), .A2(G543), .A3(new_n510), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(new_n506), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n516), .A2(new_n519), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(new_n515), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n513), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n524), .A2(new_n525), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AOI22_X1  g107(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n506), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n534), .B1(new_n514), .B2(new_n535), .C1(new_n536), .C2(new_n517), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n506), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n541), .A2(new_n517), .B1(new_n514), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT75), .B1(new_n517), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n507), .A2(KEYINPUT73), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n507), .A2(KEYINPUT73), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n556), .A2(new_n557), .B1(new_n509), .B2(G651), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n558), .A2(new_n559), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(KEYINPUT9), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n513), .A2(G65), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n506), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n515), .B2(G91), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  OAI211_X1 g141(.A(KEYINPUT75), .B(new_n566), .C1(new_n517), .C2(new_n554), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n561), .A2(new_n565), .A3(new_n567), .ZN(G299));
  NAND2_X1  g143(.A1(new_n515), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n518), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND3_X1  g147(.A1(new_n558), .A2(G48), .A3(G543), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n558), .A2(G86), .A3(new_n513), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n506), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n518), .A2(G47), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n515), .A2(G85), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n506), .C2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  INV_X1    g157(.A(G92), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT76), .B1(new_n514), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n558), .A2(new_n585), .A3(G92), .A4(new_n513), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n584), .A2(KEYINPUT10), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT10), .B1(new_n584), .B2(new_n586), .ZN(new_n588));
  INV_X1    g163(.A(G54), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n517), .A2(new_n589), .B1(new_n506), .B2(new_n590), .ZN(new_n591));
  NOR3_X1   g166(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  XNOR2_X1  g173(.A(KEYINPUT77), .B(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(G860), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT78), .ZN(G148));
  NAND2_X1  g176(.A1(new_n592), .A2(new_n599), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n547), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n473), .A2(new_n475), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n477), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(G2100), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n482), .A2(G135), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n475), .A2(G111), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(KEYINPUT80), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n613), .B2(KEYINPUT80), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n486), .A2(G123), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(G2096), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n611), .A2(new_n619), .A3(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT82), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2430), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n628), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  AND2_X1   g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(G14), .B1(new_n632), .B2(new_n635), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT83), .Z(new_n640));
  NOR2_X1   g215(.A1(G2072), .A2(G2078), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n444), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n642), .B(KEYINPUT17), .Z(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n646), .C1(new_n647), .C2(new_n640), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n642), .A2(new_n639), .A3(new_n645), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n640), .A3(new_n645), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT84), .B(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT86), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n656), .A2(new_n657), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(new_n658), .ZN(new_n666));
  MUX2_X1   g241(.A(new_n666), .B(new_n665), .S(new_n662), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1991), .B(G1996), .Z(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  XOR2_X1   g245(.A(G1981), .B(G1986), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G229));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT33), .B(G1976), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n677), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1971), .ZN(new_n685));
  NOR2_X1   g260(.A1(G6), .A2(G16), .ZN(new_n686));
  INV_X1    g261(.A(G305), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(G16), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  NOR3_X1   g265(.A1(new_n682), .A2(new_n685), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  MUX2_X1   g269(.A(G24), .B(G290), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(G1986), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n486), .A2(G119), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g275(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n701));
  OAI221_X1 g276(.A(G2104), .B1(G107), .B2(new_n475), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n482), .A2(G131), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n705), .S(G29), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n693), .A2(new_n694), .A3(new_n696), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT36), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n677), .A2(G20), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT23), .Z(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G299), .B2(G16), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT100), .B(G1956), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n547), .A2(G16), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G16), .B2(G19), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT90), .B(G1341), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n482), .A2(G141), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT26), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n478), .A2(G105), .A3(new_n475), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n723), .B(new_n724), .C1(new_n486), .C2(G129), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(G32), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT30), .B(G28), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT31), .A2(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n734), .A2(new_n728), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G34), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n738), .B2(KEYINPUT24), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(KEYINPUT24), .B2(new_n738), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n480), .B2(new_n728), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n737), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n742), .B2(new_n741), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n618), .A2(new_n728), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT98), .Z(new_n746));
  NAND4_X1  g321(.A1(new_n732), .A2(new_n733), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n677), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n677), .ZN(new_n749));
  INV_X1    g324(.A(G1966), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n677), .A2(G5), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G171), .B2(new_n677), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n755), .C1(new_n714), .C2(new_n713), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n747), .A2(new_n756), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n720), .B(new_n757), .C1(new_n717), .C2(new_n719), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n728), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n760), .B(new_n761), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n482), .A2(G140), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n475), .A2(G116), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n486), .A2(G128), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g343(.A1(new_n768), .A2(KEYINPUT91), .A3(G29), .ZN(new_n769));
  AOI21_X1  g344(.A(KEYINPUT91), .B1(new_n768), .B2(G29), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n762), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT94), .B(G2067), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(new_n475), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT25), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n775), .B(new_n777), .C1(new_n482), .C2(G139), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  NOR2_X1   g354(.A1(G29), .A2(G33), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT95), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT96), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n442), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n728), .A2(G35), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n728), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(G2090), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G2090), .B2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n783), .A2(new_n442), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT97), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n592), .A2(G16), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G4), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(G1348), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G27), .A2(G29), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G164), .B2(G29), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT99), .B(G2078), .Z(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n793), .A2(new_n794), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n795), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n789), .A2(new_n791), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n710), .A2(new_n758), .A3(new_n773), .A4(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  NAND2_X1  g380(.A1(new_n518), .A2(G55), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n515), .A2(G93), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(new_n506), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G860), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n592), .A2(G559), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n546), .A2(new_n810), .ZN(new_n816));
  INV_X1    g391(.A(new_n810), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(new_n540), .C1(new_n544), .C2(new_n545), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n815), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT102), .Z(new_n822));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n820), .B2(KEYINPUT39), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n812), .B1(new_n822), .B2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n618), .B(new_n480), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G162), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n500), .A2(KEYINPUT72), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT4), .B1(new_n500), .B2(KEYINPUT72), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n504), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n497), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n768), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n726), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n778), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n705), .B(new_n609), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n482), .A2(G142), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n486), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n475), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n836), .B(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n827), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n835), .B2(new_n842), .ZN(new_n844));
  INV_X1    g419(.A(G37), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n835), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n827), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n835), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n844), .B(new_n845), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g427(.A(new_n819), .B(new_n602), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n592), .A2(G299), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n855));
  INV_X1    g430(.A(new_n592), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(new_n596), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n592), .A2(KEYINPUT104), .A3(G299), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n859), .A2(KEYINPUT41), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n863));
  INV_X1    g438(.A(new_n854), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT105), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n857), .A2(new_n858), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(KEYINPUT105), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n862), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n861), .B1(new_n869), .B2(new_n853), .ZN(new_n870));
  XOR2_X1   g445(.A(G303), .B(G288), .Z(new_n871));
  XNOR2_X1  g446(.A(G290), .B(new_n687), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT42), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n870), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G868), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(G868), .B2(new_n817), .ZN(G295));
  OAI21_X1  g454(.A(new_n878), .B1(G868), .B2(new_n817), .ZN(G331));
  INV_X1    g455(.A(new_n875), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT110), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(G301), .A2(KEYINPUT107), .ZN(new_n884));
  NAND2_X1  g459(.A1(G301), .A2(KEYINPUT107), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(G168), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(G168), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n816), .B(new_n818), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n819), .A2(new_n890), .A3(new_n886), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n891), .A3(KEYINPUT108), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n886), .ZN(new_n893));
  INV_X1    g468(.A(new_n819), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n868), .A2(new_n863), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n859), .A2(KEYINPUT41), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n889), .A2(new_n891), .A3(KEYINPUT109), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n894), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n859), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n883), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n906), .B(new_n882), .C1(new_n869), .C2(new_n897), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n907), .A3(new_n845), .ZN(new_n908));
  XOR2_X1   g483(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  INV_X1    g487(.A(new_n897), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n901), .A2(new_n863), .A3(new_n903), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n859), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n901), .A2(new_n903), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n916), .A2(new_n863), .A3(new_n868), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n881), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n906), .B(new_n875), .C1(new_n869), .C2(new_n897), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n918), .A2(new_n845), .A3(new_n919), .A4(new_n909), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n911), .A2(new_n912), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n845), .ZN(new_n922));
  INV_X1    g497(.A(new_n914), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n860), .B1(new_n923), .B2(new_n897), .ZN(new_n924));
  INV_X1    g499(.A(new_n917), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n875), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n905), .A2(new_n907), .A3(new_n845), .A4(new_n909), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n912), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n921), .A2(new_n929), .ZN(G397));
  XOR2_X1   g505(.A(new_n705), .B(new_n707), .Z(new_n931));
  INV_X1    g506(.A(G2067), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n768), .B(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G1996), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n726), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(G290), .A2(G1986), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G290), .A2(G1986), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT111), .B(G1384), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n830), .B2(new_n831), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(KEYINPUT45), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n472), .A2(new_n476), .A3(G40), .A4(new_n479), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G1384), .B1(new_n830), .B2(new_n831), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(G8), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(G305), .A2(KEYINPUT49), .ZN(new_n954));
  INV_X1    g529(.A(G1981), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n576), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G305), .A2(KEYINPUT49), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n954), .B2(new_n958), .ZN(new_n960));
  OR3_X1    g535(.A1(new_n952), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1976), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n961), .A2(new_n962), .A3(new_n679), .ZN(new_n963));
  NOR2_X1   g538(.A1(G305), .A2(G1981), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n953), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n946), .B1(new_n950), .B2(KEYINPUT45), .ZN(new_n966));
  INV_X1    g541(.A(new_n942), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n832), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT112), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n943), .A2(new_n970), .A3(KEYINPUT45), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n966), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n832), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(new_n946), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n972), .A2(G1971), .B1(G2090), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(G303), .A2(G8), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n979), .A2(KEYINPUT113), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT113), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n980), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(G8), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT114), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n978), .A2(new_n987), .A3(G8), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT52), .B1(G288), .B2(new_n962), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n953), .B(new_n990), .C1(new_n962), .C2(G288), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n952), .B1(G1976), .B2(new_n679), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n961), .B(new_n991), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n965), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n504), .ZN(new_n996));
  AND4_X1   g571(.A1(G138), .A2(new_n467), .A3(new_n475), .A4(new_n469), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n503), .B1(new_n997), .B2(new_n498), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n996), .B1(new_n998), .B2(new_n501), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n974), .B1(new_n999), .B2(new_n497), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n945), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n970), .B1(new_n943), .B2(KEYINPUT45), .ZN(new_n1003));
  NOR4_X1   g578(.A1(G164), .A2(KEYINPUT112), .A3(new_n1001), .A4(new_n942), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1002), .B(new_n443), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1005), .A2(new_n1006), .B1(new_n754), .B2(new_n977), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n950), .A2(KEYINPUT45), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1002), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(G301), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n975), .A2(new_n976), .A3(new_n946), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1001), .B1(G164), .B2(G1384), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1008), .A2(new_n946), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1011), .A2(new_n742), .B1(new_n1013), .B2(new_n750), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G286), .A2(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(KEYINPUT123), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1015), .B(new_n1018), .C1(new_n1014), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1018), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1013), .A2(new_n750), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n975), .A2(new_n976), .A3(new_n742), .A4(new_n946), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(G8), .B(new_n1021), .C1(new_n1024), .C2(G286), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1016), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT62), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1010), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g603(.A(KEYINPUT62), .B(new_n1016), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n984), .B1(new_n978), .B2(G8), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(KEYINPUT116), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n994), .B1(new_n1031), .B2(KEYINPUT116), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n989), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n995), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  NOR4_X1   g610(.A1(new_n944), .A2(new_n1006), .A3(G2078), .A4(new_n945), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1007), .A2(G301), .A3(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(G301), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1026), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT61), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT56), .B(G2072), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1002), .B(new_n1044), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1045));
  INV_X1    g620(.A(G1956), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n977), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G299), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n561), .A2(new_n565), .A3(new_n567), .A4(new_n1048), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1045), .A2(new_n1047), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n592), .B2(new_n1057), .ZN(new_n1058));
  NOR3_X1   g633(.A1(G164), .A2(G1384), .A3(new_n945), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n932), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1058), .B(new_n1060), .C1(new_n1011), .C2(G1348), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n592), .A2(new_n1057), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n951), .A2(G2067), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n794), .B2(new_n977), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1062), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1058), .A3(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n977), .A2(new_n794), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1056), .B1(new_n1068), .B2(new_n1064), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1045), .A2(new_n1047), .A3(new_n1052), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n972), .A2(new_n1044), .B1(new_n1046), .B2(new_n977), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1052), .A2(KEYINPUT119), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT61), .B(new_n1071), .C1(new_n1072), .C2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1055), .A2(new_n1070), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n972), .A2(new_n934), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT58), .B(G1341), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT120), .B1(new_n1059), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1081), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n951), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1080), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1079), .B1(new_n1088), .B2(new_n547), .ZN(new_n1089));
  AOI211_X1 g664(.A(KEYINPUT121), .B(new_n546), .C1(new_n1080), .C2(new_n1087), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT59), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n934), .B2(new_n972), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT121), .B1(new_n1092), .B2(new_n546), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(new_n1079), .A3(new_n547), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1078), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n592), .B1(new_n1068), .B2(new_n1064), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1053), .A2(new_n1098), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1034), .B(new_n1042), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1007), .A2(G301), .A3(new_n1009), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1101), .A2(KEYINPUT54), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n977), .A2(new_n754), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1037), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1105), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT124), .B1(new_n1105), .B2(G171), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1102), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1102), .B(KEYINPUT125), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1035), .B1(new_n1100), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1031), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1014), .A2(new_n1019), .A3(G286), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n994), .A2(new_n1116), .ZN(new_n1117));
  AND4_X1   g692(.A1(new_n989), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1034), .A2(KEYINPUT117), .A3(new_n1115), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n989), .A2(new_n1032), .A3(new_n1033), .A4(new_n1115), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT63), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1118), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n949), .B1(new_n1113), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n947), .B1(new_n933), .B2(new_n727), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT126), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n947), .A2(G1996), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT46), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT47), .Z(new_n1130));
  NOR2_X1   g705(.A1(new_n937), .A2(new_n947), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n947), .A2(new_n939), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(KEYINPUT48), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(KEYINPUT48), .B2(new_n1132), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n703), .A2(new_n707), .A3(new_n704), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n936), .A2(new_n1135), .B1(G2067), .B2(new_n768), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n948), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1130), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1124), .A2(new_n1138), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g714(.A1(new_n911), .A2(new_n920), .ZN(new_n1141));
  OAI21_X1  g715(.A(G319), .B1(new_n636), .B2(new_n637), .ZN(new_n1142));
  OR2_X1    g716(.A1(G227), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n1144));
  AND2_X1   g718(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1146));
  NOR3_X1   g720(.A1(new_n1145), .A2(new_n1146), .A3(G229), .ZN(new_n1147));
  NAND3_X1  g721(.A1(new_n1141), .A2(new_n851), .A3(new_n1147), .ZN(G225));
  INV_X1    g722(.A(G225), .ZN(G308));
endmodule


