//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  AND2_X1   g003(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209));
  XNOR2_X1  g008(.A(G197gat), .B(G204gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT22), .ZN(new_n211));
  INV_X1    g010(.A(G211gat), .ZN(new_n212));
  INV_X1    g011(.A(G218gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G211gat), .B(G218gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n209), .B1(new_n217), .B2(KEYINPUT29), .ZN(new_n218));
  XOR2_X1   g017(.A(G141gat), .B(G148gat), .Z(new_n219));
  INV_X1    g018(.A(G155gat), .ZN(new_n220));
  INV_X1    g019(.A(G162gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(KEYINPUT2), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n223), .B(new_n222), .C1(new_n227), .C2(KEYINPUT2), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n218), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n228), .A3(new_n209), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n217), .B1(new_n232), .B2(KEYINPUT29), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(G22gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(G228gat), .A2(G233gat), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n236), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n208), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n237), .A2(new_n238), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n239), .B1(new_n205), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G113gat), .ZN(new_n242));
  INV_X1    g041(.A(G120gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(G113gat), .B2(G120gat), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G127gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(G134gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(G127gat), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n244), .A2(new_n247), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n255), .A3(KEYINPUT72), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n262), .A2(KEYINPUT69), .A3(KEYINPUT24), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n269));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(KEYINPUT23), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR4_X1   g076(.A1(new_n268), .A2(new_n269), .A3(new_n272), .A4(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n271), .B2(KEYINPUT23), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n276), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  OAI22_X1  g083(.A1(new_n284), .A2(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  OAI211_X1 g084(.A(G183gat), .B(G190gat), .C1(new_n265), .C2(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n261), .A2(new_n284), .A3(KEYINPUT24), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n281), .B(new_n283), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n287), .ZN(new_n291));
  INV_X1    g090(.A(new_n285), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT66), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n269), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(KEYINPUT68), .B(new_n269), .C1(new_n290), .C2(new_n294), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n278), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n262), .B1(new_n302), .B2(KEYINPUT28), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(KEYINPUT28), .B2(new_n302), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n275), .A2(KEYINPUT70), .A3(KEYINPUT26), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n271), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n308), .A3(new_n270), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n310), .A2(new_n311), .B1(new_n307), .B2(new_n271), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(KEYINPUT71), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n304), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n260), .B1(new_n299), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n278), .ZN(new_n316));
  INV_X1    g115(.A(new_n298), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n293), .A2(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n288), .A2(new_n289), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n282), .A2(new_n272), .A3(new_n280), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT68), .B1(new_n321), .B2(new_n269), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n316), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n314), .ZN(new_n324));
  INV_X1    g123(.A(new_n260), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G227gat), .ZN(new_n327));
  INV_X1    g126(.A(G233gat), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n315), .B(new_n326), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT34), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n326), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n327), .A2(new_n328), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n332), .B(KEYINPUT64), .Z(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT34), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n330), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G15gat), .B(G43gat), .Z(new_n337));
  XNOR2_X1  g136(.A(G71gat), .B(G99gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n333), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n315), .B2(new_n326), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n341), .B2(KEYINPUT33), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT32), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  AOI221_X4 g144(.A(new_n343), .B1(KEYINPUT33), .B2(new_n339), .C1(new_n331), .C2(new_n333), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n336), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n299), .A2(new_n260), .A3(new_n314), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n325), .B1(new_n323), .B2(new_n324), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n333), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n353), .A3(new_n339), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n342), .A2(new_n344), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n331), .A2(new_n335), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(KEYINPUT34), .B2(new_n329), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n241), .A2(new_n347), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g161(.A(G226gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n328), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n299), .A2(new_n364), .A3(new_n314), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(KEYINPUT29), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(new_n323), .B2(new_n324), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n217), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n366), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n299), .B2(new_n314), .ZN(new_n370));
  INV_X1    g169(.A(new_n217), .ZN(new_n371));
  INV_X1    g170(.A(new_n364), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n323), .A2(new_n324), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n362), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n368), .A2(new_n374), .A3(new_n362), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379));
  XNOR2_X1  g178(.A(G57gat), .B(G85gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n229), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(new_n258), .A3(KEYINPUT4), .A4(new_n259), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n226), .A2(new_n228), .A3(new_n250), .A4(new_n255), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n229), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(new_n256), .A3(new_n231), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT74), .B1(new_n229), .B2(KEYINPUT3), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n386), .B(new_n391), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  AND4_X1   g194(.A1(new_n228), .A2(new_n226), .A3(new_n250), .A4(new_n255), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n226), .A2(new_n228), .B1(new_n250), .B2(new_n255), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(KEYINPUT75), .A3(new_n388), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT5), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n388), .B1(new_n396), .B2(new_n397), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n394), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n405), .A2(new_n392), .A3(new_n256), .A4(new_n231), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n389), .A2(new_n390), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n385), .A2(new_n258), .A3(new_n259), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(new_n390), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n406), .A2(new_n409), .A3(new_n400), .A4(new_n387), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n384), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT6), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n384), .A3(new_n410), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n416), .B2(new_n411), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n371), .B1(new_n370), .B2(new_n373), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(KEYINPUT73), .A3(KEYINPUT30), .A4(new_n362), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n368), .A2(KEYINPUT30), .A3(new_n374), .A4(new_n362), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT73), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n378), .A2(new_n417), .A3(new_n421), .A4(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT35), .B1(new_n359), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n237), .A2(new_n205), .A3(new_n238), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n240), .B2(new_n208), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(KEYINPUT35), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n347), .A2(KEYINPUT81), .A3(new_n358), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT81), .B1(new_n347), .B2(new_n358), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n433));
  INV_X1    g232(.A(new_n375), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n377), .A2(new_n376), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n421), .A2(new_n424), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT78), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n404), .A2(new_n410), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(new_n384), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n411), .A2(KEYINPUT78), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n415), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n412), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n433), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n424), .A2(new_n434), .A3(new_n435), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n445), .A2(KEYINPUT80), .A3(new_n421), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n426), .B1(new_n432), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n440), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n387), .B1(new_n406), .B2(new_n409), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n451), .B(KEYINPUT39), .C1(new_n388), .C2(new_n398), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT39), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n383), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT40), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT40), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n449), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n428), .B1(new_n436), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n420), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n362), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n368), .A2(new_n374), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(KEYINPUT37), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT38), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n362), .B1(new_n420), .B2(new_n461), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n418), .A2(KEYINPUT79), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n468), .B(KEYINPUT37), .C1(new_n464), .C2(KEYINPUT79), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n441), .A2(new_n412), .A3(new_n377), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n460), .A2(new_n473), .B1(new_n425), .B2(new_n428), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n347), .A2(KEYINPUT36), .A3(new_n358), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT36), .B1(new_n347), .B2(new_n358), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n448), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G64gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G57gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT87), .B(G57gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n479), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(G71gat), .B(G78gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(KEYINPUT88), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n482), .B(new_n485), .C1(KEYINPUT88), .C2(new_n484), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT9), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n479), .A2(G57gat), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n480), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n489), .A2(new_n484), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G231gat), .A2(G233gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(new_n251), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT16), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(G1gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G1gat), .B2(new_n497), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n500), .B(G8gat), .Z(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n486), .A2(new_n490), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(KEYINPUT21), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n496), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(new_n220), .ZN(new_n507));
  XNOR2_X1  g306(.A(G183gat), .B(G211gat), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n507), .B(new_n508), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n505), .A2(new_n510), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516));
  INV_X1    g315(.A(G85gat), .ZN(new_n517));
  INV_X1    g316(.A(G92gat), .ZN(new_n518));
  AOI22_X1  g317(.A1(KEYINPUT8), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G99gat), .B(G106gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G43gat), .B(G50gat), .Z(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT84), .B(KEYINPUT15), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT85), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT14), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT83), .B(G29gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(G36gat), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n527), .A2(new_n529), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n529), .A2(new_n537), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n525), .B(KEYINPUT85), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n529), .A2(new_n537), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT17), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n522), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n544), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n520), .B(new_n521), .Z(new_n548));
  INV_X1    g347(.A(KEYINPUT41), .ZN(new_n549));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT89), .Z(new_n551));
  OAI22_X1  g350(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n549), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(new_n253), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(new_n221), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n562), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n557), .A2(new_n558), .A3(new_n563), .A4(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n513), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT91), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n548), .A2(new_n491), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n503), .A2(new_n522), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT10), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n503), .A2(KEYINPUT10), .A3(new_n522), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n575), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n576), .B2(new_n577), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n573), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n581), .A2(new_n583), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT92), .B1(new_n585), .B2(new_n572), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n587));
  NOR4_X1   g386(.A1(new_n581), .A2(new_n587), .A3(new_n583), .A4(new_n573), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n569), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G197gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT11), .B(G169gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(KEYINPUT86), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n544), .A2(KEYINPUT17), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n598), .B(new_n501), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n502), .B1(new_n541), .B2(new_n545), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT86), .B1(new_n547), .B2(new_n501), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n501), .B(new_n544), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n605), .B(KEYINPUT13), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT18), .B1(new_n604), .B2(new_n605), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n597), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n604), .A2(new_n605), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT18), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n597), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n606), .A4(new_n610), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n591), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n478), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n417), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n436), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n627), .A2(G8gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT16), .B(G8gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT42), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(KEYINPUT42), .B2(new_n630), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT93), .ZN(G1325gat));
  INV_X1    g432(.A(KEYINPUT94), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n475), .B2(new_n476), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT36), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n345), .A2(new_n336), .A3(new_n346), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n357), .B1(new_n354), .B2(new_n355), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n347), .A2(KEYINPUT36), .A3(new_n358), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(KEYINPUT94), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(G15gat), .B1(new_n622), .B2(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n430), .A2(new_n431), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n644), .B1(new_n622), .B2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n622), .A2(new_n241), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT95), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  NAND2_X1  g451(.A1(new_n478), .A2(new_n568), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n513), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(new_n620), .A3(new_n589), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n536), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n624), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT45), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n474), .A2(new_n635), .A3(new_n641), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n448), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT97), .B(KEYINPUT44), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n568), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n567), .B1(new_n448), .B2(new_n662), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n664), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n667), .A2(new_n669), .B1(KEYINPUT44), .B2(new_n653), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n656), .B(KEYINPUT96), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n670), .A2(new_n417), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n661), .B1(new_n673), .B2(new_n659), .ZN(G1328gat));
  NAND2_X1  g473(.A1(new_n653), .A2(KEYINPUT44), .ZN(new_n675));
  AND4_X1   g474(.A1(KEYINPUT98), .A2(new_n663), .A3(new_n568), .A4(new_n664), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT98), .B1(new_n668), .B2(new_n664), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n436), .A3(new_n671), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n531), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n680), .B2(new_n679), .ZN(new_n682));
  INV_X1    g481(.A(new_n436), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n657), .A2(G36gat), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(G1329gat));
  NOR3_X1   g485(.A1(new_n657), .A2(G43gat), .A3(new_n646), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n678), .A2(new_n642), .A3(new_n671), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G43gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n690), .A2(KEYINPUT100), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n690), .A2(G43gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n688), .B1(new_n695), .B2(new_n687), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1330gat));
  NAND3_X1  g496(.A1(new_n678), .A2(new_n428), .A3(new_n671), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G50gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n241), .A2(G50gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT101), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n658), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(KEYINPUT102), .A2(KEYINPUT48), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n699), .A2(new_n705), .A3(new_n706), .A4(new_n702), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(G1331gat));
  AND4_X1   g509(.A1(new_n620), .A2(new_n663), .A3(new_n569), .A4(new_n589), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n624), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n481), .ZN(G1332gat));
  AND2_X1   g512(.A1(new_n711), .A2(new_n436), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  AND2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n714), .B2(new_n715), .ZN(G1333gat));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n642), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n646), .A2(G71gat), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n719), .A2(G71gat), .B1(new_n711), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g521(.A1(new_n711), .A2(new_n428), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g523(.A1(new_n513), .A2(new_n620), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT103), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n590), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n678), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G85gat), .B1(new_n728), .B2(new_n417), .ZN(new_n729));
  INV_X1    g528(.A(new_n726), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n668), .A2(KEYINPUT51), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT51), .B1(new_n668), .B2(new_n730), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n590), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n517), .A3(new_n624), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n735), .ZN(G1336gat));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n518), .A3(new_n436), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n728), .A2(new_n683), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n518), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT52), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n737), .B(new_n741), .C1(new_n738), .C2(new_n518), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n728), .B2(new_n643), .ZN(new_n744));
  INV_X1    g543(.A(G99gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n734), .A2(new_n745), .A3(new_n645), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(G1338gat));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n678), .A2(new_n428), .A3(new_n727), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G106gat), .ZN(new_n750));
  INV_X1    g549(.A(new_n733), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n241), .A2(G106gat), .A3(new_n590), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT104), .Z(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n748), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n731), .B2(new_n732), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n748), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n749), .B2(G106gat), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT105), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n757), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n750), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n749), .A2(G106gat), .B1(new_n751), .B2(new_n753), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n761), .B(new_n762), .C1(new_n748), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n759), .A2(new_n764), .ZN(G1339gat));
  OR2_X1    g564(.A1(new_n586), .A2(new_n588), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n579), .A2(new_n580), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n582), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n579), .A2(new_n580), .A3(new_n575), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(KEYINPUT54), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n572), .B1(new_n581), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT55), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(KEYINPUT55), .A3(new_n772), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n766), .A2(KEYINPUT106), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n586), .B2(new_n588), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n773), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n619), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n607), .A2(new_n609), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n604), .B2(new_n605), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n595), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n618), .A2(new_n589), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n568), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n776), .A2(new_n779), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n618), .A2(new_n565), .A3(new_n566), .A4(new_n783), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n513), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n569), .A2(new_n620), .A3(new_n590), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(new_n417), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n436), .A2(new_n428), .ZN(new_n795));
  AND4_X1   g594(.A1(new_n358), .A2(new_n794), .A3(new_n347), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT108), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(new_n242), .A3(new_n619), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n645), .A3(new_n795), .ZN(new_n799));
  OAI21_X1  g598(.A(G113gat), .B1(new_n799), .B2(new_n620), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1340gat));
  NAND3_X1  g600(.A1(new_n797), .A2(new_n243), .A3(new_n589), .ZN(new_n802));
  OAI21_X1  g601(.A(G120gat), .B1(new_n799), .B2(new_n590), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1341gat));
  NAND3_X1  g603(.A1(new_n796), .A2(new_n251), .A3(new_n655), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n799), .A2(new_n513), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n251), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT109), .ZN(G1342gat));
  NAND3_X1  g607(.A1(new_n796), .A2(new_n253), .A3(new_n568), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n811));
  OAI21_X1  g610(.A(G134gat), .B1(new_n799), .B2(new_n567), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(G1343gat));
  INV_X1    g612(.A(G141gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n789), .A2(new_n791), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT107), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n816), .A2(new_n817), .A3(new_n428), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n436), .A2(new_n417), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n643), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n770), .A2(new_n772), .ZN(new_n822));
  XNOR2_X1  g621(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n778), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n619), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n784), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n618), .A2(KEYINPUT110), .A3(new_n589), .A4(new_n783), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n567), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT112), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n567), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n788), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT113), .A3(new_n513), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n791), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n655), .B1(new_n831), .B2(new_n834), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(KEYINPUT113), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n428), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n821), .B1(new_n840), .B2(KEYINPUT57), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n814), .B1(new_n841), .B2(new_n619), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n642), .A2(new_n241), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n436), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n794), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(G141gat), .A3(new_n620), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT58), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n821), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n838), .A2(KEYINPUT113), .ZN(new_n850));
  INV_X1    g649(.A(new_n791), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n851), .B1(new_n838), .B2(KEYINPUT113), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n241), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n849), .B1(new_n853), .B2(new_n817), .ZN(new_n854));
  OAI21_X1  g653(.A(G141gat), .B1(new_n854), .B2(new_n620), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  INV_X1    g655(.A(new_n847), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n848), .A2(new_n858), .ZN(G1344gat));
  INV_X1    g658(.A(new_n846), .ZN(new_n860));
  INV_X1    g659(.A(G148gat), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n589), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n792), .A2(new_n793), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(KEYINPUT114), .A3(KEYINPUT57), .A4(new_n428), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n816), .A2(KEYINPUT57), .A3(new_n428), .A4(new_n818), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n766), .A2(new_n775), .A3(new_n774), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n832), .B1(new_n870), .B2(new_n787), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n513), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n241), .B1(new_n872), .B2(new_n791), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT115), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n851), .B1(new_n871), .B2(new_n513), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n875), .B(new_n817), .C1(new_n876), .C2(new_n241), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n869), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n879), .A2(new_n589), .A3(new_n643), .A4(new_n820), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n863), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT59), .B(new_n861), .C1(new_n841), .C2(new_n589), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n862), .B1(new_n881), .B2(new_n882), .ZN(G1345gat));
  AOI21_X1  g682(.A(G155gat), .B1(new_n860), .B2(new_n655), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n513), .A2(new_n220), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT116), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n841), .B2(new_n886), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n854), .B2(new_n567), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n860), .A2(new_n221), .A3(new_n568), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n359), .A2(new_n683), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n864), .A2(new_n417), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n619), .A2(new_n273), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT117), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n683), .A2(new_n624), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n645), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT118), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n864), .A2(new_n241), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n620), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n895), .A2(KEYINPUT119), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1348gat));
  OAI21_X1  g704(.A(new_n274), .B1(new_n892), .B2(new_n590), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT120), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n899), .A2(new_n274), .A3(new_n590), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n655), .A2(new_n300), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n892), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT121), .ZN(new_n912));
  OAI21_X1  g711(.A(G183gat), .B1(new_n899), .B2(new_n513), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT60), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n899), .B2(new_n567), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n568), .A2(new_n301), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n923), .A2(new_n924), .B1(new_n892), .B2(new_n925), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n844), .A2(new_n683), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n864), .A2(new_n417), .A3(new_n927), .ZN(new_n928));
  XOR2_X1   g727(.A(KEYINPUT123), .B(G197gat), .Z(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n619), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n643), .A2(new_n896), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n869), .B2(new_n878), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n933), .A3(new_n619), .ZN(new_n934));
  INV_X1    g733(.A(new_n929), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n932), .B2(new_n619), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n930), .B1(new_n936), .B2(new_n937), .ZN(G1352gat));
  INV_X1    g737(.A(G204gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n928), .A2(new_n939), .A3(new_n589), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n941), .A2(KEYINPUT125), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(new_n945));
  AOI211_X1 g744(.A(new_n590), .B(new_n931), .C1(new_n869), .C2(new_n878), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n939), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n212), .A3(new_n655), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n949), .B(new_n212), .C1(new_n932), .C2(new_n655), .ZN(new_n950));
  INV_X1    g749(.A(new_n931), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n879), .A2(new_n655), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n948), .B1(new_n950), .B2(new_n953), .ZN(G1354gat));
  AOI21_X1  g753(.A(G218gat), .B1(new_n928), .B2(new_n568), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT126), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n957));
  AOI211_X1 g756(.A(new_n213), .B(new_n567), .C1(new_n932), .C2(new_n957), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n932), .A2(new_n957), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1355gat));
endmodule


