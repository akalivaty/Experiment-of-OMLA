//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G131), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G214), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT86), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(G237), .A2(G953), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n198), .B(G214), .C1(KEYINPUT86), .C2(G143), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n191), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT17), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n191), .A3(new_n199), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT16), .ZN(new_n209));
  OR3_X1    g023(.A1(new_n207), .A2(KEYINPUT16), .A3(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G146), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n209), .B2(new_n210), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n200), .A2(KEYINPUT17), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n197), .A2(new_n199), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT18), .A2(G131), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n206), .A2(new_n208), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n217), .A2(new_n218), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n197), .A2(new_n199), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT87), .ZN(new_n226));
  INV_X1    g040(.A(new_n218), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n226), .B1(new_n225), .B2(new_n227), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n224), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n190), .B1(new_n232), .B2(KEYINPUT93), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT93), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n216), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(KEYINPUT94), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n216), .A2(new_n231), .A3(new_n190), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT94), .B1(new_n233), .B2(new_n235), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n187), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G475), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT90), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n197), .A2(new_n191), .A3(new_n199), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n211), .B1(new_n243), .B2(new_n200), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT19), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n206), .B(new_n208), .C1(KEYINPUT88), .C2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n219), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n245), .B1(new_n249), .B2(G146), .ZN(new_n250));
  INV_X1    g064(.A(new_n248), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n222), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n252), .A2(KEYINPUT89), .A3(new_n220), .A4(new_n247), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n244), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n223), .A2(new_n221), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n225), .B2(new_n227), .ZN(new_n256));
  INV_X1    g070(.A(new_n230), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(new_n228), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n242), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n260));
  INV_X1    g074(.A(new_n190), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n250), .A2(new_n253), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n212), .B1(new_n201), .B2(new_n203), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT90), .A3(new_n231), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n260), .A3(new_n261), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n237), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n257), .A2(new_n228), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n268), .A2(new_n224), .B1(new_n262), .B2(new_n263), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n190), .B1(new_n269), .B2(KEYINPUT90), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n260), .B1(new_n270), .B2(new_n259), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT92), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT20), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n265), .A2(new_n261), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT90), .B1(new_n264), .B2(new_n231), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT91), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(new_n237), .A3(new_n266), .ZN(new_n277));
  NOR2_X1   g091(.A1(G475), .A2(G902), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n272), .A2(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT92), .ZN(new_n280));
  AND4_X1   g094(.A1(new_n280), .A2(new_n277), .A3(new_n273), .A4(new_n278), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n241), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n284), .A2(G122), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(G122), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G107), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT13), .ZN(new_n290));
  INV_X1    g104(.A(G128), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(G143), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(G143), .ZN(new_n293));
  OR3_X1    g107(.A1(new_n292), .A2(KEYINPUT95), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  INV_X1    g109(.A(new_n293), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT95), .B1(new_n296), .B2(new_n290), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n294), .B(G134), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT68), .B(G134), .ZN(new_n299));
  XNOR2_X1  g113(.A(G128), .B(G143), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n289), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n287), .A2(new_n288), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n299), .B(new_n300), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n285), .B1(new_n286), .B2(KEYINPUT14), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n306), .A2(KEYINPUT96), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(KEYINPUT96), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n303), .B(new_n304), .C1(new_n309), .C2(new_n288), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(new_n312), .A3(G953), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n302), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n302), .B2(new_n310), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT97), .B1(new_n316), .B2(G902), .ZN(new_n317));
  INV_X1    g131(.A(G478), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT15), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT97), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n320), .B(new_n187), .C1(new_n314), .C2(new_n315), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n316), .A2(G902), .A3(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n283), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G110), .B(G122), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G116), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n284), .A2(G119), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT5), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n336));
  INV_X1    g150(.A(G113), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT2), .B(G113), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n334), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n338), .A3(KEYINPUT85), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n288), .A3(G104), .ZN(new_n349));
  INV_X1    g163(.A(G101), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n189), .A2(G107), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n347), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n288), .A2(G104), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n189), .A2(G107), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT80), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(KEYINPUT81), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n352), .A2(new_n355), .A3(new_n358), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n358), .B1(new_n352), .B2(new_n355), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n346), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n344), .A2(KEYINPUT71), .ZN(new_n366));
  INV_X1    g180(.A(new_n334), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n342), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G101), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n342), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT71), .A3(new_n344), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(new_n374), .A3(G101), .ZN(new_n375));
  AND4_X1   g189(.A1(new_n368), .A2(new_n371), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n330), .B1(new_n365), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n346), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n364), .A2(new_n360), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n366), .B(new_n372), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n371), .A3(new_n375), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n382), .A3(new_n329), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n383), .A3(KEYINPUT6), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT65), .B1(new_n220), .B2(G143), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT65), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n196), .A3(G146), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n220), .A2(KEYINPUT64), .A3(G143), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT64), .B1(new_n220), .B2(G143), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n385), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(KEYINPUT0), .A2(G128), .ZN(new_n391));
  NOR2_X1   g205(.A1(KEYINPUT0), .A2(G128), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n220), .A2(G143), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT66), .B1(new_n196), .B2(G146), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT66), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n220), .A3(G143), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n390), .A2(new_n393), .B1(new_n398), .B2(new_n391), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(new_n207), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n220), .A2(G143), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n291), .B1(new_n401), .B2(KEYINPUT1), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n385), .A2(new_n387), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n220), .A2(KEYINPUT64), .A3(G143), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n402), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n398), .A2(new_n410), .A3(G128), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n207), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n400), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G224), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G953), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(new_n330), .C1(new_n365), .C2(new_n376), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n384), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n329), .B(KEYINPUT8), .Z(new_n420));
  NAND2_X1  g234(.A1(new_n346), .A2(new_n356), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n357), .A2(new_n359), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n344), .A3(new_n339), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n420), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT7), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n415), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n400), .A2(new_n412), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n400), .B2(new_n412), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n429), .B2(new_n383), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n419), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G210), .B1(G237), .B2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n419), .A2(new_n430), .A3(new_n432), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n328), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n193), .A2(G952), .ZN(new_n437));
  INV_X1    g251(.A(G234), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(new_n192), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n187), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(G898), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n436), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n326), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n312), .B1(G234), .B2(new_n187), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT75), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT22), .B(G137), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n331), .A2(G128), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n291), .A2(KEYINPUT23), .A3(G119), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n331), .A2(G128), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(KEYINPUT23), .ZN(new_n456));
  XNOR2_X1  g270(.A(G119), .B(G128), .ZN(new_n457));
  INV_X1    g271(.A(G110), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT24), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT24), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G110), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n456), .A2(G110), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n212), .B2(new_n213), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT74), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n463), .B(KEYINPUT74), .C1(new_n212), .C2(new_n213), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n291), .A2(G119), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n459), .B(new_n461), .C1(new_n469), .C2(new_n455), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n456), .B2(G110), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n471), .A2(new_n211), .A3(new_n221), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT76), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT76), .ZN(new_n475));
  AOI211_X1 g289(.A(new_n475), .B(new_n472), .C1(new_n466), .C2(new_n467), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n452), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n472), .B1(new_n466), .B2(new_n467), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n452), .B1(new_n478), .B2(KEYINPUT76), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n187), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n477), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n480), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n448), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n467), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n209), .A2(new_n210), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n220), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n211), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT74), .B1(new_n489), .B2(new_n463), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n473), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n475), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n478), .A2(KEYINPUT76), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n479), .B1(new_n494), .B2(new_n452), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n447), .A2(G902), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n485), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT11), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT67), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT11), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G137), .ZN(new_n504));
  INV_X1    g318(.A(G134), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G134), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n503), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(KEYINPUT11), .A3(G134), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n509), .B2(new_n504), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT69), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT67), .B(KEYINPUT11), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n299), .B2(G137), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n299), .A2(G137), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n516), .A2(new_n191), .A3(new_n517), .A4(new_n511), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT69), .B(G131), .C1(new_n510), .C2(new_n512), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n399), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n368), .A2(new_n373), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n409), .A2(new_n411), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n299), .A2(G137), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n504), .A2(G134), .ZN(new_n525));
  OAI21_X1  g339(.A(G131), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n518), .A3(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n521), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT28), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n198), .A2(G210), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT27), .Z(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(G101), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  NAND3_X1  g348(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT28), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n530), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n521), .A2(KEYINPUT30), .A3(new_n527), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n521), .A2(new_n527), .A3(KEYINPUT72), .A4(KEYINPUT30), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n521), .A2(new_n527), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n545), .B(new_n381), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n534), .B1(new_n552), .B2(new_n535), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n538), .A2(new_n539), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n187), .B(new_n540), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n534), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n528), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT73), .B(KEYINPUT31), .Z(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n534), .B1(new_n530), .B2(new_n537), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n557), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n546), .A2(new_n548), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT70), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n564), .A2(new_n549), .B1(new_n543), .B2(new_n544), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n565), .B2(new_n381), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT31), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n559), .B(new_n561), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(G472), .A2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT32), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n555), .A2(G472), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n569), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n571), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n498), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G469), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n187), .ZN(new_n580));
  INV_X1    g394(.A(new_n402), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n395), .A2(new_n397), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n394), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n356), .B1(new_n583), .B2(new_n411), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT79), .B1(new_n584), .B2(KEYINPUT10), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT79), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n398), .A2(new_n402), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n410), .A2(G128), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n589), .B(new_n394), .C1(new_n395), .C2(new_n397), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n586), .B(new_n587), .C1(new_n591), .C2(new_n356), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n390), .A2(new_n393), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n398), .A2(new_n391), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n375), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n369), .A2(G101), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT78), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT78), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n399), .A2(new_n371), .A3(new_n600), .A4(new_n375), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n585), .A2(new_n592), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n519), .A2(new_n520), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT10), .B1(new_n408), .B2(new_n590), .ZN(new_n604));
  AOI211_X1 g418(.A(KEYINPUT82), .B(new_n604), .C1(new_n360), .C2(new_n364), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT82), .ZN(new_n606));
  INV_X1    g420(.A(new_n604), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n379), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n602), .B(new_n603), .C1(new_n605), .C2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT83), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n362), .A2(new_n363), .A3(new_n361), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT81), .B1(new_n357), .B2(new_n359), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n607), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT82), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n379), .A2(new_n606), .A3(new_n607), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n617), .A2(KEYINPUT83), .A3(new_n603), .A4(new_n602), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n603), .ZN(new_n620));
  OAI22_X1  g434(.A1(new_n523), .A2(new_n422), .B1(new_n356), .B2(new_n591), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  NAND2_X1  g437(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(G110), .B(G140), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n193), .A2(G227), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n625), .B(new_n626), .Z(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT77), .Z(new_n628));
  OAI21_X1  g442(.A(new_n602), .B1(new_n605), .B2(new_n608), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n620), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT84), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT84), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(new_n632), .A3(new_n620), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n627), .B1(new_n611), .B2(new_n618), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n624), .A2(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n580), .B1(new_n636), .B2(G469), .ZN(new_n637));
  INV_X1    g451(.A(new_n627), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n634), .B2(new_n619), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n619), .A2(new_n638), .A3(new_n623), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n579), .B(new_n187), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n578), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n446), .A2(new_n576), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G101), .ZN(G3));
  INV_X1    g458(.A(G472), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n568), .B2(new_n187), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n552), .A2(new_n557), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n560), .B1(new_n647), .B2(KEYINPUT31), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n570), .B1(new_n648), .B2(new_n559), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n646), .A2(new_n649), .A3(new_n498), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n642), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(KEYINPUT98), .Z(new_n652));
  NAND3_X1  g466(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n316), .B(KEYINPUT33), .Z(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n187), .A2(G478), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n282), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n445), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G104), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT99), .B(KEYINPUT34), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  AOI21_X1  g477(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n277), .A2(new_n273), .A3(new_n278), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n665), .A2(new_n666), .B1(G475), .B2(new_n240), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(KEYINPUT100), .A3(new_n444), .A4(new_n324), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  INV_X1    g483(.A(new_n666), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n241), .B(new_n324), .C1(new_n670), .C2(new_n664), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n669), .B1(new_n671), .B2(new_n443), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n668), .A2(new_n672), .A3(new_n436), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n652), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT101), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT35), .B(G107), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  AOI21_X1  g491(.A(KEYINPUT25), .B1(new_n495), .B2(new_n187), .ZN(new_n678));
  INV_X1    g492(.A(new_n484), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n447), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n491), .B(KEYINPUT102), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT36), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n452), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n496), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n680), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n496), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n684), .B2(new_n685), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT103), .B1(new_n485), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n646), .A3(new_n649), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n446), .A2(new_n694), .A3(new_n642), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT37), .B(G110), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G12));
  NAND2_X1  g511(.A1(new_n568), .A2(new_n572), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n552), .A2(new_n535), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n554), .B1(new_n699), .B2(new_n556), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n187), .B1(new_n538), .B2(new_n539), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n698), .B(new_n702), .C1(new_n649), .C2(KEYINPUT32), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n441), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n439), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n671), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n689), .A2(new_n692), .A3(new_n436), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n642), .A2(new_n703), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G128), .ZN(G30));
  XNOR2_X1  g525(.A(new_n706), .B(KEYINPUT39), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n642), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT40), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT40), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n556), .B1(new_n528), .B2(new_n529), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT104), .ZN(new_n717));
  AOI21_X1  g531(.A(G902), .B1(new_n647), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n575), .B(new_n698), .C1(new_n645), .C2(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n434), .A2(new_n435), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT38), .Z(new_n721));
  NAND2_X1  g535(.A1(new_n282), .A2(new_n324), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n680), .A2(new_n687), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n328), .A3(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n714), .A2(new_n715), .A3(new_n719), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  AND3_X1   g541(.A1(new_n282), .A2(new_n657), .A3(new_n706), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n642), .A2(new_n703), .A3(new_n709), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT105), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n689), .A2(new_n692), .A3(new_n436), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n575), .B2(new_n573), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n642), .A4(new_n728), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT106), .B(G146), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G48));
  OAI21_X1  g551(.A(new_n187), .B1(new_n639), .B2(new_n640), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G469), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n577), .A3(new_n641), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n576), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n659), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n673), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR2_X1   g562(.A1(new_n326), .A2(new_n443), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n732), .A2(new_n740), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  XOR2_X1   g565(.A(new_n569), .B(KEYINPUT107), .Z(new_n752));
  NAND2_X1  g566(.A1(new_n568), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(new_n498), .A3(new_n646), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n722), .A2(new_n445), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n740), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  NAND4_X1  g572(.A1(new_n739), .A2(new_n577), .A3(new_n641), .A4(new_n436), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(G902), .B1(new_n648), .B2(new_n559), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n723), .B(new_n753), .C1(new_n761), .C2(new_n645), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n282), .A2(new_n657), .A3(new_n706), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  NOR2_X1   g580(.A1(new_n578), .A2(new_n328), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n720), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n580), .B(KEYINPUT108), .Z(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n636), .B2(G469), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n768), .B1(new_n771), .B2(new_n641), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n576), .A2(new_n772), .A3(new_n728), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT109), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n576), .A2(new_n772), .A3(new_n777), .A4(new_n728), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n773), .A2(new_n776), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT42), .B1(new_n773), .B2(KEYINPUT109), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n775), .B1(new_n782), .B2(new_n778), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G131), .ZN(G33));
  NAND3_X1  g600(.A1(new_n576), .A2(new_n772), .A3(new_n708), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  OAI21_X1  g602(.A(G469), .B1(new_n636), .B2(KEYINPUT45), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(KEYINPUT45), .B2(new_n636), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(new_n770), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n790), .A2(new_n792), .A3(new_n770), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n641), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(new_n577), .A3(new_n712), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n720), .A2(new_n327), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT112), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n283), .A2(new_n657), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT43), .B1(new_n800), .B2(KEYINPUT111), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n723), .ZN(new_n804));
  INV_X1    g618(.A(new_n646), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n804), .B1(new_n805), .B2(new_n574), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT44), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n803), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n799), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n796), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  NOR4_X1   g627(.A1(new_n703), .A2(new_n763), .A3(new_n497), .A4(new_n797), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n795), .A2(KEYINPUT47), .A3(new_n577), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT47), .B1(new_n795), .B2(new_n577), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(KEYINPUT113), .B(G140), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(G42));
  AND2_X1   g634(.A1(new_n739), .A2(new_n641), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT49), .Z(new_n822));
  NAND4_X1  g636(.A1(new_n283), .A2(new_n497), .A3(new_n657), .A4(new_n767), .ZN(new_n823));
  OR4_X1    g637(.A1(new_n719), .A2(new_n822), .A3(new_n721), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n825));
  INV_X1    g639(.A(new_n762), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n772), .A3(new_n728), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n787), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n667), .A2(new_n325), .A3(new_n706), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n693), .A3(new_n797), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n703), .A3(new_n642), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(KEYINPUT114), .A3(new_n703), .A4(new_n642), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n828), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n740), .B(new_n576), .C1(new_n673), .C2(new_n659), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n446), .B(new_n642), .C1(new_n576), .C2(new_n694), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n283), .A2(new_n324), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n445), .B1(new_n840), .B2(new_n658), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n642), .A3(new_n650), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n750), .A3(new_n757), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n835), .A2(new_n839), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n784), .B2(new_n781), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n642), .A2(new_n703), .A3(new_n709), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n847), .A2(new_n708), .B1(new_n760), .B2(new_n764), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n723), .A2(new_n578), .A3(new_n707), .ZN(new_n849));
  INV_X1    g663(.A(new_n771), .ZN(new_n850));
  INV_X1    g664(.A(new_n641), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(KEYINPUT115), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n722), .A2(new_n328), .A3(new_n720), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n719), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(KEYINPUT52), .A2(new_n735), .A3(new_n848), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n735), .A2(new_n848), .A3(new_n857), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(KEYINPUT116), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n859), .A2(new_n863), .A3(new_n860), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n846), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n728), .A2(new_n805), .A3(new_n723), .A4(new_n753), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n710), .B1(new_n759), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n734), .B2(new_n730), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(KEYINPUT52), .A3(new_n857), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n861), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n846), .A2(KEYINPUT53), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n825), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n846), .B(KEYINPUT53), .C1(new_n862), .C2(new_n864), .ZN(new_n875));
  INV_X1    g689(.A(new_n872), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n838), .A2(new_n843), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n779), .A2(new_n780), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n877), .B(new_n835), .C1(new_n878), .C2(new_n783), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n866), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n875), .A2(new_n880), .A3(new_n825), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n740), .A2(new_n755), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n721), .A2(new_n327), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n803), .A2(new_n882), .A3(new_n440), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n821), .A2(new_n440), .A3(new_n720), .A4(new_n767), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n888), .A2(new_n801), .A3(new_n802), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n719), .A3(new_n498), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n282), .A2(new_n657), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n889), .A2(new_n826), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n884), .A2(new_n886), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n817), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n821), .A2(new_n578), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n815), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n803), .A2(new_n440), .A3(new_n755), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n799), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n896), .A2(new_n897), .ZN(new_n905));
  AND4_X1   g719(.A1(KEYINPUT51), .A2(new_n898), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n890), .A2(new_n282), .A3(new_n657), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n907), .B(new_n437), .C1(new_n759), .C2(new_n902), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n889), .A2(new_n576), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n909), .A2(KEYINPUT48), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(KEYINPUT48), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n896), .B1(new_n901), .B2(new_n903), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(KEYINPUT51), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n874), .A2(new_n881), .A3(new_n906), .A4(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(G952), .A2(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n824), .B1(new_n915), .B2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n193), .A2(G952), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n384), .A2(new_n418), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n416), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n187), .B1(new_n875), .B2(new_n880), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(G210), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(KEYINPUT119), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n921), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n921), .A2(KEYINPUT120), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n923), .B(new_n926), .C1(KEYINPUT119), .C2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n918), .B1(new_n928), .B2(new_n930), .ZN(G51));
  AOI21_X1  g745(.A(new_n825), .B1(new_n875), .B2(new_n880), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n881), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n769), .B(KEYINPUT57), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n933), .A2(new_n934), .B1(new_n639), .B2(new_n640), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n922), .A2(new_n790), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n918), .B1(new_n935), .B2(new_n936), .ZN(G54));
  AND2_X1   g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n922), .A2(new_n277), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n277), .B1(new_n922), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n918), .ZN(G60));
  INV_X1    g755(.A(new_n918), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n654), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n942), .B1(new_n933), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT52), .B1(new_n870), .B2(new_n857), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n871), .B1(new_n949), .B2(new_n863), .ZN(new_n950));
  INV_X1    g764(.A(new_n864), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n879), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n873), .B1(new_n952), .B2(KEYINPUT53), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n875), .A2(new_n880), .A3(new_n825), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n944), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n948), .B1(new_n956), .B2(new_n654), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n945), .B1(new_n874), .B2(new_n881), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(KEYINPUT121), .A3(new_n655), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n947), .B1(new_n957), .B2(new_n959), .ZN(G63));
  NAND2_X1  g774(.A1(new_n875), .A2(new_n880), .ZN(new_n961));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT122), .Z(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n495), .B(KEYINPUT123), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n918), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  INV_X1    g782(.A(new_n964), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n875), .B2(new_n880), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n686), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n967), .A2(KEYINPUT124), .A3(new_n968), .A4(new_n971), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n974));
  INV_X1    g788(.A(new_n966), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n942), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n961), .A2(new_n686), .A3(new_n964), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n973), .B(new_n974), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n972), .A2(new_n978), .ZN(G66));
  OAI21_X1  g793(.A(G953), .B1(new_n442), .B2(new_n414), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n877), .B2(G953), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n919), .B1(G898), .B2(new_n193), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G69));
  XOR2_X1   g797(.A(new_n565), .B(new_n249), .Z(new_n984));
  NAND2_X1  g798(.A1(G900), .A2(G953), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n576), .A2(new_n856), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n796), .B1(new_n811), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n870), .A2(new_n787), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n818), .A2(new_n987), .A3(new_n785), .A4(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n984), .B(new_n985), .C1(new_n989), .C2(G953), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n840), .A2(new_n658), .ZN(new_n991));
  OR4_X1    g805(.A1(new_n742), .A2(new_n991), .A3(new_n713), .A4(new_n797), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n818), .A2(new_n812), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n870), .A2(new_n726), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT62), .Z(new_n995));
  AOI21_X1  g809(.A(G953), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n990), .B1(new_n996), .B2(new_n984), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n990), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n997), .B(new_n1000), .Z(G72));
  NAND3_X1  g815(.A1(new_n993), .A2(new_n877), .A3(new_n995), .ZN(new_n1002));
  XNOR2_X1  g816(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n645), .A2(new_n187), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1003), .B(new_n1004), .Z(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n556), .B1(new_n552), .B2(new_n535), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n699), .A2(new_n534), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1005), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1009), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n953), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n877), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1005), .B1(new_n989), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1009), .B(KEYINPUT127), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AND4_X1   g830(.A1(new_n942), .A2(new_n1008), .A3(new_n1012), .A4(new_n1016), .ZN(G57));
endmodule


