//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n462), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT68), .B1(new_n470), .B2(G125), .ZN(new_n471));
  OAI211_X1 g046(.A(KEYINPUT68), .B(G125), .C1(new_n463), .C2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n468), .B1(new_n474), .B2(G2105), .ZN(G160));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n464), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(new_n462), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(new_n470), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n462), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  OAI22_X1  g063(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(new_n462), .A3(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n476), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT69), .B1(new_n470), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n489), .B1(new_n497), .B2(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n506), .A2(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n504), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  AOI22_X1  g091(.A1(new_n505), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n509), .A2(new_n508), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n506), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT70), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(G51), .A2(new_n530), .B1(new_n521), .B2(new_n522), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n531), .B(new_n532), .C1(new_n518), .C2(new_n517), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n526), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n503), .ZN(new_n536));
  INV_X1    g111(.A(new_n512), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT71), .B(G90), .Z(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n537), .A2(new_n539), .B1(G52), .B2(new_n530), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n536), .A2(new_n540), .A3(KEYINPUT72), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n535), .A2(new_n503), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n506), .A2(new_n544), .B1(new_n512), .B2(new_n538), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n542), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n541), .A2(new_n546), .ZN(G171));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n506), .A2(new_n548), .B1(new_n512), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n501), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n503), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n506), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n530), .A2(new_n562), .A3(G53), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n501), .A2(G65), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT73), .Z(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n537), .A2(G91), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT72), .B1(new_n536), .B2(new_n540), .ZN(new_n572));
  NOR3_X1   g147(.A1(new_n543), .A2(new_n545), .A3(new_n542), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n541), .A2(new_n546), .A3(KEYINPUT74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  OAI21_X1  g153(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n501), .A2(new_n505), .A3(G87), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT75), .B1(new_n512), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n501), .A2(new_n505), .A3(new_n585), .A4(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n518), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G48), .B2(new_n530), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n530), .A2(G47), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT76), .B(G85), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n593), .B1(new_n512), .B2(new_n594), .C1(new_n595), .C2(new_n503), .ZN(G290));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n512), .A2(KEYINPUT77), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT77), .B1(new_n512), .B2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n598), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT78), .B(G66), .Z(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n518), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n576), .B2(G868), .ZN(G284));
  AOI21_X1  g185(.A(new_n609), .B1(new_n576), .B2(G868), .ZN(G321));
  NOR2_X1   g186(.A1(G299), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g188(.A(new_n612), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g189(.A(G860), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n608), .B1(G559), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT79), .Z(G148));
  OR2_X1    g192(.A1(new_n608), .A2(G559), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n470), .A2(new_n466), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n477), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n479), .A2(G123), .ZN(new_n630));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G2096), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n627), .A2(new_n628), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT17), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  OR3_X1    g235(.A1(new_n657), .A2(new_n655), .A3(new_n658), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n655), .A3(new_n658), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT18), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n634), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT83), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n670), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n670), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT86), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n684), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G32), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n477), .A2(G141), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT95), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n479), .A2(G129), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT26), .Z(new_n696));
  AOI21_X1  g271(.A(KEYINPUT96), .B1(new_n466), .B2(G105), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n466), .A2(KEYINPUT96), .A3(G105), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n694), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n691), .B1(new_n700), .B2(new_n690), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT97), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT27), .B(G1996), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G27), .A2(G29), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G164), .B2(G29), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT100), .B(G2078), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT24), .ZN(new_n709));
  INV_X1    g284(.A(G34), .ZN(new_n710));
  AOI21_X1  g285(.A(G29), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G160), .B2(new_n690), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n708), .B1(G2084), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n690), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n690), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT29), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  OR2_X1    g293(.A1(G29), .A2(G33), .ZN(new_n719));
  NAND2_X1  g294(.A1(G115), .A2(G2104), .ZN(new_n720));
  INV_X1    g295(.A(G127), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n476), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n462), .B1(new_n722), .B2(KEYINPUT94), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(KEYINPUT94), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n725));
  NAND2_X1  g300(.A1(G103), .A2(G2104), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G2105), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n477), .A2(G139), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n719), .B1(new_n730), .B2(new_n690), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n717), .A2(G2090), .B1(new_n718), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n477), .A2(G140), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n479), .A2(G128), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n462), .A2(G116), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n690), .A2(G26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT28), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2067), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G19), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n554), .B2(new_n743), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1341), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n633), .A2(new_n690), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(KEYINPUT99), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT31), .B(G11), .Z(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT30), .B(G28), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n690), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n747), .B2(KEYINPUT99), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n742), .A2(new_n746), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n704), .A2(new_n714), .A3(new_n732), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n743), .A2(G20), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G168), .A2(new_n743), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n743), .B2(G21), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT98), .B(G1966), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n743), .A2(G5), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G171), .B2(new_n743), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n764), .B1(G1961), .B2(new_n766), .C1(G2084), .C2(new_n713), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n743), .A2(G4), .ZN(new_n768));
  AND3_X1   g343(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n743), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT93), .B(G1348), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n702), .B2(new_n703), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n731), .A2(new_n718), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G1961), .B2(new_n766), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(G2090), .B2(new_n717), .C1(new_n762), .C2(new_n763), .ZN(new_n776));
  NOR4_X1   g351(.A1(new_n754), .A2(new_n767), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n743), .A2(G23), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n780));
  NAND2_X1  g355(.A1(G288), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(KEYINPUT91), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n779), .B1(new_n783), .B2(new_n743), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n743), .A2(G22), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G166), .B2(new_n743), .ZN(new_n788));
  INV_X1    g363(.A(G1971), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n743), .A2(G6), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G305), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT32), .B(G1981), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n792), .A2(new_n794), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n786), .A2(new_n790), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT92), .Z(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT34), .Z(new_n799));
  MUX2_X1   g374(.A(G24), .B(G290), .S(G16), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT90), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G1986), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n690), .A2(G25), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n477), .A2(G131), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n479), .A2(G119), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n462), .A2(G107), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT87), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT88), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n803), .B1(new_n812), .B2(new_n690), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT89), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n802), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n799), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n799), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n778), .B1(new_n821), .B2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n777), .ZN(G150));
  NAND2_X1  g401(.A1(new_n769), .A2(G559), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT38), .Z(new_n828));
  XOR2_X1   g403(.A(KEYINPUT102), .B(G55), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n530), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n501), .A2(new_n505), .A3(G93), .ZN(new_n831));
  AND2_X1   g406(.A1(G80), .A2(G543), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n501), .B2(G67), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n830), .B(new_n831), .C1(new_n833), .C2(new_n503), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT103), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n518), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(G651), .B1(new_n837), .B2(new_n832), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n831), .A4(new_n830), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n530), .A2(G43), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n841), .B1(new_n549), .B2(new_n512), .C1(new_n842), .C2(new_n503), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n835), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n554), .B2(new_n834), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n835), .A2(new_n840), .A3(new_n845), .A4(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n828), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(new_n615), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n835), .A2(new_n840), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(G145));
  INV_X1    g432(.A(new_n633), .ZN(new_n858));
  XNOR2_X1  g433(.A(G164), .B(new_n737), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n693), .A2(new_n699), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n862), .A3(new_n730), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n730), .A2(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n700), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  INV_X1    g441(.A(G118), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(G2105), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n479), .B2(G130), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n477), .A2(G142), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n870), .A2(KEYINPUT106), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(KEYINPUT106), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n863), .A2(new_n865), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n873), .B1(new_n863), .B2(new_n865), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n860), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n859), .A3(new_n874), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n809), .B(new_n624), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n880), .B1(new_n877), .B2(new_n879), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n858), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n877), .A2(new_n879), .ZN(new_n886));
  INV_X1    g461(.A(new_n880), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n888), .A2(new_n882), .A3(new_n633), .A4(new_n881), .ZN(new_n889));
  XNOR2_X1  g464(.A(G160), .B(G162), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n890), .B1(new_n885), .B2(new_n889), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(G395));
  INV_X1    g472(.A(G868), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n854), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n618), .B(new_n849), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n769), .A2(new_n901), .A3(G299), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n602), .A2(G299), .A3(new_n603), .A4(new_n607), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT108), .ZN(new_n904));
  INV_X1    g479(.A(G299), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n608), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n906), .A2(new_n909), .A3(new_n903), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n907), .B2(KEYINPUT41), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n908), .B1(new_n912), .B2(new_n900), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n913), .B(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n783), .B(G305), .ZN(new_n917));
  XOR2_X1   g492(.A(G303), .B(G290), .Z(new_n918));
  XOR2_X1   g493(.A(new_n917), .B(new_n918), .Z(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n914), .B2(KEYINPUT42), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n916), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n899), .B1(new_n922), .B2(new_n898), .ZN(G295));
  OAI21_X1  g498(.A(new_n899), .B1(new_n922), .B2(new_n898), .ZN(G331));
  NAND3_X1  g499(.A1(new_n574), .A2(G168), .A3(new_n575), .ZN(new_n925));
  NAND2_X1  g500(.A1(G286), .A2(G171), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n847), .A2(new_n928), .A3(new_n848), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n847), .B2(new_n848), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n849), .A2(KEYINPUT110), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n847), .A2(new_n928), .A3(new_n848), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n932), .A2(new_n933), .B1(new_n926), .B2(new_n925), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n911), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n932), .A2(new_n933), .A3(new_n926), .A4(new_n925), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n907), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n920), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n892), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n920), .B1(new_n935), .B2(new_n938), .ZN(new_n941));
  OR3_X1    g516(.A1(new_n940), .A2(KEYINPUT43), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n909), .B1(new_n936), .B2(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n906), .A2(new_n903), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n920), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n907), .B2(new_n943), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n946), .A2(new_n892), .A3(new_n939), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  OAI211_X1 g523(.A(KEYINPUT44), .B(new_n942), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n940), .B2(new_n941), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n940), .C2(new_n941), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n946), .A2(new_n948), .A3(new_n892), .A4(new_n939), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n955), .A2(KEYINPUT112), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT112), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n949), .B1(new_n957), .B2(new_n958), .ZN(G397));
  NAND2_X1  g534(.A1(new_n861), .A2(G1996), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n700), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G2067), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n737), .B(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(G164), .B2(G1384), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n465), .A2(new_n467), .A3(G40), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n469), .ZN(new_n970));
  OAI21_X1  g545(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT68), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n970), .B1(new_n973), .B2(new_n472), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n969), .B1(new_n974), .B2(new_n462), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n967), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n965), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n976), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n809), .B(new_n814), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT48), .Z(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n812), .A2(new_n977), .A3(new_n814), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n737), .A2(G2067), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n976), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT46), .B1(new_n976), .B2(new_n961), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n861), .B1(KEYINPUT46), .B2(new_n961), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n993), .A2(new_n964), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n978), .B2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n986), .B(new_n989), .C1(new_n990), .C2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n990), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n490), .B1(new_n476), .B2(new_n492), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n470), .A2(KEYINPUT69), .A3(new_n495), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n499), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n487), .A2(new_n488), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n479), .B2(G126), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n968), .B1(new_n474), .B2(G2105), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1005), .B(new_n1006), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1961), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(new_n975), .ZN(new_n1015));
  INV_X1    g590(.A(G2078), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n967), .A2(new_n1015), .A3(KEYINPUT53), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1006), .B1(G164), .B2(new_n1013), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n1003), .B2(new_n1012), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1018), .A2(new_n1019), .A3(G2078), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1011), .B(new_n1017), .C1(new_n1020), .C2(KEYINPUT53), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n576), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n967), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1023), .A2(new_n1024), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n462), .B1(new_n474), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n1026), .B2(new_n474), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1014), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n968), .A2(new_n1024), .A3(G2078), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n967), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1025), .A2(G301), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT54), .B1(new_n1022), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1007), .B1(new_n1003), .B2(new_n1012), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1035), .A2(G2084), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1966), .B1(new_n967), .B2(new_n1015), .ZN(new_n1038));
  OAI21_X1  g613(.A(G8), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G286), .A2(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G168), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT122), .ZN(new_n1045));
  INV_X1    g620(.A(G1966), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n975), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1049));
  INV_X1    g624(.A(G2084), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n1043), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1034), .A2(new_n1041), .B1(new_n1045), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1039), .A2(KEYINPUT51), .A3(new_n1040), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1033), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n530), .A2(G48), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n503), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n512), .A2(new_n583), .ZN(new_n1062));
  OAI21_X1  g637(.A(G1981), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT115), .B(G1981), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n587), .A2(new_n591), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1042), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1065), .A3(KEYINPUT49), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n781), .A2(G1976), .A3(new_n782), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(G8), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1069), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1071), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT116), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1071), .A2(new_n1075), .A3(new_n1081), .A4(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G303), .A2(G8), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1085));
  XOR2_X1   g660(.A(new_n1084), .B(new_n1085), .Z(new_n1086));
  OAI211_X1 g661(.A(KEYINPUT113), .B(new_n789), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1087));
  INV_X1    g662(.A(G2090), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1048), .A2(new_n1049), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n967), .A2(new_n1015), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT113), .B1(new_n1091), .B2(new_n789), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1086), .B(G8), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n789), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1042), .B1(new_n1094), .B2(new_n1089), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1095), .A2(new_n1086), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1083), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n1011), .A3(new_n1031), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1025), .A2(G301), .A3(new_n1017), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT54), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1057), .A2(new_n1058), .A3(new_n1098), .A4(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1034), .B(G8), .C1(new_n1052), .C2(G286), .ZN(new_n1105));
  AOI211_X1 g680(.A(KEYINPUT122), .B(new_n1040), .C1(new_n1047), .C2(new_n1051), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1053), .B1(new_n1052), .B2(new_n1043), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1056), .B(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n1109));
  AND4_X1   g684(.A1(G301), .A2(new_n1099), .A3(new_n1011), .A4(new_n1031), .ZN(new_n1110));
  AOI21_X1  g685(.A(G301), .B1(new_n1025), .B2(new_n1017), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1112), .A3(new_n1103), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT124), .B1(new_n1113), .B2(new_n1097), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT56), .B(G2072), .Z(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n967), .A2(new_n1015), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1117), .A2(new_n1118), .B1(new_n759), .B2(new_n1009), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n1120));
  XNOR2_X1  g695(.A(G299), .B(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n967), .A2(new_n1015), .A3(KEYINPUT118), .A4(new_n1116), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1126), .A2(new_n1127), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1009), .A2(new_n771), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1006), .A2(new_n1008), .A3(new_n1130), .A4(new_n963), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT119), .B1(new_n1072), .B2(G2067), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1133), .A2(new_n769), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1124), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1121), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1123), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1133), .A2(new_n769), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT60), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n608), .A2(KEYINPUT60), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n967), .A2(new_n1015), .A3(new_n961), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT58), .B(G1341), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n1072), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n843), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(KEYINPUT121), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1133), .A2(new_n1141), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1138), .A2(new_n1140), .A3(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1128), .A2(new_n1123), .A3(new_n1136), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1135), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1104), .A2(new_n1114), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n1155));
  NOR2_X1   g730(.A1(G288), .A2(G1976), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1071), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1065), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1069), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1093), .B2(new_n1079), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1042), .B(G286), .C1(new_n1047), .C2(new_n1051), .ZN(new_n1161));
  AND4_X1   g736(.A1(KEYINPUT63), .A2(new_n1071), .A3(new_n1075), .A4(new_n1078), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1093), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT113), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1094), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1165), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1086), .B1(new_n1166), .B2(G8), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT117), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1052), .A2(G8), .A3(G168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1169), .A2(new_n1079), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(G8), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1086), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1171), .A2(new_n1174), .A3(new_n1175), .A4(new_n1093), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1168), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1170), .B1(new_n1097), .B2(new_n1169), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1160), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1154), .A2(new_n1155), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1155), .B1(new_n1154), .B2(new_n1179), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1111), .B1(new_n1108), .B2(KEYINPUT62), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1097), .B(new_n1182), .C1(KEYINPUT62), .C2(new_n1108), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(G290), .B(G1986), .Z(new_n1185));
  OAI21_X1  g760(.A(new_n981), .B1(new_n978), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n997), .B1(new_n1184), .B2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g762(.A1(new_n460), .A2(G401), .A3(G227), .A4(G229), .ZN(new_n1189));
  INV_X1    g763(.A(new_n893), .ZN(new_n1190));
  INV_X1    g764(.A(new_n894), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g766(.A1(new_n1192), .A2(new_n955), .ZN(G308));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n955), .ZN(G225));
endmodule


