//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT78), .B(G469), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(G143), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT66), .B1(new_n193), .B2(G143), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G143), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n192), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT69), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n197), .A2(new_n207), .A3(KEYINPUT1), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(G128), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n201), .B2(G143), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n204), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G107), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n215), .A2(G107), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  INV_X1    g035(.A(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G104), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n220), .A2(new_n223), .A3(new_n224), .A4(new_n216), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n214), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n219), .A2(new_n225), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g043(.A(G128), .B1(new_n211), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n200), .A2(new_n203), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n228), .B1(new_n231), .B2(new_n204), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT11), .B1(new_n234), .B2(G134), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n238), .A2(new_n234), .A3(KEYINPUT11), .A4(G134), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n234), .A2(KEYINPUT11), .A3(G134), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT68), .B1(new_n241), .B2(G137), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n237), .A2(G131), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  INV_X1    g059(.A(new_n243), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n241), .A2(G137), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n236), .B1(new_n247), .B2(KEYINPUT11), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n235), .A2(KEYINPUT67), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n245), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT77), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n233), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT12), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n256));
  INV_X1    g070(.A(new_n213), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n190), .B1(new_n205), .B2(KEYINPUT69), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(new_n208), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n256), .B1(new_n259), .B2(new_n204), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n198), .B1(new_n201), .B2(G143), .ZN(new_n261));
  AND4_X1   g075(.A1(new_n202), .A2(new_n194), .A3(new_n196), .A4(G143), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n191), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n197), .A2(new_n207), .A3(KEYINPUT1), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n207), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n264), .A2(new_n265), .A3(new_n190), .ZN(new_n266));
  OAI211_X1 g080(.A(KEYINPUT71), .B(new_n263), .C1(new_n266), .C2(new_n257), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT10), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n226), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n260), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n200), .A2(new_n203), .A3(new_n230), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n226), .B1(new_n263), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n273), .B2(KEYINPUT10), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n232), .A2(KEYINPUT76), .A3(new_n268), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n220), .A2(new_n223), .A3(new_n216), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G101), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT4), .A3(new_n225), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n280), .A3(G101), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n200), .A2(new_n203), .ZN(new_n283));
  AND2_X1   g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  OR3_X1    g098(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n283), .A2(new_n284), .B1(new_n213), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n270), .A2(new_n276), .A3(new_n252), .A4(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT12), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n233), .A2(new_n253), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G227), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n255), .A2(new_n290), .A3(new_n292), .A4(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n244), .A2(new_n251), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT76), .B1(new_n232), .B2(new_n268), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n273), .A2(new_n271), .A3(KEYINPUT10), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n289), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n260), .A2(new_n267), .A3(new_n269), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n297), .B1(new_n304), .B2(new_n290), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT79), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n298), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI211_X1 g121(.A(KEYINPUT79), .B(new_n297), .C1(new_n304), .C2(new_n290), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n187), .B(new_n189), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n255), .A2(new_n290), .A3(new_n292), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n290), .A2(new_n297), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n310), .A2(new_n296), .B1(new_n311), .B2(new_n304), .ZN(new_n312));
  OAI21_X1  g126(.A(G469), .B1(new_n312), .B2(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT88), .ZN(new_n318));
  XNOR2_X1  g132(.A(G113), .B(G122), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(new_n215), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT85), .A2(G143), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT85), .A2(G143), .ZN(new_n323));
  NOR2_X1   g137(.A1(G237), .A2(G953), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n322), .A2(new_n323), .B1(new_n324), .B2(G214), .ZN(new_n325));
  INV_X1    g139(.A(G237), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(new_n294), .A3(G214), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n321), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT18), .B(G131), .C1(new_n325), .C2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(G214), .A3(new_n324), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT18), .A2(G131), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT85), .B(G143), .Z(new_n332));
  INV_X1    g146(.A(new_n327), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n330), .B(new_n331), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G125), .B(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n201), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G125), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G146), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n329), .A2(new_n334), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G131), .B1(new_n325), .B2(new_n328), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n330), .B(new_n245), .C1(new_n332), .C2(new_n333), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT17), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(KEYINPUT17), .B(G131), .C1(new_n325), .C2(new_n328), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT16), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n339), .A2(KEYINPUT16), .A3(G140), .ZN(new_n351));
  AOI21_X1  g165(.A(G146), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n351), .A3(G146), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n320), .B(new_n344), .C1(new_n348), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n354), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n345), .B2(new_n346), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT19), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n341), .A2(KEYINPUT86), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT19), .B1(new_n335), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n201), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n334), .A2(new_n343), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n358), .A2(new_n363), .B1(new_n364), .B2(new_n329), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n356), .B1(new_n365), .B2(new_n320), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT87), .ZN(new_n367));
  NOR2_X1   g181(.A1(G475), .A2(G902), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT20), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n368), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(KEYINPUT87), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n356), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(new_n353), .A3(new_n354), .A4(new_n349), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n320), .B1(new_n378), .B2(new_n344), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n187), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G475), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n318), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n371), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT20), .A3(new_n369), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n371), .A2(new_n374), .B1(new_n380), .B2(G475), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT88), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n210), .A2(G128), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n190), .A2(G143), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n241), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G116), .ZN(new_n393));
  INV_X1    g207(.A(G122), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT89), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G122), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n394), .A2(G116), .ZN(new_n399));
  OAI21_X1  g213(.A(G107), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT89), .B(G122), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n222), .B(new_n401), .C1(new_n402), .C2(new_n393), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n392), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT13), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n190), .B2(G143), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n210), .A2(KEYINPUT13), .A3(G128), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n390), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT90), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n408), .A2(new_n409), .A3(G134), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n408), .B2(G134), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n404), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT14), .B1(new_n402), .B2(new_n393), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(G107), .C1(new_n399), .C2(new_n398), .ZN(new_n414));
  OAI221_X1 g228(.A(new_n401), .B1(KEYINPUT14), .B2(new_n222), .C1(new_n402), .C2(new_n393), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT91), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n241), .B1(new_n389), .B2(new_n390), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n416), .B1(new_n392), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n417), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT91), .A3(new_n391), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n414), .A2(new_n415), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G217), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n315), .A2(new_n423), .A3(G953), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n412), .A2(new_n421), .A3(new_n424), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n187), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n388), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G119), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT2), .B(G113), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n437), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT70), .ZN(new_n443));
  OR3_X1    g257(.A1(new_n441), .A2(KEYINPUT70), .A3(new_n437), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n443), .A2(new_n279), .A3(new_n444), .A4(new_n281), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n446));
  INV_X1    g260(.A(G119), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G116), .ZN(new_n448));
  OAI211_X1 g262(.A(G113), .B(new_n448), .C1(new_n438), .C2(new_n446), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n228), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G122), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n445), .A2(new_n450), .A3(new_n452), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n457), .A3(new_n453), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n339), .B(new_n263), .C1(new_n266), .C2(new_n257), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n283), .A2(new_n284), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n213), .A2(new_n287), .ZN(new_n462));
  OAI21_X1  g276(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n294), .A2(G224), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT80), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n465), .B(KEYINPUT81), .Z(new_n466));
  NAND3_X1  g280(.A1(new_n460), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n460), .B2(new_n463), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT82), .B1(new_n459), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n460), .A2(new_n463), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n460), .A2(new_n463), .A3(KEYINPUT84), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n452), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n450), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n228), .B1(new_n442), .B2(new_n449), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n455), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n473), .B1(new_n460), .B2(new_n463), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(G902), .B1(new_n478), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n469), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n467), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(new_n490), .A3(new_n458), .A4(new_n456), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n471), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G210), .B1(G237), .B2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n471), .A2(new_n487), .A3(new_n491), .A4(new_n493), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n436), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n294), .A2(G952), .ZN(new_n498));
  NAND2_X1  g312(.A1(G234), .A2(G237), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT21), .B(G898), .Z(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(G902), .A3(G953), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(KEYINPUT92), .Z(new_n504));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n317), .A2(new_n434), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G234), .ZN(new_n507));
  OAI21_X1  g321(.A(G217), .B1(new_n507), .B2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT74), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n447), .A2(G128), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n447), .A2(G128), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n511), .B(new_n512), .C1(new_n513), .C2(KEYINPUT23), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT24), .B(G110), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n190), .A2(G119), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n517), .A2(new_n511), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n514), .A2(G110), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n352), .B2(new_n357), .ZN(new_n520));
  OAI22_X1  g334(.A1(new_n514), .A2(G110), .B1(new_n516), .B2(new_n518), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n354), .A3(new_n336), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT75), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT22), .B(G137), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n520), .A3(new_n522), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n510), .B1(new_n532), .B2(G902), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(KEYINPUT25), .A3(new_n187), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n509), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n508), .A2(new_n187), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n443), .A2(new_n444), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n288), .B1(new_n244), .B2(new_n251), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n246), .A2(new_n245), .A3(new_n250), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n234), .A2(G134), .ZN(new_n543));
  OAI21_X1  g357(.A(G131), .B1(new_n543), .B2(new_n247), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n541), .B1(new_n214), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n540), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n545), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n260), .A2(new_n267), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n541), .A2(KEYINPUT30), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n541), .A2(new_n540), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n324), .A2(G210), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n556), .B(KEYINPUT27), .Z(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT26), .B(G101), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n557), .B(new_n558), .Z(new_n559));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT31), .ZN(new_n561));
  INV_X1    g375(.A(new_n559), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT28), .ZN(new_n563));
  INV_X1    g377(.A(new_n540), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n546), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n555), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT28), .B1(new_n550), .B2(new_n554), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n562), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n548), .A2(new_n552), .B1(new_n550), .B2(new_n554), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT31), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n559), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n561), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(G472), .A2(G902), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT32), .B1(new_n572), .B2(new_n573), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n540), .B1(new_n550), .B2(new_n541), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT73), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n555), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI211_X1 g393(.A(KEYINPUT73), .B(new_n540), .C1(new_n550), .C2(new_n541), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT28), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n567), .A2(new_n582), .A3(new_n562), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n569), .B2(new_n559), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n566), .A2(new_n567), .A3(new_n562), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n553), .A2(new_n555), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n562), .ZN(new_n590));
  INV_X1    g404(.A(new_n567), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n550), .A2(new_n554), .B1(new_n546), .B2(new_n564), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n591), .B(new_n559), .C1(new_n563), .C2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n590), .A2(new_n593), .A3(KEYINPUT72), .A4(new_n582), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n584), .A2(new_n588), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n539), .B1(new_n576), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n506), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n422), .B2(new_n425), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT93), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n412), .A2(new_n421), .A3(new_n602), .A4(new_n424), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n427), .A2(KEYINPUT93), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT94), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n601), .A2(new_n604), .A3(new_n607), .A4(new_n603), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n428), .A2(new_n600), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n430), .A2(G902), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n606), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n429), .A2(new_n430), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n383), .A2(new_n387), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n497), .A2(new_n614), .A3(new_n504), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT95), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n497), .A2(new_n614), .A3(new_n617), .A4(new_n504), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n572), .A2(new_n187), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G472), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n572), .A2(new_n573), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n538), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n317), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  INV_X1    g441(.A(new_n497), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n372), .A2(new_n382), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n432), .A3(new_n504), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n630), .A2(KEYINPUT96), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(KEYINPUT96), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT98), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT35), .B(G107), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(new_n523), .Z(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n536), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n535), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n621), .A2(new_n622), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT99), .ZN(new_n645));
  INV_X1    g459(.A(new_n316), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n309), .B2(new_n313), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n505), .A2(new_n434), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n621), .A2(new_n649), .A3(new_n622), .A4(new_n643), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n645), .A2(new_n647), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  INV_X1    g467(.A(KEYINPUT32), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n622), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n596), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n385), .A2(new_n386), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n502), .A2(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n500), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n433), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n497), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n657), .A2(new_n647), .A3(new_n643), .A4(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n642), .B1(new_n576), .B2(new_n596), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(KEYINPUT100), .A3(new_n647), .A4(new_n663), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XNOR2_X1  g484(.A(new_n660), .B(KEYINPUT39), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n647), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT40), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n589), .A2(new_n559), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n187), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n579), .A2(new_n559), .A3(new_n580), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n655), .A2(new_n677), .A3(new_n656), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n495), .A2(new_n496), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n383), .A2(new_n387), .A3(new_n432), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n682), .A2(new_n436), .A3(new_n643), .A4(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n673), .A2(new_n678), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n595), .A2(G472), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n655), .A2(new_n656), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n647), .B(new_n643), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n383), .A2(new_n387), .A3(new_n613), .A4(new_n660), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n692), .A2(new_n497), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n693), .B1(new_n692), .B2(new_n497), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n688), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n383), .A2(new_n387), .A3(new_n613), .A4(new_n660), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT102), .B1(new_n628), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n692), .A2(new_n497), .A3(new_n693), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n667), .A3(KEYINPUT103), .A4(new_n647), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(new_n309), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  INV_X1    g520(.A(new_n290), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n274), .A2(new_n275), .B1(new_n288), .B2(new_n282), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n252), .B1(new_n708), .B2(new_n270), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n296), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n255), .A2(new_n292), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n710), .A2(KEYINPUT79), .B1(new_n711), .B2(new_n311), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n305), .A2(new_n306), .ZN(new_n713));
  AOI21_X1  g527(.A(G902), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(G469), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n706), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n187), .B1(new_n307), .B2(new_n308), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(KEYINPUT104), .A3(G469), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n646), .B(new_n705), .C1(new_n716), .C2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n597), .A3(new_n619), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  AOI21_X1  g536(.A(new_n705), .B1(new_n716), .B2(new_n718), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n597), .A2(new_n723), .A3(new_n316), .A4(new_n633), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  INV_X1    g539(.A(new_n504), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n434), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n719), .A2(new_n497), .A3(new_n667), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NOR3_X1   g543(.A1(new_n628), .A2(new_n684), .A3(new_n726), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT105), .B(G472), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n620), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n559), .B1(new_n581), .B2(new_n591), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n561), .A2(new_n571), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n573), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n732), .A2(new_n735), .A3(new_n538), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n723), .A2(new_n730), .A3(new_n736), .A4(new_n316), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT106), .B(G122), .Z(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G24));
  NAND2_X1  g553(.A1(new_n710), .A2(KEYINPUT79), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n713), .A3(new_n298), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n706), .B(new_n715), .C1(new_n741), .C2(new_n187), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT104), .B1(new_n717), .B2(G469), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n316), .B(new_n309), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n628), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n732), .A2(new_n735), .A3(new_n643), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n732), .A2(new_n735), .A3(KEYINPUT107), .A4(new_n643), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n698), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n339), .ZN(G27));
  NOR2_X1   g568(.A1(new_n679), .A2(new_n436), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT108), .B1(new_n317), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n647), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n656), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n572), .A2(KEYINPUT109), .A3(KEYINPUT32), .A4(new_n573), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n575), .B1(new_n595), .B2(G472), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n538), .A3(new_n692), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT42), .B1(new_n760), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n757), .A2(new_n769), .A3(new_n597), .A4(new_n759), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n245), .ZN(G33));
  NAND4_X1  g586(.A1(new_n757), .A2(new_n597), .A3(new_n662), .A4(new_n759), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  OAI21_X1  g588(.A(G469), .B1(new_n312), .B2(KEYINPUT45), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(KEYINPUT45), .B2(new_n312), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(G469), .B2(G902), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n705), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n316), .A3(new_n671), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n613), .ZN(new_n786));
  INV_X1    g600(.A(new_n388), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT43), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n787), .A2(new_n786), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n791), .B1(KEYINPUT43), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n642), .B1(new_n621), .B2(new_n622), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT44), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n755), .B(KEYINPUT113), .Z(new_n797));
  AND2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n785), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  NAND2_X1  g614(.A1(new_n782), .A2(new_n316), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n657), .A2(new_n756), .A3(new_n538), .A4(new_n698), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  XOR2_X1   g620(.A(new_n723), .B(KEYINPUT49), .Z(new_n807));
  NAND4_X1  g621(.A1(new_n790), .A2(new_n538), .A3(new_n316), .A4(new_n435), .ZN(new_n808));
  OR4_X1    g622(.A1(new_n678), .A2(new_n807), .A3(new_n681), .A4(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n793), .A2(new_n499), .A3(new_n498), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n736), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n811), .A2(new_n435), .A3(new_n681), .A4(new_n744), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT50), .Z(new_n813));
  NOR2_X1   g627(.A1(new_n744), .A2(new_n756), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n749), .A2(new_n750), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n678), .A2(new_n539), .A3(new_n500), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n388), .A2(new_n786), .ZN(new_n820));
  OAI22_X1  g634(.A1(new_n815), .A2(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n811), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n723), .A2(new_n646), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n797), .B(new_n823), .C1(new_n803), .C2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(KEYINPUT51), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n766), .A2(new_n538), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n815), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT48), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n819), .A2(new_n388), .A3(new_n786), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n498), .B1(new_n811), .B2(new_n746), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n697), .A2(new_n702), .B1(new_n666), .B2(new_n668), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n497), .A2(new_n683), .A3(new_n642), .A4(new_n660), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n835), .A2(new_n647), .A3(new_n678), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n745), .B2(new_n751), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  AND4_X1   g652(.A1(KEYINPUT52), .A2(new_n703), .A3(new_n669), .A4(new_n837), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT114), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n703), .A2(new_n669), .A3(new_n837), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n834), .A2(KEYINPUT52), .A3(new_n837), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n728), .A2(new_n720), .A3(new_n724), .A4(new_n737), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n771), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n434), .B1(new_n388), .B2(new_n613), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n505), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n506), .A2(new_n597), .B1(new_n624), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n314), .A2(new_n755), .A3(new_n316), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n658), .A2(new_n432), .A3(new_n661), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n667), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n851), .A2(new_n651), .A3(new_n773), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n751), .A2(new_n757), .A3(new_n759), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n848), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n840), .A2(new_n846), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n843), .A2(new_n844), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(KEYINPUT54), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT116), .B1(new_n855), .B2(new_n857), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n624), .A2(new_n850), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n598), .A2(new_n651), .A3(new_n854), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n773), .A4(new_n856), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n868), .A2(new_n848), .A3(new_n872), .A4(KEYINPUT53), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n838), .A2(new_n839), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n860), .B2(new_n863), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n865), .A2(new_n866), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n867), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT51), .B1(new_n822), .B2(new_n825), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n833), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(G952), .A2(G953), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n809), .B1(new_n882), .B2(new_n883), .ZN(G75));
  XNOR2_X1  g698(.A(new_n459), .B(KEYINPUT117), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n470), .B(KEYINPUT55), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n860), .A2(new_n863), .ZN(new_n889));
  INV_X1    g703(.A(new_n875), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT118), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n887), .B(new_n888), .C1(new_n893), .C2(new_n494), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  INV_X1    g709(.A(G210), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(new_n887), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n294), .A2(G952), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n894), .A2(new_n898), .A3(new_n899), .ZN(G51));
  NAND2_X1  g714(.A1(new_n893), .A2(new_n776), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n878), .ZN(new_n904));
  NAND2_X1  g718(.A1(G469), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT57), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n901), .A2(KEYINPUT120), .B1(new_n741), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n899), .B1(new_n902), .B2(new_n908), .ZN(G54));
  NAND3_X1  g723(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n910));
  INV_X1    g724(.A(new_n366), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n899), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .A4(new_n366), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(G60));
  INV_X1    g728(.A(new_n899), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n903), .A2(new_n878), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n917));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT59), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n915), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n917), .B1(new_n880), .B2(new_n919), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G63));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n876), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n929), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n848), .A2(new_n858), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n862), .B2(KEYINPUT114), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n933), .B2(new_n846), .ZN(new_n934));
  OAI211_X1 g748(.A(KEYINPUT122), .B(new_n931), .C1(new_n934), .C2(new_n875), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n930), .A2(new_n935), .A3(new_n532), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n930), .A2(new_n935), .A3(new_n938), .A4(new_n532), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n640), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT122), .B1(new_n891), .B2(new_n931), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n876), .A2(new_n927), .A3(new_n929), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(KEYINPUT61), .A3(new_n915), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n926), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n640), .B1(new_n930), .B2(new_n935), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n899), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(KEYINPUT124), .A3(new_n937), .A4(new_n939), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n944), .A2(new_n915), .A3(new_n936), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n948), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(G66));
  NAND3_X1  g768(.A1(new_n501), .A2(G224), .A3(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n847), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n651), .A3(new_n851), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n957), .B2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n885), .B1(G898), .B2(new_n294), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(G69));
  NAND2_X1  g774(.A1(new_n546), .A2(new_n547), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n552), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n360), .A2(new_n362), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(G900), .B2(G953), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n768), .A2(new_n770), .A3(new_n773), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n799), .A2(new_n805), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n834), .B1(new_n746), .B2(new_n752), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n827), .A2(new_n628), .A3(new_n684), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT126), .B1(new_n785), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n785), .A2(new_n971), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n967), .B(new_n970), .C1(new_n972), .C2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n965), .B1(new_n976), .B2(G953), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n756), .A2(new_n849), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n597), .A2(new_n672), .A3(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n799), .A2(new_n805), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n970), .A2(new_n686), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n984), .A2(new_n294), .ZN(new_n985));
  INV_X1    g799(.A(new_n964), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n977), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n976), .B2(new_n957), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n589), .A2(new_n559), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n674), .ZN(new_n995));
  INV_X1    g809(.A(new_n991), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n861), .A2(new_n864), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n915), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n991), .B1(new_n984), .B2(new_n957), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n995), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n1001), .A2(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(KEYINPUT127), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(G57));
endmodule


