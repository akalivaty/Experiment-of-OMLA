//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT65), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT65), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n220), .A2(G1), .A3(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G20), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n204), .A2(G50), .A3(new_n205), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n216), .A2(new_n217), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G116), .ZN(new_n228));
  INV_X1    g0028(.A(G270), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n231));
  INV_X1    g0031(.A(G238), .ZN(new_n232));
  INV_X1    g0032(.A(G97), .ZN(new_n233));
  INV_X1    g0033(.A(G257), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n231), .B1(new_n203), .B2(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n230), .B(new_n235), .C1(G58), .C2(G232), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n236), .A2(new_n212), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT1), .Z(new_n238));
  AOI211_X1 g0038(.A(new_n226), .B(new_n238), .C1(new_n217), .C2(new_n216), .ZN(G361));
  XOR2_X1   g0039(.A(G226), .B(G232), .Z(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G264), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n229), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  INV_X1    g0048(.A(G107), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G97), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n233), .A2(G107), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G87), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(new_n228), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT67), .ZN(new_n256));
  XNOR2_X1  g0056(.A(G50), .B(G68), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(G58), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(new_n207), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n256), .B(new_n259), .ZN(G351));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n222), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT7), .B1(new_n267), .B2(new_n211), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT7), .ZN(new_n269));
  AOI211_X1 g0069(.A(new_n269), .B(G20), .C1(new_n264), .C2(new_n266), .ZN(new_n270));
  OAI21_X1  g0070(.A(G68), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(G20), .B1(G159), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT16), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n262), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT78), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT78), .B1(new_n264), .B2(new_n266), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n211), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n270), .B1(new_n280), .B2(new_n269), .ZN(new_n281));
  OAI211_X1 g0081(.A(KEYINPUT16), .B(new_n274), .C1(new_n281), .C2(new_n203), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n211), .B2(G1), .ZN(new_n290));
  AND4_X1   g0090(.A1(new_n222), .A2(new_n261), .A3(new_n286), .A4(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n210), .A2(KEYINPUT69), .A3(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(new_n293), .B2(new_n285), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n283), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G41), .A2(G45), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT68), .B1(new_n297), .B2(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(G1), .A3(G13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT68), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n210), .C1(G41), .C2(G45), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n298), .A2(G232), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n304));
  INV_X1    g0104(.A(G274), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n219), .A2(new_n221), .A3(new_n299), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n264), .A2(new_n266), .A3(G226), .A4(G1698), .ZN(new_n310));
  INV_X1    g0110(.A(G1698), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n264), .A2(new_n266), .A3(G223), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G87), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n308), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT79), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n303), .A2(new_n307), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n309), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n315), .B2(G169), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(KEYINPUT79), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n296), .A2(new_n322), .A3(KEYINPUT18), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT18), .B1(new_n296), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(KEYINPUT80), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n318), .A2(new_n319), .A3(new_n316), .ZN(new_n326));
  AOI21_X1  g0126(.A(G169), .B1(new_n318), .B2(new_n319), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT79), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT79), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n294), .B1(new_n277), .B2(new_n282), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT18), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT80), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n318), .A2(new_n319), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G200), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n315), .A2(G190), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n332), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT17), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT17), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n332), .A2(new_n343), .A3(new_n339), .A4(new_n340), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n325), .A2(new_n337), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT3), .B(G33), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(G232), .A3(new_n311), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n267), .A2(G107), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(G1698), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n348), .C1(new_n349), .C2(new_n232), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n309), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G244), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n307), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n316), .ZN(new_n357));
  INV_X1    g0157(.A(new_n273), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n284), .A2(new_n358), .B1(new_n211), .B2(new_n207), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT70), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n211), .A2(G33), .ZN(new_n362));
  OR3_X1    g0162(.A1(new_n361), .A2(KEYINPUT71), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT70), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n364), .B1(new_n211), .B2(new_n207), .C1(new_n284), .C2(new_n358), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT71), .B1(new_n361), .B2(new_n362), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n360), .A2(new_n363), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n222), .A2(new_n261), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n367), .A2(new_n368), .B1(new_n207), .B2(new_n287), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n291), .A2(G77), .A3(new_n292), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n355), .A2(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n357), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n346), .A2(G226), .A3(new_n311), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n346), .A2(G232), .A3(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G97), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n309), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n353), .A2(G238), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n307), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT13), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n306), .B1(new_n379), .B2(new_n309), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n381), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n375), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT76), .B1(new_n293), .B2(new_n203), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n291), .A2(new_n389), .A3(G68), .A4(new_n292), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n211), .A2(G33), .A3(G77), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n203), .A2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n393), .B1(new_n392), .B2(new_n394), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n273), .A2(G50), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n262), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g0200(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n401));
  INV_X1    g0201(.A(KEYINPUT12), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n213), .A2(G1), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(G20), .A3(new_n203), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n400), .A2(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n404), .A2(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(new_n397), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n399), .A3(new_n395), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n368), .ZN(new_n409));
  INV_X1    g0209(.A(new_n401), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n391), .A2(new_n405), .A3(new_n406), .A4(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n387), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n384), .A2(new_n385), .A3(new_n381), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n385), .B1(new_n384), .B2(new_n381), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G190), .ZN(new_n417));
  OAI21_X1  g0217(.A(G169), .B1(new_n414), .B2(new_n415), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(G179), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n383), .A2(new_n386), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT14), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(G169), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT77), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n412), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n400), .A2(new_n401), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n404), .A2(new_n402), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n427), .A2(new_n411), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n429), .A2(KEYINPUT77), .A3(new_n406), .A4(new_n391), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  AOI221_X4 g0231(.A(new_n374), .B1(new_n413), .B2(new_n417), .C1(new_n424), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n345), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n273), .A2(G150), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n434), .B1(new_n284), .B2(new_n362), .C1(new_n206), .C2(new_n211), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n368), .ZN(new_n436));
  INV_X1    g0236(.A(G50), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n287), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n291), .A2(G50), .A3(new_n292), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT73), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n435), .A2(new_n368), .B1(new_n437), .B2(new_n287), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(KEYINPUT73), .A3(new_n439), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT9), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n346), .A2(G222), .A3(new_n311), .ZN(new_n447));
  INV_X1    g0247(.A(G223), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n447), .B1(new_n207), .B2(new_n346), .C1(new_n349), .C2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n306), .B1(new_n449), .B2(new_n309), .ZN(new_n450));
  INV_X1    g0250(.A(G226), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n352), .ZN(new_n452));
  INV_X1    g0252(.A(G190), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT9), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n442), .A2(new_n455), .A3(new_n444), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(G200), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n446), .A2(new_n454), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT10), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n445), .A2(KEYINPUT9), .B1(G200), .B2(new_n452), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT10), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n454), .A4(new_n456), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n452), .A2(G179), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n452), .A2(new_n372), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n440), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT72), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n355), .A2(G200), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n469), .B2(new_n371), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n356), .A2(G190), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n468), .A2(new_n369), .A3(KEYINPUT72), .A4(new_n370), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n463), .A2(new_n466), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT81), .B1(new_n433), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n466), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n476), .B(new_n477), .C1(new_n459), .C2(new_n462), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT81), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n345), .A4(new_n432), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(G41), .ZN(new_n484));
  INV_X1    g0284(.A(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(G274), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n210), .B(G45), .C1(new_n485), .C2(KEYINPUT5), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT92), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n264), .A2(new_n266), .A3(G257), .A4(G1698), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n264), .A2(new_n266), .A3(G250), .A4(new_n311), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G294), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n494), .A2(new_n309), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n483), .A2(G41), .ZN(new_n496));
  OAI211_X1 g0296(.A(G264), .B(new_n300), .C1(new_n488), .C2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT91), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n483), .A2(G41), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n485), .A2(KEYINPUT5), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(new_n210), .A4(G45), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(KEYINPUT91), .A3(G264), .A4(new_n300), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n490), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n494), .A2(new_n309), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(KEYINPUT92), .A3(new_n499), .A4(new_n503), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n489), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G179), .ZN(new_n509));
  INV_X1    g0309(.A(new_n489), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n510), .A3(new_n497), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G169), .ZN(new_n512));
  INV_X1    g0312(.A(new_n403), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n249), .A2(G20), .ZN(new_n514));
  OR3_X1    g0314(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT25), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT25), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n210), .A2(G33), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n222), .A2(new_n261), .A3(new_n286), .A4(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n515), .B(new_n516), .C1(new_n518), .C2(new_n249), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT90), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n346), .A2(new_n211), .A3(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT22), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n346), .A2(new_n524), .A3(new_n211), .A4(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n527));
  XOR2_X1   g0327(.A(new_n514), .B(KEYINPUT23), .Z(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n526), .A2(KEYINPUT24), .A3(new_n527), .A4(new_n528), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n368), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n509), .A2(new_n512), .B1(new_n521), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n499), .A2(new_n503), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT92), .B1(new_n535), .B2(new_n506), .ZN(new_n536));
  INV_X1    g0336(.A(new_n507), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n510), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(KEYINPUT93), .A3(new_n375), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT93), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n508), .B2(G200), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n511), .A2(G190), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n533), .A2(new_n521), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n534), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n286), .A2(G97), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n518), .A2(new_n233), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n358), .A2(new_n207), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n250), .A2(new_n251), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n249), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(KEYINPUT82), .B(new_n550), .C1(new_n554), .C2(new_n211), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n211), .B1(new_n552), .B2(new_n553), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n549), .ZN(new_n558));
  OAI21_X1  g0358(.A(G107), .B1(new_n268), .B2(new_n270), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI211_X1 g0360(.A(new_n547), .B(new_n548), .C1(new_n560), .C2(new_n368), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n264), .A2(new_n266), .A3(G244), .A4(new_n311), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(KEYINPUT4), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n346), .A2(G244), .A3(new_n311), .A4(new_n564), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n346), .A2(G250), .A3(G1698), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G283), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n563), .A2(KEYINPUT4), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n309), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT85), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n300), .B1(new_n488), .B2(new_n496), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(new_n234), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n502), .A2(KEYINPUT85), .A3(G257), .A4(new_n300), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n489), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(G190), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n572), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n576), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT86), .B1(new_n580), .B2(new_n510), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT86), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n582), .B(new_n489), .C1(new_n575), .C2(new_n576), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n561), .B(new_n578), .C1(new_n584), .C2(new_n375), .ZN(new_n585));
  INV_X1    g0385(.A(new_n581), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n577), .A2(KEYINPUT86), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(new_n316), .A3(new_n572), .A4(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n547), .B1(new_n560), .B2(new_n368), .ZN(new_n589));
  INV_X1    g0389(.A(new_n548), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n572), .A2(new_n577), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n372), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n588), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n346), .A2(G257), .A3(new_n311), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n346), .A2(G264), .A3(G1698), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n267), .A2(G303), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n309), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n502), .A2(G270), .A3(new_n300), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n600), .A2(new_n510), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n228), .A2(G20), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n513), .A2(new_n603), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n222), .A2(new_n261), .A3(new_n286), .A4(new_n517), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(G116), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n263), .A2(G97), .ZN(new_n607));
  AOI21_X1  g0407(.A(G20), .B1(G33), .B2(G283), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n222), .A2(new_n261), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n609), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT20), .B1(new_n609), .B2(new_n603), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n602), .A2(new_n612), .A3(KEYINPUT89), .A4(G179), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT89), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n518), .A2(new_n228), .B1(new_n513), .B2(new_n603), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n607), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n368), .A2(new_n603), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT20), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n609), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n600), .A2(G179), .A3(new_n601), .A4(new_n510), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n614), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(new_n620), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n372), .B1(new_n625), .B2(new_n606), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n600), .A2(new_n510), .A3(new_n601), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(KEYINPUT21), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n612), .A2(G169), .A3(new_n627), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(G200), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n632), .B(new_n621), .C1(new_n453), .C2(new_n627), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n624), .A2(new_n628), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n210), .A2(G45), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n300), .A2(G250), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n264), .A2(new_n266), .A3(G238), .A4(new_n311), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n264), .A2(new_n266), .A3(G244), .A4(G1698), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n638), .B(new_n639), .C1(new_n263), .C2(new_n228), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n640), .B2(new_n309), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n635), .A2(new_n305), .ZN(new_n642));
  XOR2_X1   g0442(.A(new_n642), .B(KEYINPUT87), .Z(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G190), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(G200), .ZN(new_n647));
  AND2_X1   g0447(.A1(KEYINPUT88), .A2(G87), .ZN(new_n648));
  NOR2_X1   g0448(.A1(KEYINPUT88), .A2(G87), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n233), .B(new_n249), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT19), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n211), .B1(new_n378), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n346), .A2(new_n211), .A3(G68), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n211), .A2(G33), .A3(G97), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n651), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n368), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n518), .A2(new_n253), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n361), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n286), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n658), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n646), .A2(new_n647), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n645), .A2(new_n316), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n658), .B(new_n663), .C1(new_n361), .C2(new_n518), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n644), .A2(new_n372), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n634), .A2(new_n670), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n481), .A2(new_n546), .A3(new_n595), .A4(new_n671), .ZN(G372));
  NAND2_X1  g0472(.A1(new_n323), .A2(new_n336), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n424), .A2(new_n431), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n413), .A2(new_n417), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n374), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n342), .A2(new_n344), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n673), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n476), .B1(new_n680), .B2(new_n463), .ZN(new_n681));
  INV_X1    g0481(.A(new_n481), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n543), .A2(new_n545), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n647), .A2(new_n664), .A3(KEYINPUT94), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT94), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n375), .B1(new_n641), .B2(new_n643), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n658), .A2(new_n660), .A3(new_n663), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n684), .A2(new_n688), .A3(new_n646), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n669), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI211_X1 g0491(.A(new_n316), .B(new_n489), .C1(new_n505), .C2(new_n507), .ZN(new_n692));
  INV_X1    g0492(.A(new_n512), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n544), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT21), .B1(new_n626), .B2(new_n627), .ZN(new_n695));
  AND4_X1   g0495(.A1(KEYINPUT21), .A2(new_n612), .A3(G169), .A4(new_n627), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n697), .A3(new_n624), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n683), .A2(new_n595), .A3(new_n691), .A4(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n669), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n690), .A2(new_n594), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT26), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT26), .B1(new_n670), .B2(new_n594), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n681), .B1(new_n682), .B2(new_n706), .ZN(G369));
  NAND2_X1  g0507(.A1(new_n697), .A2(new_n624), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n403), .A2(new_n211), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n711), .A2(G213), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n708), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n683), .B(new_n694), .C1(new_n545), .C2(new_n717), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n534), .A2(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT96), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT96), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n723), .A3(new_n720), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n718), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n694), .A2(new_n716), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n722), .A2(new_n724), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n717), .A2(new_n621), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n708), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n634), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n727), .A2(new_n734), .ZN(G399));
  OR2_X1    g0535(.A1(new_n650), .A2(G116), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n214), .A2(G41), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n736), .A2(new_n210), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT97), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT97), .ZN(new_n740));
  INV_X1    g0540(.A(new_n737), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n739), .B(new_n740), .C1(new_n225), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n546), .A2(new_n595), .A3(new_n671), .A4(new_n717), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n592), .A2(new_n622), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n644), .B1(new_n505), .B2(new_n507), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT30), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n627), .A2(new_n644), .A3(new_n316), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n508), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n749), .B(new_n750), .C1(new_n584), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n716), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(KEYINPUT31), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G330), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n705), .A2(new_n717), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT29), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR3_X1    g0563(.A1(new_n670), .A2(new_n594), .A3(KEYINPUT26), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n561), .B1(new_n316), .B2(new_n584), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n765), .A2(new_n593), .A3(new_n669), .A4(new_n689), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n700), .B1(new_n766), .B2(KEYINPUT26), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n585), .A2(new_n594), .A3(KEYINPUT98), .ZN(new_n768));
  AOI21_X1  g0568(.A(KEYINPUT98), .B1(new_n585), .B2(new_n594), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n683), .A2(new_n691), .A3(new_n698), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n764), .B(new_n767), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(KEYINPUT29), .A3(new_n717), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n760), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n743), .B1(new_n774), .B2(G1), .ZN(G364));
  NOR2_X1   g0575(.A1(new_n731), .A2(G330), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT99), .Z(new_n777));
  NOR2_X1   g0577(.A1(new_n213), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n210), .B1(new_n778), .B2(G45), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n741), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n732), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT78), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n267), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n346), .A2(KEYINPUT78), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n214), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n225), .A2(G45), .ZN(new_n788));
  INV_X1    g0588(.A(G45), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n787), .B(new_n788), .C1(new_n259), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n215), .A2(G355), .A3(new_n346), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n791), .C1(G116), .C2(new_n215), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n222), .B1(G20), .B2(new_n372), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n316), .A2(G200), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT101), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n211), .A2(new_n453), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n211), .A2(G190), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G179), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n346), .B(new_n804), .C1(G329), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n316), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G311), .ZN(new_n813));
  NAND3_X1  g0613(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n453), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G326), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n211), .B1(new_n806), .B2(G190), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n814), .A2(G190), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT33), .B(G317), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n801), .A2(new_n810), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n800), .A2(new_n805), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n828), .A2(G322), .B1(new_n830), .B2(G283), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n809), .A2(new_n813), .A3(new_n822), .A4(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n815), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n346), .B1(new_n833), .B2(new_n437), .ZN(new_n834));
  INV_X1    g0634(.A(new_n820), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n835), .A2(new_n203), .B1(new_n818), .B2(new_n233), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(G77), .C2(new_n812), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n802), .A2(new_n649), .A3(new_n648), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n828), .B2(G58), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n837), .B(new_n839), .C1(new_n249), .C2(new_n829), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n808), .A2(G159), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT32), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n832), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n780), .B1(new_n843), .B2(new_n793), .ZN(new_n844));
  INV_X1    g0644(.A(new_n796), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n798), .B(new_n844), .C1(new_n731), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n781), .A2(new_n846), .ZN(G396));
  NAND2_X1  g0647(.A1(new_n374), .A2(new_n716), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n371), .A2(new_n716), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n374), .A2(KEYINPUT102), .ZN(new_n850));
  AND4_X1   g0650(.A1(KEYINPUT102), .A2(new_n357), .A3(new_n371), .A4(new_n373), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n473), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n761), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n477), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n705), .A2(new_n717), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n760), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n780), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n793), .A2(new_n794), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n207), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n820), .A2(G150), .B1(new_n815), .B2(G137), .ZN(new_n862));
  INV_X1    g0662(.A(G159), .ZN(new_n863));
  INV_X1    g0663(.A(G143), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n863), .B2(new_n811), .C1(new_n827), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT34), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n829), .A2(new_n203), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n786), .B1(new_n202), .B2(new_n818), .ZN(new_n868));
  INV_X1    g0668(.A(new_n802), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n867), .B(new_n868), .C1(G50), .C2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(G132), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n866), .B(new_n870), .C1(new_n871), .C2(new_n807), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n267), .B1(new_n811), .B2(new_n228), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n828), .B2(G294), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n808), .A2(G311), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G87), .A2(new_n830), .B1(new_n869), .B2(G107), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n818), .A2(new_n233), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n833), .A2(new_n803), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n877), .B(new_n878), .C1(G283), .C2(new_n820), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n780), .B1(new_n881), .B2(new_n793), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n852), .A2(new_n848), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n861), .B(new_n882), .C1(new_n883), .C2(new_n795), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n859), .A2(new_n884), .ZN(G384));
  AND2_X1   g0685(.A1(new_n413), .A2(new_n417), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n431), .B(new_n716), .C1(new_n886), .C2(new_n424), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n431), .A2(new_n716), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n674), .A2(new_n676), .A3(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n887), .A2(new_n889), .B1(new_n852), .B2(new_n848), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n755), .A2(new_n890), .A3(new_n756), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(KEYINPUT40), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n296), .A2(new_n322), .ZN(new_n894));
  INV_X1    g0694(.A(new_n714), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n296), .A2(new_n895), .ZN(new_n896));
  AND4_X1   g0696(.A1(new_n893), .A2(new_n894), .A3(new_n896), .A4(new_n341), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n282), .A2(new_n368), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT7), .B1(new_n785), .B2(new_n211), .ZN(new_n899));
  OAI21_X1  g0699(.A(G68), .B1(new_n899), .B2(new_n270), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT16), .B1(new_n900), .B2(new_n274), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n295), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n338), .A2(new_n372), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n329), .B1(new_n903), .B2(new_n320), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n714), .B1(new_n904), .B2(new_n317), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n893), .B1(new_n906), .B2(new_n341), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n897), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n894), .A2(KEYINPUT80), .A3(new_n333), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n678), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n902), .A2(new_n895), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT103), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n894), .A2(new_n896), .A3(new_n893), .A4(new_n341), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n906), .A2(new_n341), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n893), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT38), .B(new_n918), .C1(new_n345), .C2(new_n912), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n345), .B2(new_n912), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n915), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n894), .A2(new_n896), .A3(new_n341), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(new_n893), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n896), .B1(new_n678), .B2(new_n673), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n919), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n757), .A2(new_n929), .A3(new_n890), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n892), .A2(new_n924), .B1(new_n930), .B2(KEYINPUT40), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n682), .A2(new_n758), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(G330), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT104), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n887), .A2(new_n889), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n854), .A2(new_n717), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n856), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n924), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n673), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n714), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n929), .A2(KEYINPUT39), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n924), .B2(KEYINPUT39), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n675), .A2(new_n717), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n939), .B(new_n941), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n481), .A2(new_n763), .A3(new_n773), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n681), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n945), .B(new_n947), .Z(new_n948));
  XNOR2_X1  g0748(.A(new_n935), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n210), .B2(new_n778), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT35), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n224), .B1(new_n951), .B2(new_n554), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(G116), .C1(new_n951), .C2(new_n554), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT36), .ZN(new_n954));
  OAI21_X1  g0754(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n225), .A2(new_n955), .B1(G50), .B2(new_n203), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n213), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n950), .A2(new_n954), .A3(new_n957), .ZN(G367));
  XNOR2_X1  g0758(.A(new_n737), .B(KEYINPUT41), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n722), .A2(new_n724), .A3(new_n718), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n960), .A2(new_n733), .ZN(new_n961));
  INV_X1    g0761(.A(new_n718), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n728), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n960), .A2(new_n733), .ZN(new_n964));
  AND4_X1   g0764(.A1(KEYINPUT107), .A2(new_n961), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n961), .A2(new_n964), .B1(KEYINPUT107), .B2(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n774), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n726), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n768), .A2(new_n769), .B1(new_n561), .B2(new_n717), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n765), .A2(new_n593), .A3(new_n716), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n727), .B2(new_n972), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT108), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n734), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n969), .B2(new_n973), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n725), .A2(new_n973), .A3(new_n981), .A4(new_n726), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n734), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n978), .A2(new_n980), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT45), .B1(new_n727), .B2(new_n972), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n975), .B(new_n977), .C1(new_n989), .C2(new_n983), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(new_n979), .A3(new_n734), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n967), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n774), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n959), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n779), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT42), .B1(new_n963), .B2(new_n973), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n594), .B1(new_n970), .B2(new_n694), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n717), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT42), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n725), .A2(new_n999), .A3(new_n972), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n716), .A2(new_n687), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n691), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n669), .B2(new_n1002), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1001), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n986), .A2(new_n972), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1007), .A2(new_n1008), .B1(KEYINPUT105), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(KEYINPUT105), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(KEYINPUT105), .B(new_n1009), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n995), .A2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n828), .A2(G150), .B1(new_n830), .B2(G77), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n808), .A2(G137), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n818), .A2(new_n203), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n833), .A2(new_n864), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(G159), .C2(new_n820), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n346), .B1(new_n811), .B2(new_n437), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n869), .B2(G58), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G283), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n785), .B1(new_n1025), .B2(new_n811), .C1(new_n827), .C2(new_n803), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G97), .B2(new_n830), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n869), .A2(G116), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT46), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n835), .A2(new_n817), .B1(new_n818), .B2(new_n249), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G311), .B2(new_n815), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(G317), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n807), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1024), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n780), .B1(new_n1036), .B2(new_n793), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n787), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n797), .B1(new_n215), .B2(new_n361), .C1(new_n247), .C2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(new_n845), .C2(new_n1004), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT109), .Z(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1016), .A2(new_n1042), .ZN(G387));
  OR3_X1    g0843(.A1(new_n965), .A2(new_n774), .A3(new_n966), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n737), .A3(new_n967), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n779), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n965), .B2(new_n966), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1038), .B1(new_n244), .B2(G45), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n736), .A2(new_n215), .A3(new_n346), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n284), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n789), .C1(new_n203), .C2(new_n207), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1048), .A2(new_n1049), .B1(new_n736), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n214), .A2(new_n249), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n796), .B(new_n793), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n820), .A2(G311), .B1(new_n815), .B2(G322), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n803), .B2(new_n811), .C1(new_n827), .C2(new_n1033), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT48), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n1025), .B2(new_n818), .C1(new_n817), .C2(new_n802), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT49), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n808), .A2(G326), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n786), .B1(new_n830), .B2(G116), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n827), .A2(new_n437), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n818), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n661), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n833), .B2(new_n863), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n285), .B2(new_n820), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n869), .A2(G77), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n785), .B1(G68), .B2(new_n812), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n830), .A2(G97), .B1(G150), .B2(new_n808), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1065), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n780), .B(new_n1055), .C1(new_n1075), .C2(new_n793), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT110), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n728), .B2(new_n845), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1045), .A2(new_n1047), .A3(new_n1078), .ZN(G393));
  NAND2_X1  g0879(.A1(new_n973), .A2(new_n796), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n797), .B1(new_n233), .B2(new_n215), .C1(new_n255), .C2(new_n1038), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n828), .A2(G311), .B1(G317), .B2(new_n815), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  OAI22_X1  g0883(.A1(new_n249), .A2(new_n829), .B1(new_n802), .B2(new_n1025), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n346), .B1(new_n808), .B2(G322), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n228), .B2(new_n818), .C1(new_n835), .C2(new_n803), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1083), .B(new_n1087), .C1(new_n817), .C2(new_n811), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n811), .A2(new_n284), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n828), .A2(G159), .B1(G150), .B2(new_n815), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(KEYINPUT51), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n203), .A2(new_n802), .B1(new_n829), .B2(new_n253), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n786), .B1(new_n864), .B2(new_n807), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n835), .A2(new_n437), .B1(new_n818), .B2(new_n207), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n1092), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1088), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n780), .B1(new_n1098), .B2(new_n793), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1080), .A2(new_n1081), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n988), .A2(new_n991), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n1046), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n988), .A2(new_n991), .A3(new_n967), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n737), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(new_n992), .ZN(G390));
  NAND3_X1  g0905(.A1(new_n772), .A2(new_n717), .A3(new_n855), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n937), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n936), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n944), .B(KEYINPUT111), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n929), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1108), .A2(KEYINPUT112), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT112), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n936), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1106), .B2(new_n937), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n929), .A2(new_n1109), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n924), .A2(KEYINPUT39), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n938), .A2(new_n936), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n944), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n942), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n755), .A2(new_n890), .A3(G330), .A4(new_n756), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(KEYINPUT113), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1117), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n481), .A2(G330), .A3(new_n757), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n946), .A2(new_n1128), .A3(new_n681), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT114), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT114), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n946), .A2(new_n1128), .A3(new_n1131), .A4(new_n681), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n755), .A2(new_n883), .A3(G330), .A4(new_n756), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1113), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(new_n937), .A3(new_n1106), .A4(new_n1123), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1134), .A2(new_n1123), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n938), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1130), .A2(new_n1132), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1127), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n737), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n943), .A2(new_n794), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n828), .A2(G132), .B1(G128), .B2(new_n815), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT115), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT54), .B(G143), .Z(new_n1147));
  NAND2_X1  g0947(.A1(new_n812), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(G150), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n802), .A2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT53), .ZN(new_n1151));
  INV_X1    g0951(.A(G137), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n835), .A2(new_n1152), .B1(new_n818), .B2(new_n863), .ZN(new_n1153));
  INV_X1    g0953(.A(G125), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n346), .B1(new_n807), .B2(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(new_n830), .C2(G50), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1146), .A2(new_n1148), .A3(new_n1151), .A4(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT116), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n820), .A2(G107), .B1(new_n815), .B2(G283), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n207), .B2(new_n818), .C1(new_n817), .C2(new_n807), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n867), .B(new_n1160), .C1(G116), .C2(new_n828), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n267), .B1(new_n802), .B2(new_n253), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT117), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(new_n233), .C2(new_n811), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT118), .Z(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n780), .B1(new_n1166), .B2(new_n793), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1144), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n284), .B2(new_n860), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1124), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1117), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1169), .B1(new_n1174), .B2(new_n1046), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1143), .A2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(KEYINPUT119), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT56), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT55), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n463), .A2(new_n466), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n445), .A2(new_n714), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1181), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n463), .A2(new_n466), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1179), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(new_n463), .B2(new_n466), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n476), .B(new_n1181), .C1(new_n459), .C2(new_n462), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1186), .A2(new_n1187), .A3(KEYINPUT55), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1178), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1182), .A2(new_n1179), .A3(new_n1184), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT55), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n1191), .A3(KEYINPUT56), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n931), .A2(new_n1193), .A3(new_n759), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n924), .A2(new_n892), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n929), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT40), .B1(new_n1197), .B2(new_n891), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1199), .B2(G330), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1194), .A2(new_n1200), .A3(new_n945), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n944), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1202), .A2(new_n1203), .B1(new_n940), .B2(new_n714), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1193), .B1(new_n931), .B2(new_n759), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1199), .A2(G330), .A3(new_n1195), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n939), .A2(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1177), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n945), .B1(new_n1194), .B2(new_n1200), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1204), .A2(new_n1205), .A3(new_n939), .A4(new_n1206), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(KEYINPUT119), .A3(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1046), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n860), .A2(new_n437), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n830), .A2(G58), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G41), .B1(new_n812), .B2(new_n661), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n808), .A2(G283), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1071), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n786), .A2(new_n1019), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n233), .B2(new_n835), .C1(new_n228), .C2(new_n833), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(G107), .C2(new_n828), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT58), .Z(new_n1221));
  AOI22_X1  g1021(.A1(new_n828), .A2(G128), .B1(new_n869), .B2(new_n1147), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n811), .A2(new_n1152), .B1(new_n818), .B2(new_n1149), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G132), .B2(new_n820), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(new_n1154), .C2(new_n833), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT59), .Z(new_n1226));
  AOI21_X1  g1026(.A(G41), .B1(new_n830), .B2(G159), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G33), .B1(new_n808), .B2(G124), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G41), .B1(new_n786), .B2(G33), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1221), .B(new_n1229), .C1(G50), .C2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n780), .B1(new_n1231), .B2(new_n793), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1213), .B(new_n1232), .C1(new_n1195), .C2(new_n795), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1212), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1142), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1208), .A2(new_n1211), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1235), .B1(new_n1174), .B2(new_n1138), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n737), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1234), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(G375));
  OAI221_X1 g1046(.A(new_n1068), .B1(new_n833), .B2(new_n817), .C1(new_n228), .C2(new_n835), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n827), .A2(new_n1025), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n267), .B1(new_n807), .B2(new_n803), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n829), .A2(new_n207), .B1(new_n249), .B2(new_n811), .ZN(new_n1250));
  OR4_X1    g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n802), .A2(new_n233), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n802), .A2(new_n863), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n828), .A2(G137), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n830), .A2(G58), .B1(G128), .B2(new_n808), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n833), .A2(new_n871), .B1(new_n818), .B2(new_n437), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n820), .B2(new_n1147), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n785), .B1(G150), .B2(new_n812), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1251), .A2(new_n1252), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n780), .B1(new_n1260), .B2(new_n793), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n936), .B2(new_n795), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n203), .B2(new_n860), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1138), .B2(new_n1046), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1138), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n959), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1264), .B1(new_n1267), .B2(new_n1139), .ZN(G381));
  INV_X1    g1068(.A(G378), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1245), .A2(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  INV_X1    g1071(.A(G384), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT120), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1270), .A2(new_n1274), .A3(G387), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G390), .A2(G381), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(G407));
  OAI211_X1 g1077(.A(G407), .B(G213), .C1(G343), .C2(new_n1270), .ZN(G409));
  NAND2_X1  g1078(.A1(new_n715), .A2(G213), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1208), .A2(new_n1237), .A3(new_n959), .A4(new_n1211), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1046), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1143), .A2(new_n1175), .A3(new_n1233), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1279), .B(new_n1284), .C1(new_n1245), .C2(new_n1269), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1140), .B1(new_n1266), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n737), .B1(new_n1265), .B2(KEYINPUT60), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1264), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1272), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G384), .B(new_n1264), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n715), .A2(KEYINPUT121), .A3(G213), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n715), .A2(G213), .A3(G2897), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1294), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1290), .A2(new_n1296), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1243), .B1(new_n1239), .B2(new_n1238), .ZN(new_n1300));
  OAI21_X1  g1100(.A(G378), .B1(new_n1300), .B2(new_n1234), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1282), .A2(new_n1283), .B1(G213), .B2(new_n715), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1301), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT62), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1301), .A2(new_n1302), .A3(new_n1307), .A4(new_n1304), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1299), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT124), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1271), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(G393), .A2(G396), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G390), .B1(new_n1016), .B2(new_n1042), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT122), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1311), .B(new_n1312), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1016), .A2(new_n1042), .A3(G390), .ZN(new_n1316));
  INV_X1    g1116(.A(G390), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1014), .B1(new_n994), .B2(new_n779), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(new_n1041), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1315), .A2(new_n1320), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1271), .B1(new_n1319), .B2(KEYINPUT122), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(new_n1312), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT124), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1299), .A2(new_n1306), .A3(new_n1326), .A4(new_n1308), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1310), .A2(new_n1325), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1321), .A2(new_n1324), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(KEYINPUT123), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1285), .A2(new_n1298), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1305), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  OR2_X1    g1134(.A1(new_n1305), .A2(new_n1333), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT123), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1321), .A2(new_n1324), .A3(new_n1336), .A4(new_n1329), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1331), .A2(new_n1334), .A3(new_n1335), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1328), .A2(new_n1338), .ZN(G405));
  AOI21_X1  g1139(.A(new_n1304), .B1(new_n1270), .B2(new_n1301), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT126), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1340), .B(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1270), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(KEYINPUT125), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT125), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1270), .A2(new_n1301), .A3(new_n1345), .A4(new_n1304), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1325), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1342), .A2(new_n1347), .A3(KEYINPUT127), .A4(new_n1348), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1245), .A2(new_n1269), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1300), .A2(G378), .A3(new_n1234), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1303), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1341), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1340), .A2(KEYINPUT126), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1353), .A2(new_n1354), .A3(new_n1344), .A4(new_n1346), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1321), .A2(new_n1324), .A3(KEYINPUT127), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT127), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1325), .A2(new_n1357), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1355), .A2(new_n1356), .A3(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1349), .A2(new_n1359), .ZN(G402));
endmodule


