

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751;

  NAND2_X1 U376 ( .A1(G237), .A2(G234), .ZN(n477) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n468) );
  XNOR2_X1 U378 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n402) );
  XNOR2_X1 U379 ( .A(n511), .B(KEYINPUT75), .ZN(n535) );
  INV_X1 U380 ( .A(n621), .ZN(n496) );
  XNOR2_X1 U381 ( .A(n515), .B(n514), .ZN(n630) );
  AND2_X2 U382 ( .A1(n369), .A2(n391), .ZN(n368) );
  NOR2_X2 U383 ( .A1(n550), .A2(n549), .ZN(n551) );
  AND2_X2 U384 ( .A1(n523), .A2(n603), .ZN(n555) );
  OR2_X2 U385 ( .A1(n590), .A2(KEYINPUT44), .ZN(n353) );
  XNOR2_X2 U386 ( .A(n513), .B(n512), .ZN(n365) );
  NAND2_X2 U387 ( .A1(n368), .A2(n388), .ZN(n367) );
  OR2_X2 U388 ( .A1(n732), .A2(n614), .ZN(n674) );
  NOR2_X1 U389 ( .A1(n602), .A2(n689), .ZN(n587) );
  INV_X1 U390 ( .A(G125), .ZN(n387) );
  NOR2_X1 U391 ( .A1(n716), .A2(G953), .ZN(n717) );
  NAND2_X1 U392 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U393 ( .A(n381), .B(n539), .ZN(n749) );
  XNOR2_X1 U394 ( .A(n577), .B(KEYINPUT33), .ZN(n710) );
  AND2_X1 U395 ( .A1(n603), .A2(n596), .ZN(n577) );
  XNOR2_X1 U396 ( .A(n584), .B(KEYINPUT22), .ZN(n602) );
  NAND2_X1 U397 ( .A1(n689), .A2(n688), .ZN(n694) );
  NAND2_X2 U398 ( .A1(n378), .A2(n377), .ZN(n689) );
  AND2_X1 U399 ( .A1(n380), .A2(n379), .ZN(n378) );
  XNOR2_X1 U400 ( .A(n527), .B(n526), .ZN(n576) );
  AND2_X1 U401 ( .A1(n464), .A2(n432), .ZN(n376) );
  XNOR2_X1 U402 ( .A(n410), .B(n395), .ZN(n495) );
  XNOR2_X1 U403 ( .A(G119), .B(G116), .ZN(n403) );
  XNOR2_X2 U404 ( .A(KEYINPUT64), .B(G953), .ZN(n621) );
  AND2_X4 U405 ( .A1(n617), .A2(n616), .ZN(n718) );
  NAND2_X1 U406 ( .A1(n748), .A2(n607), .ZN(n592) );
  NOR2_X1 U407 ( .A1(n719), .A2(G902), .ZN(n502) );
  XNOR2_X1 U408 ( .A(n466), .B(n465), .ZN(n492) );
  XNOR2_X1 U409 ( .A(n428), .B(G134), .ZN(n466) );
  XNOR2_X2 U410 ( .A(n586), .B(KEYINPUT32), .ZN(n750) );
  XNOR2_X2 U411 ( .A(KEYINPUT67), .B(G101), .ZN(n473) );
  XNOR2_X1 U412 ( .A(n417), .B(KEYINPUT78), .ZN(n418) );
  NAND2_X1 U413 ( .A1(n626), .A2(n374), .ZN(n380) );
  INV_X1 U414 ( .A(n464), .ZN(n374) );
  XNOR2_X1 U415 ( .A(n405), .B(n404), .ZN(n467) );
  XOR2_X1 U416 ( .A(KEYINPUT3), .B(G113), .Z(n404) );
  INV_X1 U417 ( .A(KEYINPUT45), .ZN(n366) );
  XOR2_X1 U418 ( .A(G137), .B(KEYINPUT70), .Z(n491) );
  XNOR2_X1 U419 ( .A(n435), .B(n386), .ZN(n453) );
  INV_X1 U420 ( .A(KEYINPUT10), .ZN(n386) );
  INV_X1 U421 ( .A(G472), .ZN(n360) );
  NAND2_X1 U422 ( .A1(G902), .A2(G472), .ZN(n362) );
  XNOR2_X1 U423 ( .A(G128), .B(G119), .ZN(n448) );
  NAND2_X1 U424 ( .A1(n372), .A2(KEYINPUT2), .ZN(n614) );
  INV_X1 U425 ( .A(KEYINPUT106), .ZN(n384) );
  NAND2_X1 U426 ( .A1(n376), .A2(n375), .ZN(n377) );
  XNOR2_X1 U427 ( .A(n495), .B(n393), .ZN(n392) );
  XNOR2_X1 U428 ( .A(n394), .B(KEYINPUT16), .ZN(n393) );
  INV_X1 U429 ( .A(G122), .ZN(n394) );
  INV_X1 U430 ( .A(G237), .ZN(n401) );
  XNOR2_X1 U431 ( .A(n463), .B(n462), .ZN(n464) );
  AND2_X1 U432 ( .A1(n601), .A2(n609), .ZN(n391) );
  NAND2_X1 U433 ( .A1(n353), .A2(n607), .ZN(n390) );
  NOR2_X1 U434 ( .A1(n576), .A2(n694), .ZN(n596) );
  INV_X1 U435 ( .A(G104), .ZN(n395) );
  NOR2_X1 U436 ( .A1(n682), .A2(n680), .ZN(n447) );
  NOR2_X1 U437 ( .A1(n572), .A2(n571), .ZN(n575) );
  OR2_X1 U438 ( .A1(n618), .A2(n359), .ZN(n358) );
  NAND2_X1 U439 ( .A1(n360), .A2(n432), .ZN(n359) );
  XNOR2_X1 U440 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U441 ( .A(n454), .B(KEYINPUT91), .ZN(n455) );
  XNOR2_X1 U442 ( .A(n429), .B(n466), .ZN(n430) );
  XNOR2_X1 U443 ( .A(n398), .B(n411), .ZN(n397) );
  XNOR2_X1 U444 ( .A(n676), .B(KEYINPUT81), .ZN(n715) );
  NAND2_X1 U445 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X1 U446 ( .A(n579), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n579), .B(KEYINPUT77), .ZN(n354) );
  AND2_X1 U448 ( .A1(n509), .A2(n508), .ZN(n355) );
  XOR2_X1 U449 ( .A(n618), .B(KEYINPUT62), .Z(n356) );
  XOR2_X1 U450 ( .A(KEYINPUT35), .B(KEYINPUT83), .Z(n357) );
  XNOR2_X1 U451 ( .A(n467), .B(n392), .ZN(n735) );
  NAND2_X4 U452 ( .A1(n361), .A2(n358), .ZN(n692) );
  AND2_X1 U453 ( .A1(n363), .A2(n362), .ZN(n361) );
  NAND2_X1 U454 ( .A1(n618), .A2(G472), .ZN(n363) );
  XNOR2_X1 U455 ( .A(n364), .B(n507), .ZN(n508) );
  NAND2_X1 U456 ( .A1(n692), .A2(n678), .ZN(n364) );
  NAND2_X1 U457 ( .A1(n365), .A2(n656), .ZN(n515) );
  NAND2_X1 U458 ( .A1(n365), .A2(n651), .ZN(n625) );
  XNOR2_X2 U459 ( .A(n367), .B(n366), .ZN(n732) );
  NAND2_X1 U460 ( .A1(n593), .A2(KEYINPUT44), .ZN(n369) );
  XNOR2_X2 U461 ( .A(n370), .B(n357), .ZN(n748) );
  NAND2_X1 U462 ( .A1(n371), .A2(n354), .ZN(n370) );
  XNOR2_X1 U463 ( .A(n578), .B(KEYINPUT34), .ZN(n371) );
  INV_X1 U464 ( .A(n373), .ZN(n372) );
  XNOR2_X2 U465 ( .A(n373), .B(KEYINPUT82), .ZN(n672) );
  NAND2_X1 U466 ( .A1(n564), .A2(n563), .ZN(n373) );
  XNOR2_X2 U467 ( .A(n457), .B(n400), .ZN(n626) );
  INV_X1 U468 ( .A(n626), .ZN(n375) );
  OR2_X1 U469 ( .A1(n464), .A2(n432), .ZN(n379) );
  XNOR2_X1 U470 ( .A(n385), .B(n384), .ZN(n383) );
  NAND2_X1 U471 ( .A1(n535), .A2(n559), .ZN(n385) );
  XNOR2_X2 U472 ( .A(n387), .B(G146), .ZN(n435) );
  INV_X1 U473 ( .A(n748), .ZN(n389) );
  XNOR2_X1 U474 ( .A(n396), .B(n735), .ZN(n636) );
  XNOR2_X1 U475 ( .A(n414), .B(n397), .ZN(n396) );
  XNOR2_X1 U476 ( .A(n412), .B(n435), .ZN(n398) );
  NOR2_X2 U477 ( .A1(n572), .A2(n531), .ZN(n657) );
  XNOR2_X1 U478 ( .A(n589), .B(KEYINPUT86), .ZN(n590) );
  AND2_X1 U479 ( .A1(n548), .A2(n547), .ZN(n399) );
  XOR2_X1 U480 ( .A(n452), .B(n451), .Z(n400) );
  XNOR2_X1 U481 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n725) );
  INV_X1 U483 ( .A(n729), .ZN(n622) );
  INV_X1 U484 ( .A(G902), .ZN(n432) );
  NAND2_X1 U485 ( .A1(n432), .A2(n401), .ZN(n416) );
  NAND2_X1 U486 ( .A1(n416), .A2(G214), .ZN(n678) );
  XNOR2_X1 U487 ( .A(n403), .B(n402), .ZN(n405) );
  INV_X1 U488 ( .A(G107), .ZN(n406) );
  NAND2_X1 U489 ( .A1(G110), .A2(n406), .ZN(n409) );
  INV_X1 U490 ( .A(G110), .ZN(n407) );
  NAND2_X1 U491 ( .A1(n407), .A2(G107), .ZN(n408) );
  NAND2_X1 U492 ( .A1(n409), .A2(n408), .ZN(n410) );
  XOR2_X1 U493 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n412) );
  NAND2_X1 U494 ( .A1(G224), .A2(n496), .ZN(n411) );
  XNOR2_X2 U495 ( .A(G143), .B(G128), .ZN(n428) );
  XOR2_X1 U496 ( .A(n428), .B(n473), .Z(n413) );
  XNOR2_X1 U497 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n465) );
  XNOR2_X1 U498 ( .A(n413), .B(n465), .ZN(n414) );
  INV_X1 U499 ( .A(KEYINPUT15), .ZN(n415) );
  XNOR2_X1 U500 ( .A(n415), .B(G902), .ZN(n615) );
  NOR2_X1 U501 ( .A1(n636), .A2(n615), .ZN(n419) );
  NAND2_X1 U502 ( .A1(G210), .A2(n416), .ZN(n417) );
  XNOR2_X1 U503 ( .A(n419), .B(n418), .ZN(n519) );
  BUF_X1 U504 ( .A(n519), .Z(n559) );
  XNOR2_X1 U505 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n420) );
  XNOR2_X1 U506 ( .A(n559), .B(n420), .ZN(n677) );
  NAND2_X1 U507 ( .A1(n678), .A2(n677), .ZN(n682) );
  XOR2_X1 U508 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n422) );
  XNOR2_X1 U509 ( .A(G107), .B(KEYINPUT100), .ZN(n421) );
  XNOR2_X1 U510 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U511 ( .A(n423), .B(KEYINPUT9), .Z(n425) );
  XNOR2_X1 U512 ( .A(G116), .B(G122), .ZN(n424) );
  XNOR2_X1 U513 ( .A(n425), .B(n424), .ZN(n431) );
  NAND2_X1 U514 ( .A1(n496), .A2(G234), .ZN(n427) );
  XNOR2_X1 U515 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n426) );
  XNOR2_X1 U516 ( .A(n427), .B(n426), .ZN(n450) );
  NAND2_X1 U517 ( .A1(n450), .A2(G217), .ZN(n429) );
  NAND2_X1 U518 ( .A1(n725), .A2(n432), .ZN(n434) );
  XOR2_X1 U519 ( .A(KEYINPUT101), .B(G478), .Z(n433) );
  XNOR2_X1 U520 ( .A(n434), .B(n433), .ZN(n536) );
  XNOR2_X1 U521 ( .A(KEYINPUT13), .B(G475), .ZN(n446) );
  XOR2_X1 U522 ( .A(G140), .B(G131), .Z(n493) );
  XNOR2_X1 U523 ( .A(n453), .B(n493), .ZN(n740) );
  XOR2_X1 U524 ( .A(G104), .B(G113), .Z(n437) );
  XNOR2_X1 U525 ( .A(G143), .B(G122), .ZN(n436) );
  XNOR2_X1 U526 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U527 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n439) );
  XNOR2_X1 U528 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n438) );
  XNOR2_X1 U529 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U530 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U531 ( .A1(n468), .A2(G214), .ZN(n442) );
  XNOR2_X1 U532 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U533 ( .A(n740), .B(n444), .ZN(n631) );
  NOR2_X1 U534 ( .A1(G902), .A2(n631), .ZN(n445) );
  XNOR2_X1 U535 ( .A(n446), .B(n445), .ZN(n537) );
  NOR2_X1 U536 ( .A1(n536), .A2(n537), .ZN(n580) );
  INV_X1 U537 ( .A(n580), .ZN(n680) );
  XNOR2_X1 U538 ( .A(n447), .B(KEYINPUT41), .ZN(n709) );
  XOR2_X1 U539 ( .A(G140), .B(G110), .Z(n449) );
  XNOR2_X1 U540 ( .A(n449), .B(n448), .ZN(n452) );
  NAND2_X1 U541 ( .A1(n450), .A2(G221), .ZN(n451) );
  XNOR2_X1 U542 ( .A(n453), .B(KEYINPUT24), .ZN(n456) );
  XNOR2_X1 U543 ( .A(n491), .B(KEYINPUT23), .ZN(n454) );
  INV_X1 U544 ( .A(n615), .ZN(n458) );
  NAND2_X1 U545 ( .A1(n458), .A2(G234), .ZN(n460) );
  XNOR2_X1 U546 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n460), .B(n459), .ZN(n486) );
  AND2_X1 U548 ( .A1(n486), .A2(G217), .ZN(n461) );
  XNOR2_X1 U549 ( .A(n461), .B(KEYINPUT93), .ZN(n463) );
  XNOR2_X1 U550 ( .A(KEYINPUT25), .B(KEYINPUT76), .ZN(n462) );
  XNOR2_X1 U551 ( .A(n492), .B(n467), .ZN(n476) );
  NAND2_X1 U552 ( .A1(n468), .A2(G210), .ZN(n470) );
  XNOR2_X1 U553 ( .A(G137), .B(G131), .ZN(n469) );
  XNOR2_X1 U554 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U555 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n471) );
  XNOR2_X1 U556 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U557 ( .A(n473), .B(G146), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n474), .B(n494), .ZN(n475) );
  XNOR2_X1 U559 ( .A(n476), .B(n475), .ZN(n618) );
  XNOR2_X1 U560 ( .A(n477), .B(KEYINPUT88), .ZN(n478) );
  XNOR2_X1 U561 ( .A(KEYINPUT14), .B(n478), .ZN(n480) );
  NAND2_X1 U562 ( .A1(G952), .A2(n480), .ZN(n707) );
  NOR2_X1 U563 ( .A1(G953), .A2(n707), .ZN(n479) );
  XOR2_X1 U564 ( .A(KEYINPUT89), .B(n479), .Z(n570) );
  INV_X1 U565 ( .A(n570), .ZN(n483) );
  NAND2_X1 U566 ( .A1(G902), .A2(n480), .ZN(n568) );
  NOR2_X1 U567 ( .A1(G900), .A2(n568), .ZN(n481) );
  NAND2_X1 U568 ( .A1(n481), .A2(n621), .ZN(n482) );
  NAND2_X1 U569 ( .A1(n483), .A2(n482), .ZN(n485) );
  INV_X1 U570 ( .A(KEYINPUT79), .ZN(n484) );
  XNOR2_X1 U571 ( .A(n485), .B(n484), .ZN(n509) );
  AND2_X1 U572 ( .A1(n486), .A2(G221), .ZN(n487) );
  XNOR2_X1 U573 ( .A(KEYINPUT21), .B(n487), .ZN(n688) );
  AND2_X1 U574 ( .A1(n509), .A2(n688), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n692), .A2(n520), .ZN(n488) );
  OR2_X1 U576 ( .A1(n689), .A2(n488), .ZN(n490) );
  INV_X1 U577 ( .A(KEYINPUT28), .ZN(n489) );
  XNOR2_X1 U578 ( .A(n490), .B(n489), .ZN(n503) );
  XNOR2_X1 U579 ( .A(n492), .B(n491), .ZN(n741) );
  XNOR2_X1 U580 ( .A(n741), .B(n493), .ZN(n500) );
  XOR2_X1 U581 ( .A(n495), .B(n494), .Z(n498) );
  NAND2_X1 U582 ( .A1(G227), .A2(n496), .ZN(n497) );
  XNOR2_X1 U583 ( .A(n500), .B(n499), .ZN(n719) );
  INV_X1 U584 ( .A(G469), .ZN(n501) );
  XNOR2_X2 U585 ( .A(n502), .B(n501), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n503), .A2(n527), .ZN(n531) );
  OR2_X1 U587 ( .A1(n709), .A2(n531), .ZN(n505) );
  INV_X1 U588 ( .A(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U589 ( .A(n505), .B(n504), .ZN(n751) );
  INV_X1 U590 ( .A(n751), .ZN(n516) );
  INV_X1 U591 ( .A(n694), .ZN(n506) );
  NAND2_X1 U592 ( .A1(n506), .A2(n527), .ZN(n594) );
  INV_X1 U593 ( .A(n594), .ZN(n510) );
  XNOR2_X1 U594 ( .A(KEYINPUT105), .B(KEYINPUT30), .ZN(n507) );
  NAND2_X1 U595 ( .A1(n510), .A2(n355), .ZN(n511) );
  NAND2_X1 U596 ( .A1(n535), .A2(n677), .ZN(n513) );
  XNOR2_X1 U597 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n512) );
  XNOR2_X1 U598 ( .A(n537), .B(KEYINPUT98), .ZN(n541) );
  INV_X1 U599 ( .A(n536), .ZN(n540) );
  AND2_X2 U600 ( .A1(n541), .A2(n540), .ZN(n656) );
  XNOR2_X1 U601 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n514) );
  NAND2_X1 U602 ( .A1(n516), .A2(n630), .ZN(n518) );
  INV_X1 U603 ( .A(KEYINPUT46), .ZN(n517) );
  XNOR2_X1 U604 ( .A(n518), .B(n517), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n519), .A2(n678), .ZN(n530) );
  NAND2_X1 U606 ( .A1(n656), .A2(n520), .ZN(n521) );
  NOR2_X1 U607 ( .A1(n689), .A2(n521), .ZN(n523) );
  INV_X1 U608 ( .A(KEYINPUT6), .ZN(n522) );
  XNOR2_X1 U609 ( .A(n692), .B(n522), .ZN(n603) );
  XNOR2_X1 U610 ( .A(KEYINPUT109), .B(n555), .ZN(n524) );
  NOR2_X1 U611 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U612 ( .A(n525), .B(KEYINPUT36), .ZN(n528) );
  INV_X1 U613 ( .A(KEYINPUT1), .ZN(n526) );
  INV_X1 U614 ( .A(n576), .ZN(n606) );
  NAND2_X1 U615 ( .A1(n528), .A2(n606), .ZN(n669) );
  INV_X1 U616 ( .A(KEYINPUT19), .ZN(n529) );
  XNOR2_X1 U617 ( .A(n530), .B(n529), .ZN(n572) );
  INV_X1 U618 ( .A(KEYINPUT47), .ZN(n532) );
  NOR2_X1 U619 ( .A1(n657), .A2(n532), .ZN(n533) );
  OR2_X1 U620 ( .A1(n533), .A2(KEYINPUT80), .ZN(n534) );
  NAND2_X1 U621 ( .A1(n669), .A2(n534), .ZN(n550) );
  NAND2_X1 U622 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U623 ( .A(n538), .B(KEYINPUT104), .ZN(n579) );
  INV_X1 U624 ( .A(KEYINPUT107), .ZN(n539) );
  NAND2_X1 U625 ( .A1(n657), .A2(KEYINPUT68), .ZN(n545) );
  NAND2_X1 U626 ( .A1(n545), .A2(KEYINPUT80), .ZN(n543) );
  NOR2_X1 U627 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U628 ( .A(n542), .B(KEYINPUT102), .ZN(n651) );
  INV_X1 U629 ( .A(n651), .ZN(n665) );
  INV_X1 U630 ( .A(n656), .ZN(n660) );
  NAND2_X1 U631 ( .A1(n665), .A2(n660), .ZN(n681) );
  NAND2_X1 U632 ( .A1(n543), .A2(n681), .ZN(n544) );
  NAND2_X1 U633 ( .A1(n544), .A2(KEYINPUT47), .ZN(n548) );
  NOR2_X1 U634 ( .A1(KEYINPUT47), .A2(n545), .ZN(n546) );
  NAND2_X1 U635 ( .A1(n546), .A2(n681), .ZN(n547) );
  NAND2_X1 U636 ( .A1(n749), .A2(n399), .ZN(n549) );
  NAND2_X1 U637 ( .A1(n552), .A2(n551), .ZN(n554) );
  INV_X1 U638 ( .A(KEYINPUT48), .ZN(n553) );
  XNOR2_X1 U639 ( .A(n554), .B(n553), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n555), .A2(n678), .ZN(n556) );
  NOR2_X1 U641 ( .A1(n606), .A2(n556), .ZN(n558) );
  INV_X1 U642 ( .A(KEYINPUT43), .ZN(n557) );
  XNOR2_X1 U643 ( .A(n558), .B(n557), .ZN(n561) );
  INV_X1 U644 ( .A(n559), .ZN(n560) );
  AND2_X1 U645 ( .A1(n561), .A2(n560), .ZN(n671) );
  INV_X1 U646 ( .A(n671), .ZN(n562) );
  AND2_X1 U647 ( .A1(n625), .A2(n562), .ZN(n563) );
  XNOR2_X1 U648 ( .A(n672), .B(KEYINPUT74), .ZN(n565) );
  INV_X1 U649 ( .A(n565), .ZN(n611) );
  INV_X1 U650 ( .A(G953), .ZN(n566) );
  NOR2_X1 U651 ( .A1(G898), .A2(n566), .ZN(n567) );
  XOR2_X1 U652 ( .A(KEYINPUT90), .B(n567), .Z(n737) );
  NOR2_X1 U653 ( .A1(n737), .A2(n568), .ZN(n569) );
  NOR2_X1 U654 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U655 ( .A(KEYINPUT0), .B(KEYINPUT66), .Z(n573) );
  XNOR2_X1 U656 ( .A(KEYINPUT87), .B(n573), .ZN(n574) );
  XNOR2_X1 U657 ( .A(n575), .B(n574), .ZN(n582) );
  INV_X1 U658 ( .A(n582), .ZN(n597) );
  NOR2_X1 U659 ( .A1(n597), .A2(n710), .ZN(n578) );
  NAND2_X1 U660 ( .A1(n580), .A2(n688), .ZN(n581) );
  XNOR2_X1 U661 ( .A(KEYINPUT103), .B(n581), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U663 ( .A1(n576), .A2(n603), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n587), .A2(n585), .ZN(n586) );
  NOR2_X1 U665 ( .A1(n606), .A2(n692), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n587), .A2(n588), .ZN(n650) );
  NAND2_X1 U667 ( .A1(n750), .A2(n650), .ZN(n589) );
  INV_X1 U668 ( .A(KEYINPUT85), .ZN(n607) );
  INV_X1 U669 ( .A(n590), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U671 ( .A1(n594), .A2(n692), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n582), .A2(n595), .ZN(n646) );
  NAND2_X1 U673 ( .A1(n692), .A2(n596), .ZN(n698) );
  NOR2_X1 U674 ( .A1(n597), .A2(n698), .ZN(n598) );
  XOR2_X1 U675 ( .A(KEYINPUT31), .B(n598), .Z(n599) );
  XNOR2_X1 U676 ( .A(KEYINPUT95), .B(n599), .ZN(n664) );
  NAND2_X1 U677 ( .A1(n646), .A2(n664), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n600), .A2(n681), .ZN(n601) );
  NOR2_X1 U679 ( .A1(n602), .A2(n603), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n689), .A2(n604), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n642) );
  NOR2_X1 U682 ( .A1(KEYINPUT44), .A2(n607), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n642), .A2(n608), .ZN(n609) );
  INV_X1 U684 ( .A(n732), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n613) );
  INV_X1 U686 ( .A(KEYINPUT2), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n617) );
  AND2_X2 U688 ( .A1(n674), .A2(n615), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n718), .A2(G472), .ZN(n619) );
  XNOR2_X1 U690 ( .A(n619), .B(n356), .ZN(n623) );
  INV_X1 U691 ( .A(G952), .ZN(n620) );
  AND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n729) );
  NAND2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n624), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U695 ( .A(n625), .B(G134), .ZN(G36) );
  NAND2_X1 U696 ( .A1(n718), .A2(G217), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n627), .B(n626), .ZN(n628) );
  NOR2_X2 U698 ( .A1(n628), .A2(n729), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n629), .B(KEYINPUT126), .ZN(G66) );
  XNOR2_X1 U700 ( .A(n630), .B(G131), .ZN(G33) );
  NAND2_X1 U701 ( .A1(n718), .A2(G475), .ZN(n633) );
  XOR2_X1 U702 ( .A(n631), .B(KEYINPUT59), .Z(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(n634) );
  NOR2_X2 U704 ( .A1(n634), .A2(n729), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U706 ( .A1(n718), .A2(G210), .ZN(n639) );
  XOR2_X1 U707 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n637) );
  XNOR2_X1 U708 ( .A(n636), .B(n637), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X2 U710 ( .A1(n640), .A2(n729), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U712 ( .A(G101), .B(n642), .Z(n643) );
  XNOR2_X1 U713 ( .A(KEYINPUT110), .B(n643), .ZN(G3) );
  NOR2_X1 U714 ( .A1(n660), .A2(n646), .ZN(n645) );
  XNOR2_X1 U715 ( .A(G104), .B(KEYINPUT111), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(G6) );
  NOR2_X1 U717 ( .A1(n665), .A2(n646), .ZN(n648) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U720 ( .A(G107), .B(n649), .ZN(G9) );
  XNOR2_X1 U721 ( .A(G110), .B(n650), .ZN(G12) );
  XOR2_X1 U722 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n653) );
  NAND2_X1 U723 ( .A1(n657), .A2(n651), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(n655) );
  XOR2_X1 U725 ( .A(G128), .B(KEYINPUT112), .Z(n654) );
  XNOR2_X1 U726 ( .A(n655), .B(n654), .ZN(G30) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n658), .B(KEYINPUT114), .ZN(n659) );
  XNOR2_X1 U729 ( .A(G146), .B(n659), .ZN(G48) );
  NOR2_X1 U730 ( .A1(n660), .A2(n664), .ZN(n662) );
  XNOR2_X1 U731 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U733 ( .A(G113), .B(n663), .ZN(G15) );
  NOR2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U735 ( .A(G116), .B(KEYINPUT117), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(G18) );
  XOR2_X1 U737 ( .A(KEYINPUT118), .B(KEYINPUT37), .Z(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U739 ( .A(G125), .B(n670), .ZN(G27) );
  XOR2_X1 U740 ( .A(G140), .B(n671), .Z(G42) );
  NOR2_X1 U741 ( .A1(n732), .A2(n672), .ZN(n673) );
  OR2_X1 U742 ( .A1(n673), .A2(KEYINPUT2), .ZN(n675) );
  AND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n685) );
  INV_X1 U746 ( .A(n681), .ZN(n683) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n686), .A2(n710), .ZN(n687) );
  XNOR2_X1 U750 ( .A(n687), .B(KEYINPUT120), .ZN(n703) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n691) );
  XNOR2_X1 U752 ( .A(KEYINPUT49), .B(KEYINPUT119), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n691), .B(n690), .ZN(n693) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U755 ( .A1(n576), .A2(n694), .ZN(n695) );
  XNOR2_X1 U756 ( .A(KEYINPUT50), .B(n695), .ZN(n696) );
  NAND2_X1 U757 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U758 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U759 ( .A(KEYINPUT51), .B(n700), .ZN(n701) );
  NOR2_X1 U760 ( .A1(n709), .A2(n701), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U762 ( .A(n704), .B(KEYINPUT121), .Z(n705) );
  XNOR2_X1 U763 ( .A(KEYINPUT52), .B(n705), .ZN(n706) );
  NOR2_X1 U764 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U765 ( .A(n708), .B(KEYINPUT122), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U767 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U768 ( .A(KEYINPUT123), .B(n713), .Z(n714) );
  NAND2_X1 U769 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U770 ( .A(n717), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U771 ( .A1(n718), .A2(G469), .ZN(n723) );
  XNOR2_X1 U772 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n719), .B(KEYINPUT57), .ZN(n720) );
  XNOR2_X1 U774 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U775 ( .A(n723), .B(n722), .Z(n724) );
  NOR2_X1 U776 ( .A1(n729), .A2(n724), .ZN(G54) );
  NAND2_X1 U777 ( .A1(n718), .A2(G478), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n725), .B(KEYINPUT125), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n729), .A2(n728), .ZN(G63) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U783 ( .A1(n731), .A2(G898), .ZN(n734) );
  OR2_X1 U784 ( .A1(n732), .A2(G953), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n735), .B(G101), .ZN(n736) );
  NAND2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U788 ( .A(n739), .B(n738), .Z(G69) );
  XNOR2_X1 U789 ( .A(n741), .B(n740), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n672), .B(n743), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n742), .A2(n496), .ZN(n747) );
  XNOR2_X1 U792 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U794 ( .A1(G953), .A2(n745), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n747), .A2(n746), .ZN(G72) );
  XOR2_X1 U796 ( .A(G122), .B(n748), .Z(G24) );
  XNOR2_X1 U797 ( .A(G143), .B(n749), .ZN(G45) );
  XNOR2_X1 U798 ( .A(n750), .B(G119), .ZN(G21) );
  XOR2_X1 U799 ( .A(n751), .B(G137), .Z(G39) );
endmodule

