

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U557 ( .A1(n684), .A2(n786), .ZN(n731) );
  NAND2_X1 U558 ( .A1(G8), .A2(n731), .ZN(n770) );
  NOR2_X4 U559 ( .A1(n532), .A2(n531), .ZN(G160) );
  AND2_X2 U560 ( .A1(n528), .A2(G2104), .ZN(n879) );
  NOR2_X1 U561 ( .A1(n731), .A2(n951), .ZN(n700) );
  INV_X1 U562 ( .A(KEYINPUT26), .ZN(n699) );
  NOR2_X1 U563 ( .A1(n990), .A2(n703), .ZN(n705) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n720) );
  XNOR2_X1 U565 ( .A(n721), .B(n720), .ZN(n724) );
  INV_X1 U566 ( .A(KEYINPUT97), .ZN(n725) );
  XNOR2_X1 U567 ( .A(n726), .B(n725), .ZN(n739) );
  NAND2_X1 U568 ( .A1(G160), .A2(G40), .ZN(n785) );
  NOR2_X1 U569 ( .A1(G651), .A2(n621), .ZN(n645) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U571 ( .A1(G113), .A2(n889), .ZN(n526) );
  INV_X1 U572 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U573 ( .A1(G101), .A2(n879), .ZN(n522) );
  XNOR2_X1 U574 ( .A(KEYINPUT23), .B(n522), .ZN(n524) );
  INV_X1 U575 ( .A(KEYINPUT64), .ZN(n523) );
  XNOR2_X1 U576 ( .A(n524), .B(n523), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XOR2_X2 U579 ( .A(KEYINPUT17), .B(n527), .Z(n881) );
  NAND2_X1 U580 ( .A1(G137), .A2(n881), .ZN(n530) );
  NOR2_X1 U581 ( .A1(G2104), .A2(n528), .ZN(n886) );
  NAND2_X1 U582 ( .A1(G125), .A2(n886), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n531) );
  AND2_X1 U584 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U585 ( .A1(G111), .A2(n889), .ZN(n534) );
  NAND2_X1 U586 ( .A1(G135), .A2(n881), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n886), .A2(G123), .ZN(n535) );
  XOR2_X1 U589 ( .A(KEYINPUT18), .B(n535), .Z(n536) );
  NOR2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n879), .A2(G99), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n928) );
  XNOR2_X1 U593 ( .A(G2096), .B(n928), .ZN(n540) );
  OR2_X1 U594 ( .A1(G2100), .A2(n540), .ZN(G156) );
  INV_X1 U595 ( .A(G57), .ZN(G237) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U599 ( .A1(G90), .A2(n639), .ZN(n543) );
  XNOR2_X1 U600 ( .A(G543), .B(KEYINPUT0), .ZN(n541) );
  XNOR2_X1 U601 ( .A(n541), .B(KEYINPUT65), .ZN(n621) );
  INV_X1 U602 ( .A(G651), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n621), .A2(n545), .ZN(n640) );
  NAND2_X1 U604 ( .A1(G77), .A2(n640), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n544), .B(KEYINPUT9), .ZN(n548) );
  NOR2_X1 U607 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT1), .B(n546), .Z(n638) );
  NAND2_X1 U609 ( .A1(G64), .A2(n638), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n645), .A2(G52), .ZN(n549) );
  XOR2_X1 U612 ( .A(KEYINPUT66), .B(n549), .Z(n550) );
  NOR2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT67), .B(n552), .Z(G171) );
  NAND2_X1 U615 ( .A1(n639), .A2(G89), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U617 ( .A1(G76), .A2(n640), .ZN(n554) );
  NAND2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U619 ( .A(n556), .B(KEYINPUT5), .ZN(n563) );
  XNOR2_X1 U620 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n645), .A2(G51), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(KEYINPUT74), .ZN(n559) );
  NAND2_X1 U623 ( .A1(G63), .A2(n638), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U627 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(n565) );
  XNOR2_X1 U629 ( .A(KEYINPUT76), .B(n565), .ZN(G286) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U632 ( .A(G223), .ZN(n826) );
  NAND2_X1 U633 ( .A1(n826), .A2(G567), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U635 ( .A1(G56), .A2(n638), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n568), .Z(n575) );
  NAND2_X1 U637 ( .A1(G81), .A2(n639), .ZN(n569) );
  XOR2_X1 U638 ( .A(KEYINPUT12), .B(n569), .Z(n570) );
  XNOR2_X1 U639 ( .A(n570), .B(KEYINPUT71), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G68), .A2(n640), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U642 ( .A(KEYINPUT13), .B(n573), .Z(n574) );
  NOR2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n645), .A2(G43), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n990) );
  INV_X1 U646 ( .A(G860), .ZN(n599) );
  OR2_X1 U647 ( .A1(n990), .A2(n599), .ZN(G153) );
  XOR2_X1 U648 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G54), .A2(n645), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G66), .A2(n638), .ZN(n579) );
  NAND2_X1 U652 ( .A1(G92), .A2(n639), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G79), .A2(n640), .ZN(n580) );
  XNOR2_X1 U655 ( .A(KEYINPUT73), .B(n580), .ZN(n581) );
  NOR2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT15), .ZN(n975) );
  OR2_X1 U659 ( .A1(n975), .A2(G868), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G53), .A2(n645), .ZN(n588) );
  XOR2_X1 U662 ( .A(KEYINPUT70), .B(n588), .Z(n594) );
  NAND2_X1 U663 ( .A1(n640), .A2(G78), .ZN(n589) );
  XNOR2_X1 U664 ( .A(n589), .B(KEYINPUT68), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G91), .A2(n639), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U667 ( .A(KEYINPUT69), .B(n592), .Z(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n638), .A2(G65), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(G299) );
  NAND2_X1 U671 ( .A1(G868), .A2(G286), .ZN(n598) );
  INV_X1 U672 ( .A(G868), .ZN(n657) );
  NAND2_X1 U673 ( .A1(G299), .A2(n657), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n600), .A2(n975), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT77), .ZN(n602) );
  XOR2_X1 U678 ( .A(KEYINPUT16), .B(n602), .Z(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n990), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G868), .A2(n975), .ZN(n603) );
  NOR2_X1 U681 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G559), .A2(n975), .ZN(n606) );
  XOR2_X1 U684 ( .A(n990), .B(n606), .Z(n655) );
  XOR2_X1 U685 ( .A(n655), .B(KEYINPUT78), .Z(n607) );
  NOR2_X1 U686 ( .A1(G860), .A2(n607), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G93), .A2(n639), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G80), .A2(n640), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U690 ( .A1(G67), .A2(n638), .ZN(n610) );
  XNOR2_X1 U691 ( .A(KEYINPUT79), .B(n610), .ZN(n611) );
  NOR2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n645), .A2(G55), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n658) );
  XOR2_X1 U695 ( .A(n615), .B(n658), .Z(G145) );
  NAND2_X1 U696 ( .A1(n645), .A2(G49), .ZN(n616) );
  XNOR2_X1 U697 ( .A(n616), .B(KEYINPUT80), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U700 ( .A(KEYINPUT81), .B(n619), .Z(n620) );
  NOR2_X1 U701 ( .A1(n638), .A2(n620), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n621), .A2(G87), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(G288) );
  NAND2_X1 U704 ( .A1(G88), .A2(n639), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G75), .A2(n640), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G62), .A2(n638), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G50), .A2(n645), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(G166) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n631) );
  NAND2_X1 U712 ( .A1(G73), .A2(n640), .ZN(n630) );
  XNOR2_X1 U713 ( .A(n631), .B(n630), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G61), .A2(n638), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G86), .A2(n639), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n645), .A2(G48), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(G305) );
  AND2_X1 U720 ( .A1(n638), .A2(G60), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G85), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G72), .A2(n640), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n645), .A2(G47), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(G290) );
  INV_X1 U727 ( .A(G299), .ZN(n715) );
  XNOR2_X1 U728 ( .A(n715), .B(G288), .ZN(n654) );
  XNOR2_X1 U729 ( .A(G166), .B(n658), .ZN(n651) );
  XNOR2_X1 U730 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n649) );
  XNOR2_X1 U731 ( .A(G305), .B(KEYINPUT84), .ZN(n648) );
  XNOR2_X1 U732 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U733 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n652), .B(G290), .ZN(n653) );
  XNOR2_X1 U735 ( .A(n654), .B(n653), .ZN(n902) );
  XOR2_X1 U736 ( .A(n902), .B(n655), .Z(n656) );
  NOR2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n660) );
  NOR2_X1 U738 ( .A1(G868), .A2(n658), .ZN(n659) );
  NOR2_X1 U739 ( .A1(n660), .A2(n659), .ZN(G295) );
  XOR2_X1 U740 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n664) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U743 ( .A1(n662), .A2(G2090), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U745 ( .A1(G2072), .A2(n665), .ZN(G158) );
  XNOR2_X1 U746 ( .A(KEYINPUT86), .B(G44), .ZN(n666) );
  XNOR2_X1 U747 ( .A(n666), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U748 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U751 ( .A1(G218), .A2(n668), .ZN(n669) );
  XOR2_X1 U752 ( .A(KEYINPUT87), .B(n669), .Z(n670) );
  NAND2_X1 U753 ( .A1(G96), .A2(n670), .ZN(n832) );
  NAND2_X1 U754 ( .A1(n832), .A2(G2106), .ZN(n674) );
  NAND2_X1 U755 ( .A1(G69), .A2(G120), .ZN(n671) );
  NOR2_X1 U756 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U757 ( .A1(G108), .A2(n672), .ZN(n833) );
  NAND2_X1 U758 ( .A1(n833), .A2(G567), .ZN(n673) );
  NAND2_X1 U759 ( .A1(n674), .A2(n673), .ZN(n834) );
  NOR2_X1 U760 ( .A1(n675), .A2(n834), .ZN(n676) );
  XNOR2_X1 U761 ( .A(n676), .B(KEYINPUT88), .ZN(n830) );
  NAND2_X1 U762 ( .A1(G36), .A2(n830), .ZN(G176) );
  NAND2_X1 U763 ( .A1(G138), .A2(n881), .ZN(n678) );
  NAND2_X1 U764 ( .A1(G102), .A2(n879), .ZN(n677) );
  NAND2_X1 U765 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U766 ( .A1(G114), .A2(n889), .ZN(n680) );
  NAND2_X1 U767 ( .A1(G126), .A2(n886), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U769 ( .A1(n682), .A2(n681), .ZN(G164) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n754) );
  INV_X1 U772 ( .A(KEYINPUT94), .ZN(n683) );
  XNOR2_X1 U773 ( .A(n683), .B(n785), .ZN(n684) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n786) );
  NOR2_X1 U775 ( .A1(G2084), .A2(n731), .ZN(n687) );
  NAND2_X1 U776 ( .A1(G8), .A2(n687), .ZN(n730) );
  NOR2_X1 U777 ( .A1(G1966), .A2(n770), .ZN(n728) );
  INV_X1 U778 ( .A(n731), .ZN(n706) );
  OR2_X1 U779 ( .A1(n706), .A2(G1961), .ZN(n686) );
  XNOR2_X1 U780 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U781 ( .A1(n706), .A2(n955), .ZN(n685) );
  NAND2_X1 U782 ( .A1(n686), .A2(n685), .ZN(n722) );
  NOR2_X1 U783 ( .A1(G171), .A2(n722), .ZN(n692) );
  NOR2_X1 U784 ( .A1(n728), .A2(n687), .ZN(n688) );
  NAND2_X1 U785 ( .A1(G8), .A2(n688), .ZN(n689) );
  XNOR2_X1 U786 ( .A(KEYINPUT30), .B(n689), .ZN(n690) );
  NOR2_X1 U787 ( .A1(G168), .A2(n690), .ZN(n691) );
  NOR2_X1 U788 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U789 ( .A(n693), .B(KEYINPUT31), .Z(n694) );
  XNOR2_X1 U790 ( .A(KEYINPUT98), .B(n694), .ZN(n737) );
  NAND2_X1 U791 ( .A1(n706), .A2(G2072), .ZN(n695) );
  XNOR2_X1 U792 ( .A(n695), .B(KEYINPUT27), .ZN(n697) );
  INV_X1 U793 ( .A(G1956), .ZN(n1001) );
  NOR2_X1 U794 ( .A1(n1001), .A2(n706), .ZN(n696) );
  NOR2_X1 U795 ( .A1(n697), .A2(n696), .ZN(n714) );
  NOR2_X1 U796 ( .A1(n715), .A2(n714), .ZN(n698) );
  XOR2_X1 U797 ( .A(n698), .B(KEYINPUT28), .Z(n719) );
  INV_X1 U798 ( .A(G1996), .ZN(n951) );
  XNOR2_X1 U799 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n731), .A2(G1341), .ZN(n701) );
  NAND2_X1 U801 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U802 ( .A1(n705), .A2(n975), .ZN(n704) );
  XOR2_X1 U803 ( .A(n704), .B(KEYINPUT96), .Z(n713) );
  NAND2_X1 U804 ( .A1(n705), .A2(n975), .ZN(n711) );
  AND2_X1 U805 ( .A1(n706), .A2(G2067), .ZN(n707) );
  XNOR2_X1 U806 ( .A(n707), .B(KEYINPUT95), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n731), .A2(G1348), .ZN(n708) );
  NAND2_X1 U808 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U814 ( .A1(G171), .A2(n722), .ZN(n723) );
  NAND2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n726) );
  AND2_X1 U816 ( .A1(n737), .A2(n739), .ZN(n727) );
  NOR2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n746) );
  INV_X1 U819 ( .A(G8), .ZN(n736) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n770), .ZN(n733) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n731), .ZN(n732) );
  NOR2_X1 U822 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n734), .A2(G303), .ZN(n735) );
  OR2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n740) );
  AND2_X1 U825 ( .A1(n737), .A2(n740), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n743) );
  INV_X1 U827 ( .A(n740), .ZN(n741) );
  OR2_X1 U828 ( .A1(n741), .A2(G286), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U830 ( .A(n744), .B(KEYINPUT32), .ZN(n745) );
  NAND2_X1 U831 ( .A1(n746), .A2(n745), .ZN(n766) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n747) );
  XNOR2_X1 U833 ( .A(KEYINPUT99), .B(n747), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n766), .A2(n748), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n754), .A2(n749), .ZN(n752) );
  AND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NOR2_X1 U837 ( .A1(n979), .A2(n770), .ZN(n750) );
  NAND2_X1 U838 ( .A1(KEYINPUT100), .A2(n750), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U840 ( .A1(n753), .A2(KEYINPUT33), .ZN(n758) );
  INV_X1 U841 ( .A(n754), .ZN(n982) );
  NOR2_X1 U842 ( .A1(n770), .A2(n982), .ZN(n760) );
  INV_X1 U843 ( .A(n760), .ZN(n756) );
  NAND2_X1 U844 ( .A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n763) );
  OR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n768) );
  NAND2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n768), .A2(n759), .ZN(n992) );
  NOR2_X1 U850 ( .A1(KEYINPUT100), .A2(n760), .ZN(n761) );
  NOR2_X1 U851 ( .A1(n992), .A2(n761), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n774) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n764) );
  NAND2_X1 U854 ( .A1(G8), .A2(n764), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  AND2_X1 U856 ( .A1(n767), .A2(n770), .ZN(n772) );
  XNOR2_X1 U857 ( .A(n768), .B(KEYINPUT24), .ZN(n769) );
  NOR2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  AND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n807) );
  NAND2_X1 U861 ( .A1(G140), .A2(n881), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G104), .A2(n879), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n778) );
  XOR2_X1 U864 ( .A(KEYINPUT34), .B(KEYINPUT89), .Z(n777) );
  XNOR2_X1 U865 ( .A(n778), .B(n777), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G116), .A2(n889), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G128), .A2(n886), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U869 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n784), .ZN(n873) );
  XNOR2_X1 U872 ( .A(KEYINPUT37), .B(G2067), .ZN(n819) );
  NOR2_X1 U873 ( .A1(n873), .A2(n819), .ZN(n931) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n821) );
  NAND2_X1 U875 ( .A1(n931), .A2(n821), .ZN(n817) );
  XNOR2_X1 U876 ( .A(KEYINPUT91), .B(G1991), .ZN(n956) );
  NAND2_X1 U877 ( .A1(G119), .A2(n886), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G95), .A2(n879), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n881), .A2(G131), .ZN(n789) );
  XOR2_X1 U881 ( .A(KEYINPUT90), .B(n789), .Z(n790) );
  NOR2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n889), .A2(G107), .ZN(n792) );
  AND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n893) );
  OR2_X1 U885 ( .A1(n956), .A2(n893), .ZN(n803) );
  NAND2_X1 U886 ( .A1(G117), .A2(n889), .ZN(n795) );
  NAND2_X1 U887 ( .A1(G129), .A2(n886), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n879), .A2(G105), .ZN(n796) );
  XOR2_X1 U890 ( .A(KEYINPUT38), .B(n796), .Z(n797) );
  NOR2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U892 ( .A(n799), .B(KEYINPUT92), .ZN(n801) );
  NAND2_X1 U893 ( .A1(G141), .A2(n881), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n894) );
  NAND2_X1 U895 ( .A1(G1996), .A2(n894), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n924) );
  NAND2_X1 U897 ( .A1(n924), .A2(n821), .ZN(n804) );
  XNOR2_X1 U898 ( .A(n804), .B(KEYINPUT93), .ZN(n813) );
  INV_X1 U899 ( .A(n813), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n817), .A2(n805), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n809) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U903 ( .A1(n978), .A2(n821), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n824) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n894), .ZN(n939) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n893), .A2(n956), .ZN(n810) );
  XNOR2_X1 U908 ( .A(n810), .B(KEYINPUT101), .ZN(n927) );
  NOR2_X1 U909 ( .A1(n811), .A2(n927), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U911 ( .A(n814), .B(KEYINPUT102), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n939), .A2(n815), .ZN(n816) );
  XNOR2_X1 U913 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n873), .A2(n819), .ZN(n923) );
  NAND2_X1 U916 ( .A1(n820), .A2(n923), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n826), .ZN(G217) );
  NAND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n827) );
  XOR2_X1 U922 ( .A(KEYINPUT104), .B(n827), .Z(n828) );
  NAND2_X1 U923 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U926 ( .A(KEYINPUT105), .B(n831), .Z(G188) );
  NOR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G325) );
  XOR2_X1 U928 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  INV_X1 U933 ( .A(n834), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT42), .B(G2090), .Z(n836) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2084), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U937 ( .A(n837), .B(G2100), .Z(n839) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2072), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(G2096), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U941 ( .A(KEYINPUT107), .B(G2678), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n843), .B(n842), .Z(G227) );
  XOR2_X1 U944 ( .A(G1976), .B(G1956), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1991), .B(G1996), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n855) );
  XOR2_X1 U947 ( .A(KEYINPUT108), .B(KEYINPUT110), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1981), .B(G2474), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U950 ( .A(G1971), .B(G1961), .Z(n849) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1966), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G124), .A2(n886), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n889), .A2(G112), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G136), .A2(n881), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G100), .A2(n879), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U964 ( .A1(n862), .A2(n861), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G139), .A2(n881), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G103), .A2(n879), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n886), .A2(G127), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n865), .B(KEYINPUT114), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G115), .A2(n889), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U972 ( .A(KEYINPUT47), .B(n868), .ZN(n869) );
  XNOR2_X1 U973 ( .A(KEYINPUT115), .B(n869), .ZN(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(KEYINPUT116), .B(n872), .Z(n934) );
  XNOR2_X1 U976 ( .A(G160), .B(n873), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(n928), .ZN(n878) );
  XOR2_X1 U978 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n876) );
  XNOR2_X1 U979 ( .A(G164), .B(KEYINPUT46), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U981 ( .A(n878), .B(n877), .Z(n899) );
  NAND2_X1 U982 ( .A1(n879), .A2(G106), .ZN(n880) );
  XNOR2_X1 U983 ( .A(KEYINPUT112), .B(n880), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n881), .A2(G142), .ZN(n882) );
  XOR2_X1 U985 ( .A(KEYINPUT113), .B(n882), .Z(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n885), .B(KEYINPUT45), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G130), .A2(n886), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U990 ( .A1(G118), .A2(n889), .ZN(n890) );
  XNOR2_X1 U991 ( .A(KEYINPUT111), .B(n890), .ZN(n891) );
  NOR2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n897) );
  XOR2_X1 U993 ( .A(G162), .B(n893), .Z(n895) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(n934), .B(n900), .Z(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U999 ( .A(n990), .B(n902), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(G171), .B(n975), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1002 ( .A(n905), .B(G286), .Z(n906) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U1004 ( .A(G2454), .B(G2435), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G2438), .B(G2427), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n915) );
  XOR2_X1 U1007 ( .A(KEYINPUT103), .B(G2446), .Z(n910) );
  XNOR2_X1 U1008 ( .A(G2443), .B(G2430), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1010 ( .A(n911), .B(G2451), .Z(n913) );
  XNOR2_X1 U1011 ( .A(G1348), .B(G1341), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n916), .A2(G14), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  INV_X1 U1023 ( .A(n922), .ZN(G401) );
  INV_X1 U1024 ( .A(n923), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n933) );
  XOR2_X1 U1026 ( .A(G2084), .B(G160), .Z(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n944) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n936) );
  XNOR2_X1 U1032 ( .A(G2072), .B(n934), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(KEYINPUT50), .B(n937), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n940), .Z(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1040 ( .A(KEYINPUT52), .B(n945), .Z(n946) );
  NOR2_X1 U1041 ( .A1(KEYINPUT55), .A2(n946), .ZN(n948) );
  INV_X1 U1042 ( .A(G29), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n1031) );
  XNOR2_X1 U1044 ( .A(G29), .B(KEYINPUT121), .ZN(n972) );
  XOR2_X1 U1045 ( .A(KEYINPUT119), .B(G34), .Z(n950) );
  XNOR2_X1 U1046 ( .A(G2084), .B(KEYINPUT54), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n950), .B(n949), .ZN(n968) );
  XOR2_X1 U1048 ( .A(G2090), .B(G35), .Z(n966) );
  XNOR2_X1 U1049 ( .A(G32), .B(n951), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n952), .A2(G28), .ZN(n962) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1054 ( .A(n955), .B(G27), .Z(n958) );
  XOR2_X1 U1055 ( .A(n956), .B(G25), .Z(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1059 ( .A(KEYINPUT53), .B(n963), .Z(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(KEYINPUT118), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n970), .B(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(G11), .ZN(n1028) );
  INV_X1 U1067 ( .A(G16), .ZN(n1024) );
  XOR2_X1 U1068 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n974) );
  XNOR2_X1 U1069 ( .A(n1024), .B(n974), .ZN(n1000) );
  XOR2_X1 U1070 ( .A(G1348), .B(n975), .Z(n977) );
  XNOR2_X1 U1071 ( .A(G303), .B(G1971), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1075 ( .A(KEYINPUT124), .B(n982), .Z(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n988) );
  XOR2_X1 U1077 ( .A(G171), .B(G1961), .Z(n986) );
  XNOR2_X1 U1078 ( .A(G299), .B(G1956), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(n989), .ZN(n998) );
  XNOR2_X1 U1082 ( .A(n990), .B(G1341), .ZN(n996) );
  XOR2_X1 U1083 ( .A(G168), .B(G1966), .Z(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1085 ( .A(KEYINPUT57), .B(n993), .Z(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT123), .B(n994), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  XNOR2_X1 U1090 ( .A(G20), .B(n1001), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(KEYINPUT59), .B(G1348), .Z(n1006) );
  XNOR2_X1 U1096 ( .A(G4), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1009), .ZN(n1019) );
  XNOR2_X1 U1099 ( .A(G1961), .B(KEYINPUT126), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(G5), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(G21), .B(G1966), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1115 ( .A(n1029), .B(KEYINPUT127), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1032), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

