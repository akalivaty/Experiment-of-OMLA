//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936;
  XOR2_X1   g000(.A(KEYINPUT72), .B(KEYINPUT73), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G43gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT28), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n210));
  OR2_X1    g009(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212));
  NAND2_X1  g011(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI211_X1 g013(.A(new_n208), .B(G190gat), .C1(new_n210), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n218));
  OR2_X1    g017(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n207), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n210), .A2(new_n214), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT28), .A3(new_n216), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(KEYINPUT68), .A3(new_n220), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT69), .ZN(new_n232));
  INV_X1    g031(.A(new_n229), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(KEYINPUT26), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n222), .A2(new_n224), .A3(new_n227), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G183gat), .B2(G190gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND3_X1   g039(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n229), .B(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n236), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n239), .B(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n236), .B(new_n244), .C1(new_n247), .C2(new_n238), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(KEYINPUT65), .B2(new_n236), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n245), .B1(new_n249), .B2(new_n228), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G120gat), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n253));
  INV_X1    g052(.A(G127gat), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n254), .A2(G134gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(G134gat), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT70), .B(G134gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G127gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n255), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(KEYINPUT71), .A3(G127gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n257), .B1(new_n263), .B2(new_n253), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n251), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n253), .ZN(new_n266));
  INV_X1    g065(.A(new_n257), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n235), .A2(new_n250), .A3(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n265), .A2(G227gat), .A3(G233gat), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT33), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n206), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(KEYINPUT32), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n270), .B(KEYINPUT32), .C1(new_n271), .C2(new_n206), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n269), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n268), .B1(new_n235), .B2(new_n250), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n269), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n277), .B1(new_n283), .B2(new_n278), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT76), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n276), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT31), .B(G50gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(G106gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G22gat), .B(G78gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT86), .ZN(new_n297));
  OR2_X1    g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT81), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT82), .B(G155gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G162gat), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n301), .A2(new_n303), .B1(new_n305), .B2(KEYINPUT2), .ZN(new_n306));
  XNOR2_X1  g105(.A(G141gat), .B(G148gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT80), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n307), .A2(KEYINPUT2), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n300), .ZN(new_n311));
  INV_X1    g110(.A(new_n300), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n312), .B(KEYINPUT80), .C1(KEYINPUT2), .C2(new_n307), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n306), .A2(new_n308), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT77), .B(KEYINPUT22), .Z(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n325), .ZN(new_n327));
  INV_X1    g126(.A(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n297), .B1(new_n316), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n313), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n301), .A2(new_n303), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n308), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n322), .A2(new_n323), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n324), .A2(new_n337), .A3(KEYINPUT29), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n338), .B2(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(new_n315), .A3(new_n335), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n329), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(KEYINPUT86), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n331), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G228gat), .A2(G233gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n346), .B(KEYINPUT85), .Z(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT87), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n346), .B1(new_n342), .B2(new_n343), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT3), .B1(new_n330), .B2(new_n341), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(new_n314), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n296), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n345), .A2(new_n350), .A3(new_n347), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n350), .B1(new_n345), .B2(new_n347), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n296), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n294), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n295), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(new_n293), .A3(new_n359), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n274), .A2(new_n285), .A3(new_n275), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT75), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n274), .A2(new_n285), .A3(new_n368), .A4(new_n275), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n291), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  INV_X1    g171(.A(G64gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G92gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G226gat), .ZN(new_n377));
  INV_X1    g176(.A(G233gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n235), .A2(new_n250), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n235), .B2(new_n250), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n379), .A2(KEYINPUT29), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n251), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n343), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n383), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(new_n381), .A3(new_n385), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n251), .A2(new_n377), .A3(new_n378), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n343), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n376), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n389), .A2(new_n381), .A3(new_n385), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n330), .B1(new_n395), .B2(new_n391), .ZN(new_n396));
  INV_X1    g195(.A(new_n376), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n387), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n398), .A3(KEYINPUT30), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n396), .A2(new_n387), .A3(new_n400), .A4(new_n397), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(new_n268), .A3(new_n340), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n264), .A2(new_n314), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n264), .B2(new_n314), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n403), .B(new_n405), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n403), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n264), .A2(new_n314), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n264), .A2(new_n314), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n410), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n417), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT89), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n264), .B1(KEYINPUT3), .B2(new_n336), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n428), .A2(new_n407), .B1(new_n429), .B2(new_n340), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT5), .B1(new_n430), .B2(new_n403), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n424), .B1(new_n410), .B2(new_n415), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n423), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT84), .B(KEYINPUT6), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n425), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(new_n422), .ZN(new_n439));
  INV_X1    g238(.A(new_n426), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n436), .A2(new_n439), .B1(new_n440), .B2(new_n437), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n402), .A2(new_n441), .A3(KEYINPUT35), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n371), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n437), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n433), .B2(new_n423), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(new_n440), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n287), .A2(new_n366), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n399), .A2(new_n401), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n365), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(KEYINPUT36), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(KEYINPUT74), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT74), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n288), .A2(new_n290), .B1(new_n367), .B2(new_n369), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(KEYINPUT36), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  INV_X1    g256(.A(new_n398), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT37), .B1(new_n388), .B2(new_n393), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n396), .A2(new_n387), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n461), .A3(new_n376), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n458), .B1(new_n462), .B2(KEYINPUT38), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n343), .B1(new_n395), .B2(new_n391), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n384), .A2(new_n330), .A3(new_n386), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(KEYINPUT37), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n461), .A3(new_n467), .A4(new_n376), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n441), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n430), .A2(KEYINPUT88), .A3(new_n403), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n411), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT88), .B1(new_n430), .B2(new_n403), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n472), .A3(new_n411), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n413), .A2(new_n414), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n470), .B1(new_n478), .B2(new_n403), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n480), .A3(KEYINPUT40), .A4(new_n422), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n434), .B1(new_n433), .B2(new_n423), .ZN(new_n482));
  NOR4_X1   g281(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT89), .A4(new_n422), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n476), .A2(new_n477), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n423), .B1(new_n485), .B2(new_n470), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT40), .B1(new_n486), .B2(new_n480), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n402), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n489), .A3(new_n365), .ZN(new_n490));
  INV_X1    g289(.A(new_n365), .ZN(new_n491));
  INV_X1    g290(.A(new_n446), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n402), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n451), .B1(new_n457), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT92), .B(G29gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT14), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n498), .A2(G29gat), .A3(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504));
  INV_X1    g303(.A(G43gat), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT93), .B1(new_n505), .B2(G50gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n503), .B(new_n504), .C1(new_n507), .C2(new_n501), .ZN(new_n508));
  OR3_X1    g307(.A1(new_n501), .A2(new_n507), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT17), .ZN(new_n511));
  XOR2_X1   g310(.A(G99gat), .B(G106gat), .Z(new_n512));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT8), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(G85gat), .B2(G92gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(KEYINPUT98), .ZN(new_n517));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT98), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n518), .B(KEYINPUT99), .C1(new_n519), .C2(KEYINPUT7), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(KEYINPUT98), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT99), .B1(new_n522), .B2(new_n518), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n517), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n519), .B2(KEYINPUT7), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT99), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n517), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(new_n520), .ZN(new_n529));
  AOI211_X1 g328(.A(new_n512), .B(new_n515), .C1(new_n524), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n512), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n529), .ZN(new_n532));
  INV_X1    g331(.A(new_n515), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n511), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n531), .A3(new_n533), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n521), .A2(new_n523), .A3(new_n517), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n528), .B1(new_n527), .B2(new_n520), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n512), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n510), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT100), .B(G190gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G218gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n543), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT97), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT101), .ZN(new_n549));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(KEYINPUT97), .A3(new_n551), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  OR2_X1    g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G57gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(G64gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT95), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n560), .B2(G64gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n373), .A2(G57gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT9), .B1(new_n566), .B2(new_n561), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n556), .A3(new_n557), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n254), .ZN(new_n573));
  XOR2_X1   g372(.A(G15gat), .B(G22gat), .Z(new_n574));
  INV_X1    g373(.A(G1gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n577));
  AOI21_X1  g376(.A(G8gat), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT16), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(G1gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n576), .B1(new_n580), .B2(new_n574), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n578), .B(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n571), .B2(new_n570), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n573), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT96), .B(G155gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n588), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n555), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n511), .A2(new_n582), .ZN(new_n595));
  INV_X1    g394(.A(new_n510), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n596), .A2(new_n582), .ZN(new_n597));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT18), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n510), .B(new_n582), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n598), .B(KEYINPUT13), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n595), .A2(KEYINPUT18), .A3(new_n597), .A4(new_n598), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT91), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT90), .B(G197gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT11), .B(G169gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618));
  INV_X1    g417(.A(G176gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n620), .B(G204gat), .Z(new_n621));
  OAI21_X1  g420(.A(new_n570), .B1(new_n534), .B2(new_n530), .ZN(new_n622));
  INV_X1    g421(.A(new_n570), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n540), .A2(new_n623), .A3(new_n536), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n540), .A2(new_n536), .A3(KEYINPUT10), .A4(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n629), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n626), .B2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n629), .B1(new_n622), .B2(new_n624), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n621), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n634), .A2(new_n637), .A3(new_n621), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n617), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n495), .A2(new_n594), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n492), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g445(.A1(new_n644), .A2(new_n402), .ZN(new_n647));
  INV_X1    g446(.A(G8gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n579), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n647), .A2(new_n648), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n651), .A2(KEYINPUT103), .A3(new_n652), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT103), .B1(new_n651), .B2(new_n652), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n653), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n644), .B2(new_n455), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n457), .A2(G15gat), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n644), .B2(new_n659), .ZN(G1326gat));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n491), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  NAND2_X1  g464(.A1(new_n495), .A2(new_n555), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n643), .A2(new_n593), .ZN(new_n667));
  NOR4_X1   g466(.A1(new_n666), .A2(new_n446), .A3(new_n496), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n495), .B(new_n555), .C1(KEYINPUT107), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n371), .A2(new_n442), .B1(new_n449), .B2(KEYINPUT35), .ZN(new_n675));
  INV_X1    g474(.A(new_n452), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n454), .ZN(new_n677));
  INV_X1    g476(.A(new_n290), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n289), .B1(new_n276), .B2(new_n286), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n370), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT36), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT74), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n677), .B1(new_n682), .B2(new_n676), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n365), .B1(new_n446), .B2(new_n448), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n439), .B1(new_n482), .B2(new_n483), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n440), .A2(new_n437), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n685), .A2(new_n468), .A3(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n687), .A2(new_n463), .B1(new_n488), .B2(new_n402), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n684), .B1(new_n688), .B2(new_n365), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n675), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n555), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n674), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n672), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n667), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n496), .B1(new_n695), .B2(new_n446), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n670), .A2(new_n696), .ZN(G1328gat));
  OAI21_X1  g496(.A(G36gat), .B1(new_n695), .B2(new_n448), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n666), .A2(G36gat), .A3(new_n448), .A4(new_n667), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n700), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n701), .B2(new_n703), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n698), .B1(new_n704), .B2(new_n705), .ZN(G1329gat));
  NOR2_X1   g505(.A1(new_n666), .A2(new_n667), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n505), .A3(new_n455), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n695), .A2(new_n683), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(new_n505), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT47), .B1(new_n708), .B2(KEYINPUT109), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI221_X1 g511(.A(new_n708), .B1(KEYINPUT109), .B2(KEYINPUT47), .C1(new_n709), .C2(new_n505), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1330gat));
  NAND2_X1  g513(.A1(new_n491), .A2(G50gat), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n666), .A2(new_n365), .A3(new_n667), .ZN(new_n716));
  OAI22_X1  g515(.A1(new_n695), .A2(new_n715), .B1(G50gat), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g517(.A1(new_n594), .A2(new_n642), .A3(new_n617), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT110), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n495), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n446), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(new_n560), .ZN(G1332gat));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n448), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n721), .B2(new_n683), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n721), .A2(G71gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n680), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g531(.A1(new_n721), .A2(new_n365), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT111), .B(G78gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n616), .A2(new_n592), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n642), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT112), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n672), .B2(new_n692), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n446), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n641), .A2(G85gat), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n495), .A2(new_n555), .A3(new_n736), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n745), .A2(new_n746), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(KEYINPUT113), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n743), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n742), .B1(new_n752), .B2(new_n446), .ZN(G1336gat));
  NOR3_X1   g552(.A1(new_n448), .A2(G92gat), .A3(new_n641), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n749), .B2(new_n751), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n671), .A2(KEYINPUT107), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n690), .A2(new_n691), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n673), .B1(new_n495), .B2(new_n555), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n402), .B(new_n738), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n755), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n746), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n754), .B1(new_n750), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT114), .B1(new_n765), .B2(KEYINPUT52), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n767), .B(new_n756), .C1(new_n761), .C2(new_n764), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n766), .B2(new_n768), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n741), .B2(new_n683), .ZN(new_n770));
  INV_X1    g569(.A(G99gat), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n771), .B(new_n455), .C1(new_n749), .C2(new_n751), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n772), .B2(new_n641), .ZN(G1338gat));
  NOR3_X1   g572(.A1(new_n365), .A2(G106gat), .A3(new_n641), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n749), .B2(new_n751), .ZN(new_n775));
  INV_X1    g574(.A(G106gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n740), .B2(new_n491), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n774), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n747), .B2(new_n748), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT53), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(G1339gat));
  NOR2_X1   g582(.A1(new_n402), .A2(new_n446), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n626), .A2(new_n633), .A3(new_n627), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT54), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n621), .B1(new_n788), .B2(new_n634), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n636), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n786), .B1(new_n791), .B2(KEYINPUT55), .ZN(new_n792));
  INV_X1    g591(.A(new_n789), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n794));
  AOI211_X1 g593(.A(new_n631), .B(new_n633), .C1(new_n626), .C2(new_n627), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n790), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND4_X1   g595(.A1(new_n786), .A2(new_n793), .A3(new_n796), .A4(KEYINPUT55), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n796), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n639), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n616), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n602), .A2(new_n603), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT116), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n598), .B1(new_n595), .B2(new_n597), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n612), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n601), .A2(new_n604), .A3(new_n605), .A4(new_n613), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n641), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n555), .B1(new_n802), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n808), .B(KEYINPUT117), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n801), .B1(new_n792), .B2(new_n797), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n691), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n593), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n594), .A2(new_n641), .A3(new_n617), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n785), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n365), .A2(new_n447), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT118), .ZN(new_n820));
  INV_X1    g619(.A(G113gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n616), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n816), .A2(new_n371), .ZN(new_n823));
  OAI21_X1  g622(.A(G113gat), .B1(new_n823), .B2(new_n617), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1340gat));
  INV_X1    g624(.A(G120gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n820), .A2(new_n826), .A3(new_n642), .ZN(new_n827));
  OAI21_X1  g626(.A(G120gat), .B1(new_n823), .B2(new_n641), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1341gat));
  AOI21_X1  g628(.A(G127gat), .B1(new_n819), .B2(new_n592), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n823), .A2(new_n254), .A3(new_n593), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(G1342gat));
  NAND3_X1  g631(.A1(new_n819), .A2(new_n258), .A3(new_n555), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT56), .Z(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n823), .B2(new_n691), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1343gat));
  INV_X1    g635(.A(G141gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n683), .A2(new_n784), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n812), .A2(KEYINPUT120), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(new_n801), .C1(new_n792), .C2(new_n797), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n616), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n555), .B1(new_n842), .B2(new_n809), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n593), .B1(new_n843), .B2(new_n813), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT121), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n846), .B(new_n593), .C1(new_n843), .C2(new_n813), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n815), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n491), .A2(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n814), .A2(new_n815), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n491), .ZN(new_n852));
  XNOR2_X1  g651(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n838), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n837), .B1(new_n855), .B2(new_n616), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n852), .A2(new_n838), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n837), .A3(new_n616), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT122), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT58), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n859), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n617), .B(new_n838), .C1(new_n850), .C2(new_n854), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n837), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1344gat));
  INV_X1    g664(.A(G148gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n857), .A2(new_n866), .A3(new_n642), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT59), .B(new_n866), .C1(new_n855), .C2(new_n642), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  INV_X1    g668(.A(new_n838), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n852), .A2(new_n853), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n844), .A2(new_n815), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n491), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n642), .B(new_n870), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n869), .B1(new_n874), .B2(G148gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n867), .B1(new_n868), .B2(new_n875), .ZN(G1345gat));
  AOI21_X1  g675(.A(new_n304), .B1(new_n857), .B2(new_n592), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n592), .A2(new_n304), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n855), .B2(new_n878), .ZN(G1346gat));
  INV_X1    g678(.A(G162gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n857), .A2(new_n880), .A3(new_n555), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n855), .A2(new_n555), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n880), .ZN(G1347gat));
  AOI21_X1  g682(.A(new_n492), .B1(new_n814), .B2(new_n815), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n402), .A3(new_n371), .ZN(new_n885));
  OAI21_X1  g684(.A(G169gat), .B1(new_n885), .B2(new_n617), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n887), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n818), .A2(new_n402), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT124), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n617), .A2(G169gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(G1348gat));
  NOR3_X1   g694(.A1(new_n885), .A2(new_n619), .A3(new_n641), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n890), .A2(new_n642), .A3(new_n892), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n619), .ZN(G1349gat));
  OAI21_X1  g697(.A(G183gat), .B1(new_n885), .B2(new_n593), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n888), .A2(new_n225), .A3(new_n889), .A4(new_n892), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n593), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g701(.A1(new_n691), .A2(G190gat), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n889), .A3(new_n892), .A4(new_n903), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n884), .A2(new_n555), .A3(new_n402), .A4(new_n371), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(G190gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n905), .B2(G190gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n909), .B(new_n910), .ZN(G1351gat));
  OR2_X1    g710(.A1(new_n871), .A2(new_n873), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n457), .A2(new_n492), .A3(new_n448), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n617), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n457), .A2(new_n448), .ZN(new_n916));
  AND4_X1   g715(.A1(new_n491), .A2(new_n888), .A3(new_n889), .A4(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n617), .A2(G197gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1352gat));
  XOR2_X1   g719(.A(KEYINPUT126), .B(G204gat), .Z(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n642), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n912), .A2(new_n642), .A3(new_n913), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n921), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n917), .A2(new_n927), .A3(new_n642), .A4(new_n922), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n917), .A2(new_n319), .A3(new_n592), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n592), .B(new_n913), .C1(new_n871), .C2(new_n873), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n931), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT63), .B1(new_n931), .B2(G211gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(G1354gat));
  NOR3_X1   g733(.A1(new_n914), .A2(new_n320), .A3(new_n691), .ZN(new_n935));
  AOI21_X1  g734(.A(G218gat), .B1(new_n917), .B2(new_n555), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(G1355gat));
endmodule


