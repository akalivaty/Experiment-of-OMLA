//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT27), .B(G183gat), .Z(new_n211));
  OAI21_X1  g010(.A(KEYINPUT28), .B1(new_n211), .B2(G190gat), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n211), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n209), .A2(new_n210), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT64), .B1(new_n216), .B2(new_n205), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(new_n210), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n219), .B2(new_n210), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n217), .A2(KEYINPUT25), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT25), .B1(new_n217), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n214), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G127gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n233), .ZN(new_n235));
  INV_X1    g034(.A(G127gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G134gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI22_X1  g037(.A1(new_n227), .A2(new_n230), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n226), .A2(new_n232), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n242), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(new_n214), .C1(new_n222), .C2(new_n223), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT70), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G15gat), .B(G43gat), .Z(new_n250));
  XNOR2_X1  g049(.A(G71gat), .B(G99gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n247), .B1(new_n243), .B2(new_n245), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT33), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT32), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(new_n252), .C1(new_n253), .C2(new_n255), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT34), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n248), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n252), .A2(KEYINPUT33), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(KEYINPUT32), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n260), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n261), .B1(new_n260), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n249), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n267), .ZN(new_n269));
  INV_X1    g068(.A(new_n249), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n265), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT87), .B(KEYINPUT35), .Z(new_n275));
  NAND3_X1  g074(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT86), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  INV_X1    g077(.A(G85gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G57gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n284));
  XNOR2_X1  g083(.A(G141gat), .B(G148gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT2), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT78), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT78), .B(KEYINPUT2), .C1(new_n287), .C2(new_n288), .ZN(new_n292));
  XNOR2_X1  g091(.A(G155gat), .B(G162gat), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n286), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n293), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n285), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n244), .B1(KEYINPUT3), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n298), .B2(KEYINPUT3), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n294), .A2(new_n297), .A3(KEYINPUT79), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OR3_X1    g103(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n298), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT4), .B1(new_n242), .B2(new_n298), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n299), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n308), .B(KEYINPUT80), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n242), .B(new_n298), .Z(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(new_n310), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n284), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT5), .B1(new_n307), .B2(new_n310), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n283), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n316), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n313), .B1(new_n310), .B2(new_n307), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n318), .B(new_n282), .C1(new_n319), .C2(new_n284), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT6), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n315), .A2(new_n316), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT6), .A3(new_n282), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n224), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n224), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n329), .B2(new_n326), .ZN(new_n330));
  XOR2_X1   g129(.A(G211gat), .B(G218gat), .Z(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT71), .ZN(new_n332));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333));
  INV_X1    g132(.A(G211gat), .ZN(new_n334));
  INV_X1    g133(.A(G218gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n333), .B1(KEYINPUT22), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n332), .B(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G8gat), .B(G36gat), .Z(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n338), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n327), .B(new_n346), .C1(new_n329), .C2(new_n326), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n339), .A2(KEYINPUT30), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n339), .A2(new_n347), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n349), .A2(new_n350), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n351), .B2(new_n344), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n339), .A2(KEYINPUT75), .A3(new_n345), .A4(new_n347), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT30), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT76), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359));
  AOI211_X1 g158(.A(new_n359), .B(KEYINPUT30), .C1(new_n354), .C2(new_n355), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n325), .B(new_n352), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n363));
  INV_X1    g162(.A(G228gat), .ZN(new_n364));
  INV_X1    g163(.A(G233gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n302), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n366));
  AOI211_X1 g165(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(new_n298), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n301), .B2(new_n303), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(new_n346), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n369), .B2(KEYINPUT81), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n368), .A2(new_n371), .A3(new_n346), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n368), .A2(new_n346), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n371), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n376));
  INV_X1    g175(.A(new_n372), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .A4(new_n367), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n337), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n380), .A2(new_n331), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n328), .B1(new_n380), .B2(new_n331), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n302), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n298), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n374), .A2(new_n384), .B1(G228gat), .B2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n363), .B1(new_n379), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI211_X1 g187(.A(KEYINPUT83), .B(new_n385), .C1(new_n373), .C2(new_n378), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G50gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(G50gat), .B1(new_n387), .B2(new_n389), .ZN(new_n393));
  XOR2_X1   g192(.A(G78gat), .B(G106gat), .Z(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(G22gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT31), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n393), .ZN(new_n398));
  INV_X1    g197(.A(new_n396), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n362), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n202), .B1(new_n277), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n397), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n403), .A2(new_n361), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT86), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT86), .B1(new_n268), .B2(new_n271), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n405), .A2(new_n408), .A3(KEYINPUT88), .A4(new_n275), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n268), .A2(new_n271), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT35), .B1(new_n401), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n402), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n397), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n352), .B1(new_n358), .B2(new_n360), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT39), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n312), .B2(new_n310), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n417), .A2(KEYINPUT84), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(KEYINPUT84), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n418), .B(new_n419), .C1(new_n310), .C2(new_n307), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n307), .A2(new_n310), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n282), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(KEYINPUT40), .A3(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n420), .A2(new_n422), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n424), .A2(KEYINPUT40), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n415), .A2(new_n320), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n351), .A2(KEYINPUT37), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT38), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n345), .B1(new_n351), .B2(KEYINPUT37), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n325), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n354), .B2(new_n355), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n431), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n432), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n414), .A2(new_n426), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n413), .A2(new_n361), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n272), .B(KEYINPUT36), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n412), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(G57gat), .B(G64gat), .Z(new_n443));
  NAND2_X1  g242(.A1(G71gat), .A2(G78gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT9), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G71gat), .ZN(new_n448));
  INV_X1    g247(.A(G78gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT99), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT99), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(G71gat), .B2(G78gat), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT98), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n444), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(KEYINPUT98), .A2(G71gat), .A3(G78gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT100), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n450), .A2(new_n452), .ZN(new_n459));
  AND3_X1   g258(.A1(KEYINPUT98), .A2(G71gat), .A3(G78gat), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT98), .B1(G71gat), .B2(G78gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT100), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n447), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n443), .A2(new_n446), .ZN(new_n466));
  INV_X1    g265(.A(new_n444), .ZN(new_n467));
  NOR2_X1   g266(.A1(G71gat), .A2(G78gat), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT21), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(KEYINPUT21), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT96), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT16), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(G1gat), .ZN(new_n478));
  INV_X1    g277(.A(G8gat), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(new_n479), .C1(G1gat), .C2(new_n476), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n476), .A2(G1gat), .ZN(new_n481));
  INV_X1    g280(.A(G1gat), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n475), .B1(KEYINPUT16), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(G8gat), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  MUX2_X1   g284(.A(new_n472), .B(new_n473), .S(new_n485), .Z(new_n486));
  NAND2_X1  g285(.A1(G231gat), .A2(G233gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT101), .Z(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G183gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(new_n334), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n486), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G127gat), .B(G155gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n491), .B(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(G134gat), .B(G162gat), .Z(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT91), .B(G29gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT92), .B(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(G43gat), .A2(G50gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(G43gat), .A2(G50gat), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT15), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OR3_X1    g302(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT94), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n501), .A2(KEYINPUT15), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT93), .B(G43gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n511), .B2(G50gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n507), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n512), .A2(new_n508), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n504), .A2(KEYINPUT90), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n505), .B1(new_n504), .B2(KEYINPUT90), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n500), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n503), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT95), .B1(new_n522), .B2(KEYINPUT17), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n521), .A2(new_n525), .ZN(new_n528));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529));
  INV_X1    g328(.A(G92gat), .ZN(new_n530));
  AOI22_X1  g329(.A1(KEYINPUT8), .A2(new_n529), .B1(new_n279), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n279), .B2(new_n530), .ZN(new_n533));
  NAND3_X1  g332(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n529), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n535), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT102), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n528), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n527), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n521), .A2(new_n538), .B1(KEYINPUT41), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n497), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n542), .A2(KEYINPUT41), .ZN(new_n546));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n497), .A3(new_n543), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n545), .B2(new_n549), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OR3_X1    g351(.A1(new_n495), .A2(new_n552), .A3(KEYINPUT103), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT103), .B1(new_n495), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n528), .A2(new_n485), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n527), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n485), .A2(new_n521), .ZN(new_n558));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n561), .B2(new_n562), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n557), .A2(new_n566), .A3(new_n558), .A4(new_n563), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n485), .B(new_n522), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n559), .B(KEYINPUT13), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n572));
  XNOR2_X1  g371(.A(G113gat), .B(G141gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT12), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n565), .A2(new_n570), .A3(new_n579), .A4(new_n567), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n538), .B1(new_n465), .B2(new_n469), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n463), .B1(new_n459), .B2(new_n462), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n466), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OR3_X1    g388(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n535), .A2(new_n529), .A3(new_n536), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n531), .A2(new_n537), .A3(new_n533), .A4(new_n534), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n584), .A2(KEYINPUT104), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT104), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n470), .A2(new_n596), .A3(new_n593), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT10), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n586), .B1(new_n598), .B2(KEYINPUT105), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT105), .ZN(new_n600));
  AOI211_X1 g399(.A(new_n600), .B(KEYINPUT10), .C1(new_n595), .C2(new_n597), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n583), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n595), .A2(new_n597), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n583), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n607), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n555), .A2(new_n582), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n442), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(new_n325), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n482), .ZN(G1324gat));
  INV_X1    g415(.A(new_n415), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT42), .B1(new_n618), .B2(new_n479), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT16), .B(G8gat), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  MUX2_X1   g420(.A(KEYINPUT42), .B(new_n619), .S(new_n621), .Z(G1325gat));
  INV_X1    g421(.A(new_n614), .ZN(new_n623));
  INV_X1    g422(.A(new_n440), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n623), .A2(G15gat), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(G15gat), .B1(new_n623), .B2(new_n408), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(G1326gat));
  NOR2_X1   g426(.A1(new_n614), .A2(new_n414), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT43), .B(G22gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1327gat));
  INV_X1    g429(.A(new_n552), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n412), .B2(new_n441), .ZN(new_n632));
  INV_X1    g431(.A(new_n495), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n582), .A2(new_n633), .A3(new_n612), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n635), .A2(new_n325), .A3(new_n498), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT45), .Z(new_n637));
  INV_X1    g436(.A(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n442), .A2(new_n552), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT44), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n638), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n498), .B1(new_n644), .B2(new_n325), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n637), .A2(new_n645), .ZN(G1328gat));
  INV_X1    g445(.A(new_n635), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n617), .A2(new_n499), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT106), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n651), .A3(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n499), .B1(new_n644), .B2(new_n617), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n650), .A2(KEYINPUT46), .A3(new_n652), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(G1329gat));
  INV_X1    g457(.A(new_n408), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n635), .A2(new_n659), .A3(new_n511), .ZN(new_n660));
  INV_X1    g459(.A(new_n642), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n632), .A2(new_n641), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n624), .B(new_n634), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n660), .B1(new_n663), .B2(new_n511), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT47), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n510), .B1(new_n643), .B2(new_n624), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(new_n660), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(G1330gat));
  NOR3_X1   g468(.A1(new_n635), .A2(G50gat), .A3(new_n414), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n413), .B(new_n634), .C1(new_n661), .C2(new_n662), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(G50gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT48), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT48), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n391), .B1(new_n643), .B2(new_n413), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(new_n670), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(G1331gat));
  NOR3_X1   g476(.A1(new_n555), .A2(new_n581), .A3(new_n611), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n442), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n433), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G57gat), .ZN(G1332gat));
  INV_X1    g480(.A(KEYINPUT49), .ZN(new_n682));
  INV_X1    g481(.A(G64gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n415), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT107), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n688));
  AND4_X1   g487(.A1(new_n682), .A2(new_n687), .A3(new_n683), .A4(new_n688), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n687), .A2(new_n688), .B1(new_n682), .B2(new_n683), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(G1333gat));
  AOI21_X1  g490(.A(new_n448), .B1(new_n679), .B2(new_n624), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n659), .A2(G71gat), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n679), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n413), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g496(.A1(new_n633), .A2(new_n581), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n611), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n640), .B2(new_n642), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G85gat), .B1(new_n703), .B2(new_n325), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n611), .A2(G85gat), .A3(new_n325), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT110), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n699), .B1(new_n639), .B2(KEYINPUT109), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n632), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT51), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n698), .B1(new_n632), .B2(new_n708), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT51), .ZN(new_n712));
  AOI211_X1 g511(.A(KEYINPUT109), .B(new_n631), .C1(new_n412), .C2(new_n441), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n706), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n704), .A2(new_n715), .ZN(G1336gat));
  NOR3_X1   g515(.A1(new_n617), .A2(G92gat), .A3(new_n611), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT111), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n712), .B1(new_n711), .B2(new_n713), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n639), .A2(KEYINPUT109), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n720), .A2(KEYINPUT51), .A3(new_n698), .A4(new_n709), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n718), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n530), .B1(new_n702), .B2(new_n415), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT52), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n415), .B(new_n700), .C1(new_n661), .C2(new_n662), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT52), .B1(new_n725), .B2(G92gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n717), .B1(new_n710), .B2(new_n714), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(G1337gat));
  OAI21_X1  g528(.A(G99gat), .B1(new_n703), .B2(new_n440), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n659), .A2(G99gat), .A3(new_n611), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n710), .B2(new_n714), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1338gat));
  NOR3_X1   g532(.A1(new_n414), .A2(G106gat), .A3(new_n611), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT112), .Z(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n719), .B2(new_n721), .ZN(new_n736));
  INV_X1    g535(.A(G106gat), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n702), .B2(new_n413), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT53), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n413), .B(new_n700), .C1(new_n661), .C2(new_n662), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT53), .B1(new_n740), .B2(G106gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n734), .B1(new_n710), .B2(new_n714), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(G1339gat));
  NAND2_X1  g543(.A1(new_n603), .A2(new_n585), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n600), .ZN(new_n746));
  INV_X1    g545(.A(new_n583), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n598), .A2(KEYINPUT105), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n586), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n602), .A2(new_n749), .A3(KEYINPUT54), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n583), .C1(new_n599), .C2(new_n601), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n750), .A2(KEYINPUT55), .A3(new_n607), .A4(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n607), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n757), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n750), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n602), .A2(new_n749), .A3(KEYINPUT54), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n756), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n755), .A2(new_n609), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT114), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n757), .A2(new_n750), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n608), .B1(new_n764), .B2(new_n759), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n765), .A2(new_n766), .A3(new_n758), .A4(new_n755), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n582), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g567(.A(new_n485), .B(new_n528), .C1(new_n523), .C2(new_n526), .ZN(new_n769));
  INV_X1    g568(.A(new_n558), .ZN(new_n770));
  OAI211_X1 g569(.A(KEYINPUT115), .B(new_n560), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n568), .A2(new_n569), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n557), .A2(new_n558), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT115), .B1(new_n774), .B2(new_n560), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n576), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n580), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n611), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n631), .B1(new_n768), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n767), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT116), .B1(new_n776), .B2(new_n580), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n776), .A2(KEYINPUT116), .A3(new_n580), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n781), .B(new_n552), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n633), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n553), .A2(new_n582), .A3(new_n554), .A4(new_n611), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n325), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n659), .A2(new_n413), .A3(new_n415), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G113gat), .B1(new_n791), .B2(new_n582), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n780), .A2(new_n784), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n495), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n786), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n413), .A2(new_n415), .A3(new_n410), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n433), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n582), .A2(G113gat), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(G1340gat));
  OAI21_X1  g598(.A(G120gat), .B1(new_n791), .B2(new_n611), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n611), .A2(G120gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n797), .B2(new_n801), .ZN(G1341gat));
  NOR3_X1   g601(.A1(new_n791), .A2(new_n236), .A3(new_n495), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n789), .A2(new_n633), .A3(new_n796), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n236), .B2(new_n804), .ZN(G1342gat));
  NAND2_X1  g604(.A1(new_n552), .A2(new_n231), .ZN(new_n806));
  OR3_X1    g605(.A1(new_n797), .A2(KEYINPUT56), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G134gat), .B1(new_n791), .B2(new_n631), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT56), .B1(new_n797), .B2(new_n806), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT117), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n807), .A2(new_n808), .A3(new_n812), .A4(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1343gat));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n789), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT118), .B1(new_n788), .B2(new_n325), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n440), .A2(new_n413), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n415), .B1(new_n819), .B2(KEYINPUT119), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(KEYINPUT119), .B2(new_n819), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n582), .A2(G141gat), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT120), .Z(new_n824));
  NAND3_X1  g623(.A1(new_n818), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n795), .A2(new_n826), .A3(new_n413), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n581), .A2(new_n758), .A3(new_n765), .A4(new_n755), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n552), .B1(new_n778), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n633), .B1(new_n784), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n413), .B1(new_n831), .B2(new_n787), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT57), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n624), .A2(new_n325), .A3(new_n415), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n827), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G141gat), .B1(new_n835), .B2(new_n582), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT58), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n825), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1344gat));
  INV_X1    g640(.A(G148gat), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n818), .A2(new_n842), .A3(new_n612), .A4(new_n822), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n552), .B1(new_n783), .B2(new_n782), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n762), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n495), .B1(new_n846), .B2(new_n829), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n786), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n848), .B2(new_n413), .ZN(new_n849));
  OAI211_X1 g648(.A(KEYINPUT57), .B(new_n413), .C1(new_n785), .C2(new_n787), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n795), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n413), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n612), .A3(new_n834), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n844), .B1(new_n855), .B2(G148gat), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n835), .A2(new_n611), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(KEYINPUT59), .A3(new_n842), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n843), .B1(new_n856), .B2(new_n858), .ZN(G1345gat));
  NOR3_X1   g658(.A1(new_n835), .A2(new_n287), .A3(new_n495), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n818), .A2(new_n633), .A3(new_n822), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n287), .ZN(G1346gat));
  OAI21_X1  g661(.A(G162gat), .B1(new_n835), .B2(new_n631), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n818), .A2(new_n822), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n552), .A2(new_n288), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(G1347gat));
  NAND2_X1  g665(.A1(new_n415), .A2(new_n325), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n659), .A2(new_n413), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n795), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869), .B2(new_n582), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT122), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n413), .A2(new_n617), .A3(new_n410), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n795), .A2(new_n325), .A3(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n582), .A2(G169gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(G1348gat));
  NAND4_X1  g674(.A1(new_n795), .A2(G176gat), .A3(new_n612), .A4(new_n868), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(G176gat), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n788), .A2(new_n433), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n612), .A3(new_n872), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(G1349gat));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n495), .A2(new_n211), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n873), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n879), .A2(KEYINPUT123), .A3(new_n872), .A4(new_n883), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G183gat), .B1(new_n869), .B2(new_n495), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT60), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1350gat));
  OR3_X1    g692(.A1(new_n873), .A2(G190gat), .A3(new_n631), .ZN(new_n894));
  OAI21_X1  g693(.A(G190gat), .B1(new_n869), .B2(new_n631), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(KEYINPUT61), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(KEYINPUT61), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n819), .A2(new_n617), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  XOR2_X1   g700(.A(KEYINPUT124), .B(G197gat), .Z(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n581), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n624), .A2(new_n867), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n905), .B1(new_n852), .B2(new_n853), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n582), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n903), .B1(new_n908), .B2(new_n902), .ZN(G1352gat));
  XNOR2_X1  g708(.A(KEYINPUT125), .B(G204gat), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n611), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n900), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT62), .ZN(new_n913));
  AOI211_X1 g712(.A(new_n611), .B(new_n905), .C1(new_n852), .C2(new_n853), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND4_X1   g715(.A1(new_n915), .A2(new_n854), .A3(new_n612), .A4(new_n904), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(G1353gat));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n334), .A3(new_n633), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n920), .B(new_n334), .C1(new_n906), .C2(new_n633), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n850), .A2(new_n851), .ZN(new_n922));
  INV_X1    g721(.A(new_n849), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n850), .A2(new_n851), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n633), .B(new_n904), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT63), .B1(new_n926), .B2(G211gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n919), .B1(new_n921), .B2(new_n927), .ZN(G1354gat));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n335), .B1(new_n900), .B2(new_n631), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n631), .A2(new_n335), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n905), .B(new_n933), .C1(new_n852), .C2(new_n853), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(KEYINPUT127), .B(new_n930), .C1(new_n907), .C2(new_n933), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1355gat));
endmodule


