//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  INV_X1    g000(.A(KEYINPUT31), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G128), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n188), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT68), .A4(G128), .ZN(new_n200));
  INV_X1    g014(.A(new_n190), .ZN(new_n201));
  OAI21_X1  g015(.A(G128), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n190), .A2(new_n192), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n195), .A2(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G137), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n207), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n205), .A2(G134), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT65), .A3(new_n211), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n209), .A2(new_n210), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n208), .A3(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n219), .B(G131), .C1(new_n218), .C2(new_n215), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n204), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR3_X1   g037(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n203), .B(new_n223), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n199), .A2(KEYINPUT0), .A3(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT11), .B1(new_n205), .B2(G134), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n206), .B(new_n208), .C1(new_n230), .C2(KEYINPUT65), .ZN(new_n231));
  INV_X1    g045(.A(new_n216), .ZN(new_n232));
  OAI21_X1  g046(.A(G131), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n229), .B1(new_n217), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT30), .B1(new_n222), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n195), .A2(new_n200), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n202), .A2(new_n203), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n217), .A2(new_n220), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT30), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n233), .A2(new_n217), .ZN(new_n242));
  INV_X1    g056(.A(new_n229), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n235), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT69), .B1(new_n248), .B2(G119), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  INV_X1    g064(.A(G119), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(G119), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n249), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n249), .A2(new_n252), .A3(new_n253), .ZN(new_n257));
  INV_X1    g071(.A(new_n255), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT70), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n254), .A2(new_n260), .A3(new_n255), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n256), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n246), .A2(new_n247), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n257), .A2(KEYINPUT70), .A3(new_n258), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n260), .B1(new_n254), .B2(new_n255), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n264), .A2(new_n265), .B1(new_n255), .B2(new_n254), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n235), .B2(new_n245), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n240), .A2(new_n266), .A3(new_n244), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n263), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G953), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT72), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G953), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G237), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(G210), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT27), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G101), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n187), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n280), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n240), .A2(new_n244), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n262), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n240), .A2(KEYINPUT73), .A3(new_n244), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT28), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n262), .B1(new_n222), .B2(new_n234), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(new_n268), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n283), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n269), .B1(new_n246), .B2(new_n262), .ZN(new_n293));
  AOI211_X1 g107(.A(KEYINPUT71), .B(new_n266), .C1(new_n235), .C2(new_n245), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n187), .B(new_n280), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G472), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n285), .B1(new_n222), .B2(new_n234), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n287), .A3(new_n266), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n289), .ZN(new_n302));
  INV_X1    g116(.A(new_n291), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT29), .A4(new_n280), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n298), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n263), .B(new_n283), .C1(new_n267), .C2(new_n269), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n291), .B1(new_n289), .B2(new_n301), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT29), .B1(new_n307), .B2(new_n280), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n305), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT74), .B1(new_n309), .B2(new_n297), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n295), .A2(new_n292), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n297), .B(new_n298), .C1(new_n311), .C2(new_n281), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n308), .A2(new_n306), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n315), .B(G472), .C1(new_n316), .C2(new_n305), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n299), .A2(new_n310), .A3(new_n314), .A4(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G217), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(G234), .B2(new_n298), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G140), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT16), .B(new_n324), .C1(new_n328), .C2(new_n322), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G146), .ZN(new_n333));
  INV_X1    g147(.A(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n251), .A2(G128), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT75), .A2(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT75), .B(KEYINPUT23), .Z(new_n342));
  OAI211_X1 g156(.A(new_n336), .B(new_n341), .C1(new_n342), .C2(new_n335), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n339), .B1(new_n343), .B2(G110), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT77), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n189), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n333), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n337), .A2(new_n338), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(new_n343), .B2(G110), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n329), .A2(new_n189), .A3(new_n331), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n189), .B1(new_n329), .B2(new_n331), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(G221), .A2(G234), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n272), .A2(new_n274), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n361), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n359), .A3(new_n355), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n354), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n348), .A3(new_n353), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n298), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n367), .A2(KEYINPUT25), .A3(new_n298), .A4(new_n368), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n321), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n365), .A2(new_n348), .A3(new_n353), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n365), .B1(new_n353), .B2(new_n348), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n320), .A2(G902), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n318), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G469), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G107), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n382), .A2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT80), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n390), .A3(KEYINPUT3), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n386), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G101), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n243), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n389), .A2(new_n391), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  INV_X1    g213(.A(new_n386), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT81), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n392), .A2(new_n403), .A3(new_n399), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT4), .B1(new_n392), .B2(new_n399), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n397), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n383), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(KEYINPUT82), .B2(new_n385), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(KEYINPUT82), .B2(new_n385), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G101), .ZN(new_n413));
  INV_X1    g227(.A(new_n192), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n203), .A2(new_n334), .B1(new_n414), .B2(KEYINPUT1), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n236), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n401), .A2(KEYINPUT81), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n403), .B1(new_n392), .B2(new_n399), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n413), .B(new_n416), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT10), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n242), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n405), .A2(KEYINPUT10), .A3(new_n238), .A4(new_n413), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n409), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n275), .A2(G227), .ZN(new_n425));
  XOR2_X1   g239(.A(G110), .B(G140), .Z(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n402), .A2(new_n404), .B1(G101), .B2(new_n412), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n419), .B1(new_n430), .B2(new_n238), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT12), .A3(new_n242), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n242), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n429), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n405), .A2(new_n413), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n238), .A2(KEYINPUT10), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n406), .B1(new_n402), .B2(new_n404), .ZN(new_n439));
  OAI22_X1  g253(.A1(new_n437), .A2(new_n438), .B1(new_n439), .B2(new_n396), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT10), .B1(new_n430), .B2(new_n416), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n242), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n428), .B1(new_n442), .B2(new_n424), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n381), .B(new_n298), .C1(new_n436), .C2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n381), .A2(new_n298), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n424), .A2(new_n428), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n442), .ZN(new_n448));
  INV_X1    g262(.A(new_n424), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n432), .B2(new_n435), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n448), .B(G469), .C1(new_n450), .C2(new_n428), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G221), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT9), .B(G234), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT79), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n453), .B1(new_n456), .B2(new_n298), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G214), .B1(G237), .B2(G902), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT83), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n249), .A2(new_n252), .A3(KEYINPUT5), .A4(new_n253), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n248), .A2(KEYINPUT5), .A3(G119), .ZN(new_n463));
  INV_X1    g277(.A(G113), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n264), .A2(new_n265), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n413), .B(new_n466), .C1(new_n417), .C2(new_n418), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n262), .A2(new_n395), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n467), .B1(new_n439), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G122), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n467), .B(new_n470), .C1(new_n439), .C2(new_n468), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(KEYINPUT6), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n475), .A3(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n229), .A2(G125), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n238), .B2(G125), .ZN(new_n478));
  INV_X1    g292(.A(G224), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(G953), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n478), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(new_n479), .B2(G953), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n483), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n477), .B(new_n485), .C1(new_n238), .C2(G125), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n262), .A2(new_n395), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n408), .A2(new_n488), .B1(new_n430), .B2(new_n466), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n489), .B2(new_n470), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n470), .B(KEYINPUT8), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n430), .A2(new_n466), .ZN(new_n492));
  INV_X1    g306(.A(new_n467), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n482), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G210), .B1(G237), .B2(G902), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n498), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n482), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n461), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n459), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT20), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n382), .ZN(new_n507));
  INV_X1    g321(.A(new_n324), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n345), .B2(KEYINPUT76), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G146), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n347), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n275), .A2(G143), .A3(G214), .A4(new_n276), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n272), .A2(new_n274), .A3(G214), .A4(new_n276), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n191), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT85), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT18), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(new_n210), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n511), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(G131), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n517), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n515), .A2(G131), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n210), .B1(new_n512), .B2(new_n514), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n351), .A2(new_n352), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n530), .A3(KEYINPUT17), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n525), .B2(KEYINPUT17), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n351), .A2(new_n352), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT87), .B1(new_n520), .B2(new_n527), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(new_n531), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(KEYINPUT88), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n507), .B(new_n523), .C1(new_n536), .C2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n526), .A2(new_n352), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT19), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n346), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n509), .A2(KEYINPUT19), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT86), .B1(new_n547), .B2(new_n189), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT86), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n546), .A2(new_n549), .A3(G146), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n542), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n523), .ZN(new_n552));
  INV_X1    g366(.A(new_n507), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n541), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(G475), .A2(G902), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n505), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n556), .ZN(new_n558));
  AOI211_X1 g372(.A(KEYINPUT20), .B(new_n558), .C1(new_n541), .C2(new_n554), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n523), .B1(new_n536), .B2(new_n540), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n553), .ZN(new_n561));
  AOI21_X1  g375(.A(G902), .B1(new_n561), .B2(new_n541), .ZN(new_n562));
  INV_X1    g376(.A(G475), .ZN(new_n563));
  OAI22_X1  g377(.A1(new_n557), .A2(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n271), .A2(G952), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G234), .B2(G237), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n298), .B(new_n275), .C1(G234), .C2(G237), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n455), .A2(new_n319), .A3(G953), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G128), .B(G143), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n572), .A2(G134), .ZN(new_n573));
  AND2_X1   g387(.A1(KEYINPUT89), .A2(G122), .ZN(new_n574));
  NOR2_X1   g388(.A1(KEYINPUT89), .A2(G122), .ZN(new_n575));
  OAI21_X1  g389(.A(G116), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n248), .A2(G122), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n384), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(G134), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n577), .A2(KEYINPUT14), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT90), .ZN(new_n582));
  INV_X1    g396(.A(G122), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n582), .B(KEYINPUT14), .C1(new_n583), .C2(G116), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n582), .B1(new_n577), .B2(KEYINPUT14), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n576), .B(new_n581), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G107), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT91), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n590), .A3(G107), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n580), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n576), .A2(new_n577), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G107), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n578), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT13), .B1(new_n334), .B2(G143), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n207), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(new_n572), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n592), .A2(KEYINPUT92), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT92), .ZN(new_n602));
  INV_X1    g416(.A(new_n580), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n587), .A2(new_n590), .A3(G107), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n590), .B1(new_n587), .B2(G107), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n606), .B2(new_n599), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n571), .B1(new_n601), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT92), .B1(new_n592), .B2(new_n600), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(new_n602), .A3(new_n599), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n570), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n298), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT93), .ZN(new_n613));
  INV_X1    g427(.A(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(KEYINPUT15), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n608), .A2(new_n616), .A3(new_n298), .A4(new_n611), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n613), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n612), .B2(new_n615), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n564), .A2(new_n569), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n380), .A2(new_n504), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  OAI21_X1  g436(.A(new_n298), .B1(new_n311), .B2(new_n281), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n312), .ZN(new_n625));
  INV_X1    g439(.A(new_n379), .ZN(new_n626));
  INV_X1    g440(.A(new_n461), .ZN(new_n627));
  INV_X1    g441(.A(new_n569), .ZN(new_n628));
  INV_X1    g442(.A(new_n501), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n500), .B1(new_n482), .B2(new_n495), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  NOR4_X1   g445(.A1(new_n459), .A2(new_n625), .A3(new_n626), .A4(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT95), .B(G478), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n613), .A2(new_n617), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n601), .A2(new_n607), .A3(new_n571), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n570), .B1(new_n609), .B2(new_n610), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n608), .A2(KEYINPUT33), .A3(new_n611), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n614), .A2(G902), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT94), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n644));
  INV_X1    g458(.A(new_n642), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n644), .B(new_n645), .C1(new_n639), .C2(new_n640), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n635), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n564), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n633), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT34), .B(G104), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  AOI22_X1  g465(.A1(new_n539), .A2(KEYINPUT88), .B1(new_n527), .B2(new_n526), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n534), .A2(new_n535), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n522), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n507), .ZN(new_n655));
  INV_X1    g469(.A(new_n541), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n298), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G475), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(new_n619), .C1(new_n557), .C2(new_n559), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n633), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  AND2_X1   g476(.A1(new_n624), .A2(new_n312), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n371), .A2(new_n372), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n320), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT36), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n365), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n354), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n365), .A2(new_n348), .A3(new_n353), .A4(new_n667), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n377), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT96), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n669), .A2(KEYINPUT96), .A3(new_n377), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n664), .B1(new_n666), .B2(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n373), .A2(new_n675), .A3(KEYINPUT97), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n504), .A2(new_n620), .A3(new_n663), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT37), .B(G110), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT98), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(G12));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n567), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n566), .B(KEYINPUT99), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n659), .A2(new_n687), .ZN(new_n688));
  AND4_X1   g502(.A1(new_n502), .A2(new_n452), .A3(new_n679), .A4(new_n458), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n689), .A3(new_n318), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  NOR2_X1   g505(.A1(new_n629), .A2(new_n630), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT38), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n564), .A2(new_n619), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n373), .A2(new_n675), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n627), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n459), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n687), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  INV_X1    g515(.A(new_n314), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n312), .A2(new_n313), .ZN(new_n703));
  INV_X1    g517(.A(new_n270), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n280), .ZN(new_n705));
  INV_X1    g519(.A(new_n290), .ZN(new_n706));
  INV_X1    g520(.A(new_n268), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(G902), .B1(new_n708), .B2(new_n283), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n297), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n702), .A2(new_n703), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n699), .ZN(new_n713));
  OR3_X1    g527(.A1(new_n459), .A2(KEYINPUT40), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n697), .A2(new_n701), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  INV_X1    g530(.A(KEYINPUT100), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n689), .A2(new_n318), .ZN(new_n718));
  INV_X1    g532(.A(new_n687), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n647), .A2(new_n564), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n717), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n720), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n689), .A3(KEYINPUT100), .A4(new_n318), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  NOR2_X1   g539(.A1(new_n648), .A2(new_n631), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n435), .A2(new_n432), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n447), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n442), .A2(new_n424), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n427), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n731), .B(new_n298), .C1(KEYINPUT101), .C2(new_n381), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n381), .A2(KEYINPUT101), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n443), .B1(new_n727), .B2(new_n447), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n733), .B1(new_n734), .B2(G902), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n457), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n726), .A2(new_n318), .A3(new_n379), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT102), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n738), .B(new_n740), .ZN(G15));
  NOR2_X1   g555(.A1(new_n659), .A2(new_n631), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n318), .A3(new_n379), .A4(new_n737), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  NAND4_X1  g558(.A1(new_n502), .A2(new_n458), .A3(new_n732), .A4(new_n735), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n318), .A3(new_n620), .A4(new_n679), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G119), .ZN(G21));
  XNOR2_X1  g562(.A(new_n379), .B(KEYINPUT103), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n663), .A2(KEYINPUT104), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n751));
  INV_X1    g565(.A(new_n749), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n625), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n745), .A2(new_n694), .A3(new_n569), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT105), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n754), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  NAND2_X1  g575(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n762));
  INV_X1    g576(.A(new_n695), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n624), .A2(new_n312), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n745), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n647), .A2(new_n564), .A3(new_n766), .A4(new_n719), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n629), .A2(new_n461), .A3(new_n630), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT107), .B1(new_n459), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n771), .A2(new_n452), .A3(new_n774), .A4(new_n458), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n318), .A3(new_n379), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n762), .A2(new_n767), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n770), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n762), .A2(new_n767), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n773), .A2(new_n775), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT42), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n299), .A2(new_n317), .A3(new_n310), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n312), .B2(new_n313), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n312), .A2(new_n783), .A3(new_n313), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n752), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n778), .B1(new_n781), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NAND3_X1  g604(.A1(new_n780), .A2(new_n380), .A3(new_n688), .ZN(new_n791));
  XNOR2_X1  g605(.A(KEYINPUT109), .B(G134), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(G36));
  INV_X1    g607(.A(new_n635), .ZN(new_n794));
  INV_X1    g608(.A(new_n640), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT33), .B1(new_n608), .B2(new_n611), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n642), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n644), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n641), .A2(KEYINPUT94), .A3(new_n642), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT43), .B1(new_n800), .B2(new_n564), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n541), .A2(new_n554), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT20), .B1(new_n802), .B2(new_n558), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n555), .A2(new_n505), .A3(new_n556), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n803), .A2(new_n804), .B1(new_n657), .B2(G475), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n647), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n695), .B1(new_n624), .B2(new_n312), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n801), .A2(new_n807), .A3(KEYINPUT44), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n771), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n812), .A3(new_n771), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n801), .A2(new_n807), .A3(new_n808), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n811), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT111), .ZN(new_n818));
  INV_X1    g632(.A(new_n444), .ZN(new_n819));
  INV_X1    g633(.A(new_n432), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT12), .B1(new_n431), .B2(new_n242), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n424), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n822), .A2(new_n427), .B1(new_n442), .B2(new_n447), .ZN(new_n823));
  OAI21_X1  g637(.A(G469), .B1(new_n823), .B2(KEYINPUT45), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n448), .B(KEYINPUT45), .C1(new_n450), .C2(new_n428), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n446), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT46), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n819), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT46), .B(new_n446), .C1(new_n824), .C2(new_n826), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n457), .B(new_n713), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n811), .A2(new_n813), .A3(new_n832), .A4(new_n816), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n818), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G137), .ZN(G39));
  AOI21_X1  g649(.A(new_n457), .B1(new_n829), .B2(new_n830), .ZN(new_n836));
  XNOR2_X1  g650(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n318), .A2(new_n720), .A3(new_n379), .A4(new_n772), .ZN(new_n839));
  NOR2_X1   g653(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n838), .B(new_n839), .C1(new_n836), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  AND3_X1   g656(.A1(new_n801), .A2(new_n686), .A3(new_n807), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n843), .A2(new_n754), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n737), .A2(KEYINPUT119), .A3(new_n461), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n737), .A2(new_n461), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(new_n693), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT50), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n772), .A2(new_n736), .A3(new_n457), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n764), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n379), .A2(new_n566), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n711), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n711), .A2(new_n852), .A3(KEYINPUT120), .A4(new_n855), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n647), .A2(new_n564), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n844), .A2(new_n771), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n736), .A2(new_n458), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n836), .A2(new_n840), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n865), .B2(new_n838), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n862), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n851), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n868), .A2(KEYINPUT51), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n565), .B1(new_n844), .B2(new_n746), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n858), .A2(new_n859), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n648), .B2(new_n871), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n788), .A2(new_n853), .A3(KEYINPUT48), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT48), .B1(new_n788), .B2(new_n853), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n868), .B2(KEYINPUT51), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT50), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n850), .B(new_n878), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n866), .A2(new_n863), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(KEYINPUT51), .A3(new_n880), .A4(new_n862), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(KEYINPUT121), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n869), .B(new_n875), .C1(new_n877), .C2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n738), .A2(new_n743), .A3(new_n747), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n757), .B2(new_n759), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n789), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n764), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n779), .A2(new_n780), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n619), .A2(new_n687), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n890), .A2(new_n805), .A3(new_n679), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(new_n318), .A3(new_n698), .A4(new_n771), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n791), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n648), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n647), .A2(new_n564), .A3(KEYINPUT115), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n659), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n632), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n621), .A2(new_n899), .A3(new_n680), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n893), .A2(new_n894), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n887), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n768), .A2(new_n690), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n694), .A2(new_n503), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n763), .A2(new_n687), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n712), .A2(new_n698), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n724), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(KEYINPUT52), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n768), .A2(new_n690), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n909), .A2(KEYINPUT116), .B1(new_n721), .B2(new_n723), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT116), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n768), .A2(new_n690), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n906), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n908), .B1(KEYINPUT52), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n885), .A2(new_n789), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT117), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n902), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n907), .B(KEYINPUT52), .ZN(new_n918));
  INV_X1    g732(.A(new_n893), .ZN(new_n919));
  INV_X1    g733(.A(new_n900), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n885), .A3(new_n789), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n894), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n923));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n921), .A2(KEYINPUT53), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n914), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT53), .B1(new_n918), .B2(new_n921), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT54), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n883), .A2(new_n929), .B1(G952), .B2(G953), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n749), .A2(new_n627), .A3(new_n458), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(KEYINPUT49), .B2(new_n736), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n805), .A3(new_n647), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT113), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n736), .A2(KEYINPUT49), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n934), .A2(new_n711), .A3(new_n693), .A4(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT114), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n930), .A2(new_n937), .ZN(G75));
  NAND2_X1  g752(.A1(new_n917), .A2(new_n922), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(G902), .A3(new_n498), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT56), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n474), .A2(new_n476), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n481), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n940), .B2(new_n941), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n275), .A2(G952), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(G51));
  XNOR2_X1  g762(.A(new_n445), .B(KEYINPUT57), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n917), .A2(new_n922), .A3(new_n923), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n923), .B1(new_n917), .B2(new_n922), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n731), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n824), .A2(new_n826), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n939), .A2(G902), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n947), .B1(new_n953), .B2(new_n955), .ZN(G54));
  NAND4_X1  g770(.A1(new_n939), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n802), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n802), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n947), .ZN(G60));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT59), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n641), .B1(new_n929), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n641), .A2(new_n963), .ZN(new_n965));
  INV_X1    g779(.A(new_n951), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n924), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n964), .A2(new_n967), .A3(new_n947), .ZN(G63));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n917), .B2(new_n922), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n669), .A2(new_n670), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n947), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n972), .B2(new_n376), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n969), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n972), .A2(new_n376), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n979), .A2(KEYINPUT61), .A3(new_n974), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(G66));
  OAI21_X1  g795(.A(G953), .B1(new_n568), .B2(new_n479), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n885), .A2(new_n920), .ZN(new_n983));
  INV_X1    g797(.A(new_n275), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n942), .B1(G898), .B2(new_n275), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT122), .Z(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(G69));
  NAND3_X1  g802(.A1(new_n564), .A2(new_n502), .A3(new_n619), .ZN(new_n989));
  AOI211_X1 g803(.A(new_n752), .B(new_n989), .C1(new_n785), .C2(new_n786), .ZN(new_n990));
  INV_X1    g804(.A(new_n776), .ZN(new_n991));
  AOI22_X1  g805(.A1(new_n990), .A2(new_n831), .B1(new_n991), .B2(new_n688), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n789), .A2(new_n992), .A3(new_n841), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n910), .A2(new_n912), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n995), .A2(new_n275), .A3(new_n834), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n246), .B(new_n547), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n996), .B(new_n997), .C1(new_n684), .C2(new_n275), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n909), .A2(KEYINPUT116), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n999), .A2(new_n715), .A3(new_n724), .A4(new_n912), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n910), .A2(new_n1002), .A3(new_n715), .A4(new_n912), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n700), .A2(new_n772), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n898), .A3(new_n380), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n841), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1001), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n833), .A2(new_n831), .ZN(new_n1008));
  AOI22_X1  g822(.A1(new_n810), .A2(KEYINPUT110), .B1(new_n815), .B2(new_n814), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n832), .B1(new_n1009), .B2(new_n813), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT123), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n841), .A2(new_n1005), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(KEYINPUT62), .B2(new_n1000), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT123), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1014), .A2(new_n834), .A3(new_n1015), .A4(new_n1003), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n984), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n998), .B1(new_n1017), .B2(new_n997), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n275), .B1(G227), .B2(G900), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT124), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1018), .B(new_n1021), .ZN(G72));
  NAND3_X1  g836(.A1(new_n1012), .A2(new_n983), .A3(new_n1016), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n705), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1025), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n704), .A2(new_n280), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n926), .A2(new_n927), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n995), .A2(new_n983), .A3(new_n834), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1034), .A2(KEYINPUT125), .A3(new_n1025), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1030), .B(KEYINPUT126), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(KEYINPUT125), .B1(new_n1034), .B2(new_n1025), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n976), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(KEYINPUT127), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT127), .ZN(new_n1041));
  OAI211_X1 g855(.A(new_n1041), .B(new_n976), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1033), .B1(new_n1040), .B2(new_n1042), .ZN(G57));
endmodule


