

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(n717), .ZN(n709) );
  XNOR2_X1 U551 ( .A(n680), .B(n679), .ZN(n717) );
  NOR2_X1 U552 ( .A1(n792), .A2(n794), .ZN(n680) );
  NAND2_X1 U553 ( .A1(n690), .A2(n689), .ZN(n692) );
  INV_X1 U554 ( .A(KEYINPUT30), .ZN(n720) );
  XNOR2_X1 U555 ( .A(n735), .B(KEYINPUT32), .ZN(n761) );
  INV_X1 U556 ( .A(n952), .ZN(n756) );
  NAND2_X1 U557 ( .A1(n887), .A2(G137), .ZN(n534) );
  XOR2_X1 U558 ( .A(KEYINPUT74), .B(n519), .Z(n516) );
  OR2_X1 U559 ( .A1(n753), .A2(KEYINPUT33), .ZN(n517) );
  INV_X1 U560 ( .A(KEYINPUT97), .ZN(n691) );
  XNOR2_X1 U561 ( .A(n692), .B(n691), .ZN(n697) );
  NAND2_X1 U562 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U563 ( .A1(n734), .A2(G8), .ZN(n735) );
  INV_X1 U564 ( .A(KEYINPUT64), .ZN(n679) );
  INV_X1 U565 ( .A(KEYINPUT17), .ZN(n532) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  NOR2_X1 U567 ( .A1(G651), .A2(n635), .ZN(n644) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n539), .ZN(n895) );
  NOR2_X1 U569 ( .A1(n538), .A2(n537), .ZN(n542) );
  NOR2_X1 U570 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U571 ( .A(KEYINPUT76), .B(KEYINPUT7), .ZN(n531) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n640) );
  NAND2_X1 U573 ( .A1(n640), .A2(G89), .ZN(n518) );
  XOR2_X1 U574 ( .A(KEYINPUT4), .B(n518), .Z(n520) );
  XOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .Z(n635) );
  INV_X1 U576 ( .A(G651), .ZN(n523) );
  NOR2_X1 U577 ( .A1(n635), .A2(n523), .ZN(n641) );
  NAND2_X1 U578 ( .A1(n641), .A2(G76), .ZN(n519) );
  NOR2_X1 U579 ( .A1(n520), .A2(n516), .ZN(n521) );
  XNOR2_X1 U580 ( .A(KEYINPUT5), .B(n521), .ZN(n522) );
  XNOR2_X1 U581 ( .A(n522), .B(KEYINPUT75), .ZN(n529) );
  NAND2_X1 U582 ( .A1(G51), .A2(n644), .ZN(n526) );
  NOR2_X1 U583 ( .A1(G543), .A2(n523), .ZN(n524) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n524), .Z(n638) );
  NAND2_X1 U585 ( .A1(G63), .A2(n638), .ZN(n525) );
  NAND2_X1 U586 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U587 ( .A(KEYINPUT6), .B(n527), .Z(n528) );
  NAND2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U589 ( .A(n531), .B(n530), .ZN(G168) );
  XNOR2_X2 U590 ( .A(n533), .B(n532), .ZN(n887) );
  XNOR2_X1 U591 ( .A(n534), .B(KEYINPUT67), .ZN(n538) );
  INV_X1 U592 ( .A(G2105), .ZN(n539) );
  AND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U594 ( .A1(G113), .A2(n893), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G125), .A2(n895), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n537) );
  AND2_X1 U597 ( .A1(n539), .A2(G2104), .ZN(n889) );
  NAND2_X1 U598 ( .A1(G101), .A2(n889), .ZN(n540) );
  XOR2_X1 U599 ( .A(KEYINPUT23), .B(n540), .Z(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n544) );
  INV_X1 U601 ( .A(KEYINPUT66), .ZN(n543) );
  XNOR2_X2 U602 ( .A(n544), .B(n543), .ZN(G160) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U604 ( .A1(G135), .A2(n887), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G111), .A2(n893), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n895), .A2(G123), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT18), .B(n547), .Z(n548) );
  NOR2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n889), .A2(G99), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n1002) );
  XNOR2_X1 U612 ( .A(G2096), .B(n1002), .ZN(n552) );
  OR2_X1 U613 ( .A1(G2100), .A2(n552), .ZN(G156) );
  NAND2_X1 U614 ( .A1(G53), .A2(n644), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G65), .A2(n638), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G91), .A2(n640), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G78), .A2(n641), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n945) );
  INV_X1 U621 ( .A(n945), .ZN(G299) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  INV_X1 U625 ( .A(G108), .ZN(G238) );
  INV_X1 U626 ( .A(G120), .ZN(G236) );
  NAND2_X1 U627 ( .A1(G90), .A2(n640), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G77), .A2(n641), .ZN(n559) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(KEYINPUT9), .B(n561), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n644), .A2(G52), .ZN(n563) );
  NAND2_X1 U632 ( .A1(G64), .A2(n638), .ZN(n562) );
  AND2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(G301) );
  INV_X1 U635 ( .A(G301), .ZN(G171) );
  NAND2_X1 U636 ( .A1(n887), .A2(G138), .ZN(n567) );
  NAND2_X1 U637 ( .A1(G102), .A2(n889), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U639 ( .A1(G114), .A2(n893), .ZN(n569) );
  NAND2_X1 U640 ( .A1(G126), .A2(n895), .ZN(n568) );
  NAND2_X1 U641 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U642 ( .A1(n571), .A2(n570), .ZN(G164) );
  XOR2_X1 U643 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U645 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n574) );
  INV_X1 U647 ( .A(G223), .ZN(n829) );
  NAND2_X1 U648 ( .A1(G567), .A2(n829), .ZN(n573) );
  XNOR2_X1 U649 ( .A(n574), .B(n573), .ZN(G234) );
  NAND2_X1 U650 ( .A1(G81), .A2(n640), .ZN(n575) );
  XNOR2_X1 U651 ( .A(n575), .B(KEYINPUT72), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U653 ( .A1(G68), .A2(n641), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U655 ( .A(KEYINPUT13), .B(n579), .Z(n583) );
  NAND2_X1 U656 ( .A1(G56), .A2(n638), .ZN(n580) );
  XNOR2_X1 U657 ( .A(n580), .B(KEYINPUT14), .ZN(n581) );
  XNOR2_X1 U658 ( .A(n581), .B(KEYINPUT71), .ZN(n582) );
  NOR2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n644), .A2(G43), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n958) );
  INV_X1 U662 ( .A(n958), .ZN(n651) );
  NAND2_X1 U663 ( .A1(n651), .A2(G860), .ZN(G153) );
  NAND2_X1 U664 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G79), .A2(n641), .ZN(n587) );
  NAND2_X1 U666 ( .A1(G54), .A2(n644), .ZN(n586) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n592) );
  NAND2_X1 U668 ( .A1(G92), .A2(n640), .ZN(n589) );
  NAND2_X1 U669 ( .A1(G66), .A2(n638), .ZN(n588) );
  NAND2_X1 U670 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U671 ( .A(KEYINPUT73), .B(n590), .Z(n591) );
  NOR2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U673 ( .A(KEYINPUT15), .B(n593), .Z(n955) );
  OR2_X1 U674 ( .A1(n955), .A2(G868), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U676 ( .A1(G868), .A2(G286), .ZN(n597) );
  INV_X1 U677 ( .A(G868), .ZN(n660) );
  NAND2_X1 U678 ( .A1(G299), .A2(n660), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n597), .A2(n596), .ZN(G297) );
  INV_X1 U680 ( .A(G559), .ZN(n598) );
  NOR2_X1 U681 ( .A1(G860), .A2(n598), .ZN(n599) );
  XNOR2_X1 U682 ( .A(KEYINPUT77), .B(n599), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n600), .A2(n955), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n958), .ZN(n602) );
  XNOR2_X1 U686 ( .A(KEYINPUT78), .B(n602), .ZN(n605) );
  NAND2_X1 U687 ( .A1(G868), .A2(n955), .ZN(n603) );
  NOR2_X1 U688 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U689 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G93), .A2(n640), .ZN(n607) );
  NAND2_X1 U691 ( .A1(G80), .A2(n641), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U693 ( .A1(G55), .A2(n644), .ZN(n609) );
  NAND2_X1 U694 ( .A1(G67), .A2(n638), .ZN(n608) );
  NAND2_X1 U695 ( .A1(n609), .A2(n608), .ZN(n610) );
  OR2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n661) );
  NAND2_X1 U697 ( .A1(n955), .A2(G559), .ZN(n658) );
  XNOR2_X1 U698 ( .A(n958), .B(n658), .ZN(n612) );
  NOR2_X1 U699 ( .A1(G860), .A2(n612), .ZN(n613) );
  XOR2_X1 U700 ( .A(KEYINPUT79), .B(n613), .Z(n614) );
  XOR2_X1 U701 ( .A(n661), .B(n614), .Z(G145) );
  NAND2_X1 U702 ( .A1(G88), .A2(n640), .ZN(n616) );
  NAND2_X1 U703 ( .A1(G75), .A2(n641), .ZN(n615) );
  NAND2_X1 U704 ( .A1(n616), .A2(n615), .ZN(n621) );
  NAND2_X1 U705 ( .A1(G50), .A2(n644), .ZN(n618) );
  NAND2_X1 U706 ( .A1(G62), .A2(n638), .ZN(n617) );
  NAND2_X1 U707 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U708 ( .A(KEYINPUT82), .B(n619), .ZN(n620) );
  NOR2_X1 U709 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U710 ( .A(n622), .B(KEYINPUT83), .ZN(G303) );
  INV_X1 U711 ( .A(G303), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G86), .A2(n640), .ZN(n624) );
  NAND2_X1 U713 ( .A1(G61), .A2(n638), .ZN(n623) );
  NAND2_X1 U714 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U715 ( .A1(n641), .A2(G73), .ZN(n625) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U717 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U718 ( .A(KEYINPUT80), .B(n628), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n644), .A2(G48), .ZN(n629) );
  XOR2_X1 U720 ( .A(KEYINPUT81), .B(n629), .Z(n630) );
  NAND2_X1 U721 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G49), .A2(n644), .ZN(n633) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U724 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U725 ( .A1(n638), .A2(n634), .ZN(n637) );
  NAND2_X1 U726 ( .A1(n635), .A2(G87), .ZN(n636) );
  NAND2_X1 U727 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U728 ( .A1(n638), .A2(G60), .ZN(n639) );
  XNOR2_X1 U729 ( .A(n639), .B(KEYINPUT68), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G85), .A2(n640), .ZN(n643) );
  NAND2_X1 U731 ( .A1(G72), .A2(n641), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U733 ( .A1(G47), .A2(n644), .ZN(n645) );
  XNOR2_X1 U734 ( .A(KEYINPUT69), .B(n645), .ZN(n646) );
  NOR2_X1 U735 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U736 ( .A1(n649), .A2(n648), .ZN(G290) );
  XNOR2_X1 U737 ( .A(G166), .B(G305), .ZN(n657) );
  XOR2_X1 U738 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n650) );
  XNOR2_X1 U739 ( .A(G288), .B(n650), .ZN(n654) );
  XNOR2_X1 U740 ( .A(n661), .B(n651), .ZN(n652) );
  XNOR2_X1 U741 ( .A(n652), .B(G299), .ZN(n653) );
  XNOR2_X1 U742 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U743 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U744 ( .A(n657), .B(n656), .ZN(n905) );
  XNOR2_X1 U745 ( .A(n905), .B(n658), .ZN(n659) );
  NOR2_X1 U746 ( .A1(n660), .A2(n659), .ZN(n663) );
  NOR2_X1 U747 ( .A1(G868), .A2(n661), .ZN(n662) );
  NOR2_X1 U748 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n664) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U756 ( .A1(G236), .A2(G238), .ZN(n668) );
  NAND2_X1 U757 ( .A1(G69), .A2(n668), .ZN(n669) );
  NOR2_X1 U758 ( .A1(n669), .A2(G237), .ZN(n670) );
  XNOR2_X1 U759 ( .A(n670), .B(KEYINPUT85), .ZN(n834) );
  NAND2_X1 U760 ( .A1(n834), .A2(G567), .ZN(n675) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U763 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U764 ( .A1(G96), .A2(n673), .ZN(n835) );
  NAND2_X1 U765 ( .A1(n835), .A2(G2106), .ZN(n674) );
  NAND2_X1 U766 ( .A1(n675), .A2(n674), .ZN(n836) );
  NOR2_X1 U767 ( .A1(n676), .A2(n836), .ZN(n677) );
  XNOR2_X1 U768 ( .A(n677), .B(KEYINPUT86), .ZN(n833) );
  NAND2_X1 U769 ( .A1(G36), .A2(n833), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G40), .A2(G160), .ZN(n792) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n678) );
  XNOR2_X1 U772 ( .A(KEYINPUT65), .B(n678), .ZN(n794) );
  NAND2_X1 U773 ( .A1(n709), .A2(G1996), .ZN(n681) );
  OR2_X1 U774 ( .A1(n681), .A2(KEYINPUT26), .ZN(n683) );
  NAND2_X1 U775 ( .A1(n681), .A2(KEYINPUT26), .ZN(n682) );
  NAND2_X1 U776 ( .A1(n683), .A2(n682), .ZN(n694) );
  AND2_X1 U777 ( .A1(n717), .A2(G1341), .ZN(n684) );
  NOR2_X1 U778 ( .A1(n684), .A2(n958), .ZN(n693) );
  AND2_X1 U779 ( .A1(n955), .A2(n693), .ZN(n685) );
  NAND2_X1 U780 ( .A1(n694), .A2(n685), .ZN(n686) );
  XNOR2_X1 U781 ( .A(n686), .B(KEYINPUT96), .ZN(n690) );
  NOR2_X1 U782 ( .A1(G1348), .A2(n709), .ZN(n688) );
  NOR2_X1 U783 ( .A1(G2067), .A2(n717), .ZN(n687) );
  NOR2_X1 U784 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  OR2_X1 U786 ( .A1(n955), .A2(n695), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n702) );
  NAND2_X1 U788 ( .A1(G2072), .A2(n709), .ZN(n698) );
  XNOR2_X1 U789 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U790 ( .A(G1956), .ZN(n970) );
  NOR2_X1 U791 ( .A1(n709), .A2(n970), .ZN(n699) );
  NOR2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n945), .A2(n703), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U795 ( .A1(n945), .A2(n703), .ZN(n704) );
  XOR2_X1 U796 ( .A(n704), .B(KEYINPUT28), .Z(n705) );
  XOR2_X1 U797 ( .A(KEYINPUT29), .B(n707), .Z(n738) );
  XOR2_X1 U798 ( .A(KEYINPUT25), .B(G2078), .Z(n925) );
  NOR2_X1 U799 ( .A1(n717), .A2(n925), .ZN(n708) );
  XNOR2_X1 U800 ( .A(n708), .B(KEYINPUT95), .ZN(n711) );
  OR2_X1 U801 ( .A1(n709), .A2(G1961), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n724) );
  NAND2_X1 U803 ( .A1(n724), .A2(G171), .ZN(n739) );
  NOR2_X1 U804 ( .A1(n717), .A2(G2090), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n717), .A2(G8), .ZN(n771) );
  NOR2_X1 U806 ( .A1(G1971), .A2(n771), .ZN(n712) );
  NOR2_X1 U807 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n714), .A2(G303), .ZN(n729) );
  INV_X1 U809 ( .A(n729), .ZN(n715) );
  OR2_X1 U810 ( .A1(n715), .A2(G286), .ZN(n730) );
  AND2_X1 U811 ( .A1(n739), .A2(n730), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n738), .A2(n716), .ZN(n733) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n771), .ZN(n743) );
  NOR2_X1 U814 ( .A1(n717), .A2(G2084), .ZN(n745) );
  INV_X1 U815 ( .A(n745), .ZN(n718) );
  NAND2_X1 U816 ( .A1(G8), .A2(n718), .ZN(n719) );
  OR2_X1 U817 ( .A1(n743), .A2(n719), .ZN(n721) );
  XNOR2_X1 U818 ( .A(n721), .B(n720), .ZN(n723) );
  INV_X1 U819 ( .A(G168), .ZN(n722) );
  AND2_X1 U820 ( .A1(n723), .A2(n722), .ZN(n726) );
  NOR2_X1 U821 ( .A1(G171), .A2(n724), .ZN(n725) );
  NOR2_X1 U822 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U823 ( .A(n727), .B(KEYINPUT31), .Z(n728) );
  XNOR2_X1 U824 ( .A(n728), .B(KEYINPUT98), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n740), .A2(n729), .ZN(n731) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n950) );
  INV_X1 U829 ( .A(n771), .ZN(n736) );
  NAND2_X1 U830 ( .A1(n950), .A2(n736), .ZN(n750) );
  INV_X1 U831 ( .A(n750), .ZN(n737) );
  AND2_X1 U832 ( .A1(n761), .A2(n737), .ZN(n748) );
  NAND2_X1 U833 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U835 ( .A(KEYINPUT99), .B(n742), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U837 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n762) );
  NAND2_X1 U839 ( .A1(n748), .A2(n762), .ZN(n752) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U842 ( .A1(n754), .A2(n749), .ZN(n965) );
  OR2_X1 U843 ( .A1(n750), .A2(n965), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U845 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n771), .A2(n755), .ZN(n757) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n952) );
  NOR2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n517), .A2(n758), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n759) );
  XNOR2_X1 U851 ( .A(n759), .B(KEYINPUT100), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n760), .A2(G8), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n765), .A2(n771), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n815) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XOR2_X1 U858 ( .A(n768), .B(KEYINPUT94), .Z(n769) );
  XNOR2_X1 U859 ( .A(KEYINPUT24), .B(n769), .ZN(n770) );
  NOR2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n813) );
  NAND2_X1 U861 ( .A1(n889), .A2(G105), .ZN(n773) );
  XNOR2_X1 U862 ( .A(KEYINPUT38), .B(KEYINPUT92), .ZN(n772) );
  XNOR2_X1 U863 ( .A(n773), .B(n772), .ZN(n780) );
  NAND2_X1 U864 ( .A1(G141), .A2(n887), .ZN(n775) );
  NAND2_X1 U865 ( .A1(G129), .A2(n895), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G117), .A2(n893), .ZN(n776) );
  XNOR2_X1 U868 ( .A(KEYINPUT91), .B(n776), .ZN(n777) );
  NOR2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n879) );
  NOR2_X1 U871 ( .A1(G1996), .A2(n879), .ZN(n1009) );
  NAND2_X1 U872 ( .A1(G119), .A2(n895), .ZN(n781) );
  XNOR2_X1 U873 ( .A(n781), .B(KEYINPUT88), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G95), .A2(n889), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G107), .A2(n893), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G131), .A2(n887), .ZN(n784) );
  XNOR2_X1 U878 ( .A(KEYINPUT89), .B(n784), .ZN(n785) );
  NOR2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n882) );
  NAND2_X1 U881 ( .A1(G1991), .A2(n882), .ZN(n789) );
  XOR2_X1 U882 ( .A(KEYINPUT90), .B(n789), .Z(n791) );
  AND2_X1 U883 ( .A1(n879), .A2(G1996), .ZN(n790) );
  NOR2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n1007) );
  INV_X1 U885 ( .A(n792), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n799) );
  NOR2_X1 U887 ( .A1(n1007), .A2(n799), .ZN(n818) );
  NOR2_X1 U888 ( .A1(G1986), .A2(G290), .ZN(n795) );
  NOR2_X1 U889 ( .A1(G1991), .A2(n882), .ZN(n1001) );
  NOR2_X1 U890 ( .A1(n795), .A2(n1001), .ZN(n796) );
  NOR2_X1 U891 ( .A1(n818), .A2(n796), .ZN(n797) );
  NOR2_X1 U892 ( .A1(n1009), .A2(n797), .ZN(n798) );
  XNOR2_X1 U893 ( .A(KEYINPUT39), .B(n798), .ZN(n809) );
  INV_X1 U894 ( .A(n799), .ZN(n816) );
  XNOR2_X1 U895 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NAND2_X1 U896 ( .A1(G140), .A2(n887), .ZN(n801) );
  NAND2_X1 U897 ( .A1(G104), .A2(n889), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U899 ( .A(KEYINPUT34), .B(n802), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G116), .A2(n893), .ZN(n804) );
  NAND2_X1 U901 ( .A1(G128), .A2(n895), .ZN(n803) );
  NAND2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U903 ( .A(KEYINPUT35), .B(n805), .Z(n806) );
  NOR2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n808), .ZN(n901) );
  NOR2_X1 U906 ( .A1(n810), .A2(n901), .ZN(n1005) );
  NAND2_X1 U907 ( .A1(n816), .A2(n1005), .ZN(n820) );
  NAND2_X1 U908 ( .A1(n809), .A2(n820), .ZN(n811) );
  NAND2_X1 U909 ( .A1(n810), .A2(n901), .ZN(n1022) );
  NAND2_X1 U910 ( .A1(n811), .A2(n1022), .ZN(n812) );
  AND2_X1 U911 ( .A1(n812), .A2(n816), .ZN(n825) );
  OR2_X1 U912 ( .A1(n813), .A2(n825), .ZN(n814) );
  NOR2_X1 U913 ( .A1(n815), .A2(n814), .ZN(n827) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n949) );
  NAND2_X1 U915 ( .A1(n816), .A2(n949), .ZN(n817) );
  XNOR2_X1 U916 ( .A(KEYINPUT87), .B(n817), .ZN(n823) );
  INV_X1 U917 ( .A(n818), .ZN(n819) );
  NAND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U919 ( .A(KEYINPUT93), .B(n821), .Z(n822) );
  NOR2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U922 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n829), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT101), .B(n830), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n831), .A2(G661), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  NOR2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G325) );
  XOR2_X1 U930 ( .A(KEYINPUT102), .B(G325), .Z(G261) );
  INV_X1 U931 ( .A(n836), .ZN(G319) );
  XOR2_X1 U932 ( .A(G2096), .B(G2090), .Z(n838) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n848) );
  XOR2_X1 U935 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT105), .B(G2678), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U938 ( .A(G2100), .B(KEYINPUT103), .Z(n842) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2084), .B(G2078), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U944 ( .A(n848), .B(n847), .Z(G227) );
  XOR2_X1 U945 ( .A(G1971), .B(G1956), .Z(n850) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1961), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U948 ( .A(G1976), .B(G1966), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U952 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U954 ( .A(G1981), .B(G2474), .Z(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n895), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(KEYINPUT108), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U959 ( .A1(G112), .A2(n893), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G136), .A2(n887), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G100), .A2(n889), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U964 ( .A1(n866), .A2(n865), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G118), .A2(n893), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G130), .A2(n895), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U968 ( .A1(n889), .A2(G106), .ZN(n869) );
  XOR2_X1 U969 ( .A(KEYINPUT109), .B(n869), .Z(n871) );
  NAND2_X1 U970 ( .A1(n887), .A2(G142), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U972 ( .A(n872), .B(KEYINPUT45), .Z(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(G160), .ZN(n886) );
  XOR2_X1 U975 ( .A(KEYINPUT110), .B(KEYINPUT114), .Z(n877) );
  XNOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(n878), .B(G162), .Z(n881) );
  XOR2_X1 U979 ( .A(G164), .B(n879), .Z(n880) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n884), .B(n1002), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n903) );
  NAND2_X1 U984 ( .A1(n887), .A2(G139), .ZN(n888) );
  XOR2_X1 U985 ( .A(KEYINPUT111), .B(n888), .Z(n891) );
  NAND2_X1 U986 ( .A1(n889), .A2(G103), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(KEYINPUT112), .B(n892), .ZN(n900) );
  NAND2_X1 U989 ( .A1(n893), .A2(G115), .ZN(n894) );
  XOR2_X1 U990 ( .A(KEYINPUT113), .B(n894), .Z(n897) );
  NAND2_X1 U991 ( .A1(n895), .A2(G127), .ZN(n896) );
  NAND2_X1 U992 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U994 ( .A1(n900), .A2(n899), .ZN(n1015) );
  XNOR2_X1 U995 ( .A(n901), .B(n1015), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U997 ( .A1(G37), .A2(n904), .ZN(G395) );
  XOR2_X1 U998 ( .A(KEYINPUT115), .B(n905), .Z(n907) );
  XNOR2_X1 U999 ( .A(G171), .B(n955), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1001 ( .A(n908), .B(G286), .Z(n909) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1003 ( .A(G2451), .B(G2430), .Z(n911) );
  XNOR2_X1 U1004 ( .A(G2438), .B(G2443), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n917) );
  XOR2_X1 U1006 ( .A(G2435), .B(G2454), .Z(n913) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G1348), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n915) );
  XOR2_X1 U1009 ( .A(G2446), .B(G2427), .Z(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1011 ( .A(n917), .B(n916), .Z(n918) );
  NAND2_X1 U1012 ( .A1(G14), .A2(n918), .ZN(n924) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n924), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(G225) );
  XOR2_X1 U1019 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1021 ( .A(G96), .ZN(G221) );
  INV_X1 U1022 ( .A(G69), .ZN(G235) );
  INV_X1 U1023 ( .A(n924), .ZN(G401) );
  XOR2_X1 U1024 ( .A(n925), .B(G27), .Z(n936) );
  XOR2_X1 U1025 ( .A(G1991), .B(G25), .Z(n926) );
  NAND2_X1 U1026 ( .A1(G28), .A2(n926), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(n927), .B(KEYINPUT121), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(G2067), .B(G26), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(G32), .B(G1996), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(KEYINPUT122), .B(G2072), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(G33), .B(n932), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(n937), .B(KEYINPUT53), .ZN(n940) );
  XOR2_X1 U1037 ( .A(G2084), .B(G34), .Z(n938) );
  XNOR2_X1 U1038 ( .A(KEYINPUT54), .B(n938), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G35), .B(G2090), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1042 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n1025) );
  XNOR2_X1 U1043 ( .A(n943), .B(n1025), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(G29), .A2(n944), .ZN(n998) );
  XNOR2_X1 U1045 ( .A(KEYINPUT56), .B(G16), .ZN(n968) );
  XNOR2_X1 U1046 ( .A(n945), .B(G1956), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(G1971), .A2(G303), .ZN(n946) );
  NAND2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n964) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(KEYINPUT57), .B(n954), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n955), .B(G1348), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(G171), .B(G1961), .ZN(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(G1341), .B(n958), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT123), .ZN(n995) );
  XNOR2_X1 U1064 ( .A(n970), .B(G20), .ZN(n978) );
  XOR2_X1 U1065 ( .A(G1341), .B(G19), .Z(n973) );
  XOR2_X1 U1066 ( .A(G6), .B(KEYINPUT124), .Z(n971) );
  XNOR2_X1 U1067 ( .A(G1981), .B(n971), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT59), .B(G1348), .Z(n974) );
  XNOR2_X1 U1070 ( .A(G4), .B(n974), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n979), .B(KEYINPUT60), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(G1986), .B(G24), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(G1976), .B(KEYINPUT125), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(n982), .B(G23), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n985), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G21), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(G1961), .B(G5), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT61), .B(n992), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n993), .A2(G16), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(G11), .A2(n996), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT126), .B(n999), .ZN(n1029) );
  XOR2_X1 U1092 ( .A(G2084), .B(G160), .Z(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G2090), .B(G162), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1008), .B(KEYINPUT117), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT51), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(KEYINPUT118), .B(n1014), .Z(n1020) );
  XOR2_X1 U1103 ( .A(G2072), .B(n1015), .Z(n1017) );
  XOR2_X1 U1104 ( .A(G164), .B(G2078), .Z(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1106 ( .A(KEYINPUT50), .B(n1018), .Z(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(n1023), .B(KEYINPUT119), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT52), .B(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(G29), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1114 ( .A(n1030), .B(KEYINPUT62), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1031), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

