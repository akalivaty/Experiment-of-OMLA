//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(G143), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n189), .B1(new_n194), .B2(KEYINPUT1), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n193), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(new_n196), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n188), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n197), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G143), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n202), .B2(G143), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT69), .B(new_n203), .C1(new_n205), .C2(new_n189), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n190), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n194), .A2(new_n204), .A3(G128), .A4(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT67), .B1(new_n212), .B2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G134), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(KEYINPUT67), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(G137), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT68), .B(G131), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n219), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n211), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT71), .ZN(new_n227));
  INV_X1    g041(.A(G113), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  XOR2_X1   g047(.A(new_n232), .B(new_n233), .Z(new_n234));
  INV_X1    g048(.A(KEYINPUT0), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n189), .A3(KEYINPUT64), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(KEYINPUT0), .B2(G128), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n236), .A2(new_n238), .B1(KEYINPUT0), .B2(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n203), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT66), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n219), .B1(new_n213), .B2(KEYINPUT11), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n217), .B1(new_n216), .B2(KEYINPUT67), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n221), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n203), .A2(new_n246), .A3(new_n239), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n208), .B1(new_n202), .B2(G143), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT0), .A3(G128), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n241), .A2(new_n245), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n226), .A2(new_n227), .A3(new_n234), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n210), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n200), .B2(new_n206), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n250), .B(new_n234), .C1(new_n253), .C2(new_n224), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n234), .B1(new_n226), .B2(new_n250), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT28), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n264), .B(KEYINPUT27), .Z(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XOR2_X1   g080(.A(new_n265), .B(new_n266), .Z(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n261), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G902), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n211), .A2(KEYINPUT70), .A3(new_n225), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n253), .B2(new_n224), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .A4(new_n250), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n253), .A2(new_n224), .ZN(new_n276));
  INV_X1    g090(.A(new_n250), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT30), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n234), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n256), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n268), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n277), .B1(new_n276), .B2(KEYINPUT70), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n234), .B1(new_n284), .B2(new_n273), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT28), .B1(new_n285), .B2(new_n256), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n260), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n283), .B(new_n262), .C1(new_n268), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n187), .B1(new_n270), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n279), .A2(new_n280), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  INV_X1    g105(.A(new_n256), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n267), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n281), .A2(KEYINPUT72), .A3(new_n291), .A4(new_n267), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n267), .A3(new_n292), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n287), .A2(new_n268), .B1(new_n298), .B2(KEYINPUT31), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n187), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT32), .ZN(new_n303));
  AOI21_X1  g117(.A(G902), .B1(new_n297), .B2(new_n299), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n187), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n289), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT75), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT16), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(G125), .A2(G140), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n312), .B2(G140), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n317), .B2(new_n313), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(G146), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT24), .B(G110), .Z(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT73), .ZN(new_n321));
  XNOR2_X1  g135(.A(G119), .B(G128), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G128), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(G119), .C2(new_n189), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT74), .ZN(new_n329));
  INV_X1    g143(.A(G110), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n319), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT76), .B(G110), .Z(new_n333));
  OAI22_X1  g147(.A1(new_n321), .A2(new_n322), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G125), .B(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n202), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(G146), .B(new_n315), .C1(new_n317), .C2(new_n313), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G137), .ZN(new_n340));
  INV_X1    g154(.A(G953), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(G221), .A3(G234), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n340), .B(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n343), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n332), .B2(new_n338), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT25), .B1(new_n347), .B2(G902), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n301), .C1(new_n344), .C2(new_n346), .ZN(new_n350));
  INV_X1    g164(.A(G217), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(G234), .B2(new_n301), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(G902), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n344), .B2(new_n346), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT77), .B1(new_n307), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n289), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n304), .A2(new_n305), .A3(new_n187), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n305), .B1(new_n304), .B2(new_n187), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n362));
  INV_X1    g176(.A(new_n356), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n220), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n263), .A2(G143), .A3(G214), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G143), .B1(new_n263), .B2(G214), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n366), .B(KEYINPUT17), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n371));
  INV_X1    g185(.A(new_n369), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n220), .A3(new_n367), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n374), .A2(KEYINPUT17), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n319), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT18), .A2(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n367), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(KEYINPUT18), .B(G131), .C1(new_n368), .C2(new_n369), .ZN(new_n379));
  INV_X1    g193(.A(new_n316), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT75), .B(G125), .ZN(new_n381));
  OAI211_X1 g195(.A(G146), .B(new_n380), .C1(new_n381), .C2(new_n314), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n382), .A2(KEYINPUT89), .A3(new_n336), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT89), .B1(new_n382), .B2(new_n336), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n378), .B(new_n379), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G113), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n376), .A2(new_n385), .A3(new_n389), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n301), .B1(new_n391), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g209(.A(G475), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT81), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G116), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G122), .ZN(new_n403));
  INV_X1    g217(.A(G122), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G116), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(G107), .ZN(new_n408));
  XNOR2_X1  g222(.A(G116), .B(G122), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT93), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n189), .A2(G143), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT13), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n212), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G128), .B(G143), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n401), .A2(new_n406), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n408), .A2(new_n409), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n411), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT9), .B(G234), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT78), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n423), .A2(new_n351), .A3(G953), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT14), .B1(new_n404), .B2(G116), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(new_n402), .B2(G122), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n403), .A2(KEYINPUT14), .ZN(new_n427));
  OAI21_X1  g241(.A(G107), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n415), .A2(G134), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n415), .A2(G134), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n418), .A4(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n421), .A2(new_n424), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT94), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n421), .A2(new_n424), .A3(new_n431), .A4(KEYINPUT94), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n421), .A2(new_n431), .ZN(new_n436));
  INV_X1    g250(.A(new_n424), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n301), .ZN(new_n440));
  AND2_X1   g254(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n441));
  NOR2_X1   g255(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n442));
  OAI21_X1  g256(.A(G478), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n440), .B(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n335), .A2(KEYINPUT19), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n380), .B1(new_n381), .B2(new_n314), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n446), .B2(KEYINPUT19), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n337), .B(new_n374), .C1(new_n447), .C2(new_n198), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n385), .A2(KEYINPUT90), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n390), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT90), .B1(new_n385), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT91), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n385), .A2(new_n448), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n449), .A4(new_n390), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n452), .A2(new_n457), .A3(new_n393), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n459));
  NOR2_X1   g273(.A1(G475), .A2(G902), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n458), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n396), .B(new_n444), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(KEYINPUT96), .A2(G952), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(KEYINPUT96), .A2(G952), .ZN(new_n466));
  AOI21_X1  g280(.A(G953), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G234), .ZN(new_n468));
  INV_X1    g282(.A(G237), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G898), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n301), .B(new_n341), .C1(G234), .C2(G237), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n245), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(G104), .B2(new_n397), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n388), .A2(KEYINPUT85), .A3(G107), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G104), .B1(new_n398), .B2(new_n400), .ZN(new_n481));
  OAI21_X1  g295(.A(G101), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT82), .B1(new_n397), .B2(G104), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n388), .A3(G107), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n398), .A3(new_n400), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT83), .B(G101), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT3), .B1(new_n388), .B2(G107), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n486), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n253), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n492), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n189), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n210), .B1(new_n248), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n476), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(KEYINPUT12), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n496), .A2(new_n491), .A3(new_n482), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n253), .B2(new_n492), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT12), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n501), .A2(new_n502), .A3(new_n476), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT86), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n211), .A2(KEYINPUT10), .A3(new_n494), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n241), .A2(new_n247), .A3(new_n249), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n507));
  AND2_X1   g321(.A1(KEYINPUT84), .A2(G101), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(KEYINPUT4), .A3(new_n508), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n491), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT10), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n497), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n505), .A2(new_n514), .A3(new_n516), .A4(new_n476), .ZN(new_n517));
  XOR2_X1   g331(.A(G110), .B(G140), .Z(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT80), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n341), .A2(G227), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n498), .A2(KEYINPUT12), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n502), .B1(new_n501), .B2(new_n476), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n504), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n505), .A2(new_n514), .A3(new_n516), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n245), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n517), .ZN(new_n531));
  INV_X1    g345(.A(new_n521), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G469), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n301), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n524), .A2(new_n525), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n532), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n523), .A2(new_n530), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(G469), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n535), .A2(new_n301), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n536), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G221), .B1(new_n423), .B2(G902), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT79), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n475), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AND4_X1   g364(.A1(new_n241), .A2(new_n247), .A3(new_n249), .A4(new_n312), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n551), .B1(new_n381), .B2(new_n211), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n341), .A2(G224), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n509), .A2(new_n510), .B1(new_n556), .B2(new_n489), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n234), .B1(new_n557), .B2(new_n512), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n402), .A2(G119), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT5), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n228), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n325), .A2(G116), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n402), .A2(G119), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT5), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n561), .A2(new_n564), .B1(new_n233), .B2(new_n232), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n482), .A2(new_n491), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT87), .B1(new_n558), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT87), .ZN(new_n568));
  INV_X1    g382(.A(new_n566), .ZN(new_n569));
  INV_X1    g383(.A(new_n512), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT4), .B1(new_n507), .B2(new_n508), .ZN(new_n571));
  INV_X1    g385(.A(new_n491), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n568), .B(new_n569), .C1(new_n573), .C2(new_n234), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n555), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n555), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n558), .A2(new_n566), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT6), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n513), .A2(new_n280), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n568), .B1(new_n579), .B2(new_n569), .ZN(new_n580));
  AOI211_X1 g394(.A(KEYINPUT87), .B(new_n566), .C1(new_n513), .C2(new_n280), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n576), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT6), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n554), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n552), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n586), .A2(KEYINPUT7), .A3(new_n553), .ZN(new_n587));
  INV_X1    g401(.A(new_n577), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n553), .A2(KEYINPUT7), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n552), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n555), .B(KEYINPUT8), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n494), .A2(new_n565), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n566), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n301), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n550), .B1(new_n585), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n554), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n583), .B1(new_n582), .B2(new_n588), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n575), .A2(KEYINPUT6), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n594), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n586), .A2(KEYINPUT7), .A3(new_n553), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n603), .A3(new_n549), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n596), .A2(new_n604), .A3(KEYINPUT88), .ZN(new_n605));
  OAI21_X1  g419(.A(G214), .B1(G237), .B2(G902), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT88), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n600), .A2(new_n607), .A3(new_n603), .A4(new_n549), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n548), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n365), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n611), .B(new_n489), .Z(G3));
  XNOR2_X1  g426(.A(new_n304), .B(G472), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n544), .A2(new_n547), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n356), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT97), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n600), .A2(new_n603), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n550), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n618), .B(new_n550), .C1(new_n585), .C2(new_n595), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n604), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n606), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n585), .A2(new_n595), .A3(new_n550), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n596), .A2(KEYINPUT98), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n627), .B2(new_n621), .ZN(new_n628));
  INV_X1    g442(.A(new_n606), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT99), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n474), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n458), .A2(new_n460), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT20), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n439), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n438), .A2(KEYINPUT33), .A3(new_n432), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(G478), .A3(new_n301), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT100), .B(G478), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT101), .B1(new_n440), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n643), .B(new_n640), .C1(new_n439), .C2(new_n301), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n639), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT102), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n647), .B(new_n639), .C1(new_n642), .C2(new_n644), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n635), .A2(new_n396), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n625), .A2(new_n630), .A3(new_n631), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n617), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  INV_X1    g468(.A(new_n444), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n655), .B(new_n396), .C1(new_n461), .C2(new_n462), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n625), .A2(new_n630), .A3(new_n631), .A4(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n617), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n345), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n339), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n354), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n353), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n613), .A2(new_n610), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  AND3_X1   g483(.A1(new_n625), .A2(new_n630), .A3(new_n666), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n361), .ZN(new_n671));
  INV_X1    g485(.A(new_n473), .ZN(new_n672));
  OR3_X1    g486(.A1(new_n672), .A2(KEYINPUT103), .A3(G900), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT103), .B1(new_n672), .B2(G900), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n470), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n657), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n614), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT104), .B(G128), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G30));
  NAND2_X1  g494(.A1(new_n635), .A2(new_n396), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n444), .ZN(new_n683));
  INV_X1    g497(.A(new_n666), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n606), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT106), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n605), .A2(new_n608), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n268), .B1(new_n256), .B2(new_n257), .ZN(new_n690));
  AOI21_X1  g504(.A(G902), .B1(new_n298), .B2(new_n690), .ZN(new_n691));
  OAI22_X1  g505(.A1(new_n359), .A2(new_n360), .B1(new_n187), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT105), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n675), .B(KEYINPUT39), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n614), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT40), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n689), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NAND2_X1  g513(.A1(new_n646), .A2(new_n648), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n681), .A2(new_n700), .A3(new_n675), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n614), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n671), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  AOI21_X1  g519(.A(new_n522), .B1(new_n537), .B2(KEYINPUT86), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n706), .A2(new_n527), .B1(new_n532), .B2(new_n531), .ZN(new_n707));
  OAI21_X1  g521(.A(G469), .B1(new_n707), .B2(G902), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n536), .A3(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(KEYINPUT107), .B(G469), .C1(new_n707), .C2(G902), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n546), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n361), .A2(new_n363), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n650), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT41), .B(G113), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NOR2_X1   g530(.A1(new_n713), .A2(new_n658), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n402), .ZN(G18));
  AND4_X1   g532(.A1(new_n625), .A2(new_n630), .A3(new_n666), .A4(new_n712), .ZN(new_n719));
  INV_X1    g533(.A(new_n475), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n307), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n361), .A2(new_n475), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n625), .A2(new_n630), .A3(new_n666), .A4(new_n712), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT108), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT109), .B(G119), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G21));
  NAND3_X1  g543(.A1(new_n625), .A2(new_n630), .A3(new_n683), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n187), .A2(new_n301), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n268), .A2(new_n261), .B1(new_n298), .B2(KEYINPUT31), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n731), .B1(new_n297), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n300), .A2(new_n301), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n733), .B1(new_n734), .B2(G472), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n631), .A3(new_n712), .A4(new_n363), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n404), .ZN(G24));
  AND3_X1   g552(.A1(new_n625), .A2(new_n630), .A3(new_n712), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n666), .A3(new_n701), .A4(new_n735), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n307), .B2(new_n356), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n361), .A2(KEYINPUT111), .A3(new_n363), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n629), .B1(new_n605), .B2(new_n608), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n541), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n541), .A2(new_n746), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n536), .B(new_n543), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n745), .A2(new_n701), .A3(new_n749), .A4(new_n547), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n743), .A2(new_n744), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n745), .A2(new_n547), .A3(new_n749), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n361), .A2(new_n754), .A3(new_n363), .A4(new_n701), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n751), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  INV_X1    g572(.A(new_n676), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n361), .A2(new_n754), .A3(new_n363), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  AND2_X1   g575(.A1(new_n646), .A2(new_n648), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n681), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT43), .ZN(new_n764));
  INV_X1    g578(.A(new_n613), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n666), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT112), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  INV_X1    g584(.A(new_n536), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n539), .A2(new_n540), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT45), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n542), .B1(new_n773), .B2(G469), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n771), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(KEYINPUT46), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n547), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n695), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n745), .B(KEYINPUT113), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n769), .A2(new_n770), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  NOR2_X1   g595(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n784), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n687), .A2(new_n606), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n702), .A2(new_n788), .A3(new_n363), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n307), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n631), .B1(new_n649), .B2(new_n657), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n609), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n613), .A3(new_n615), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n795), .B(new_n667), .C1(new_n730), .C2(new_n736), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n714), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n717), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n727), .A3(new_n611), .A4(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n547), .A2(new_n745), .A3(new_n701), .A4(new_n749), .ZN(new_n800));
  INV_X1    g614(.A(new_n733), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n801), .B(new_n666), .C1(new_n187), .C2(new_n304), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT115), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n750), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n666), .A2(new_n675), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n614), .A2(new_n808), .A3(new_n463), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n361), .A2(new_n745), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n760), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n757), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n792), .B1(new_n799), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n760), .B(new_n810), .C1(new_n804), .C2(new_n806), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n756), .B2(new_n753), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n714), .A2(new_n717), .A3(new_n796), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n723), .A2(new_n726), .B1(new_n365), .B2(new_n610), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(KEYINPUT116), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n670), .B(new_n361), .C1(new_n677), .C2(new_n703), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n625), .A2(new_n630), .A3(new_n683), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n547), .A2(new_n749), .A3(new_n684), .A4(new_n675), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n692), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n740), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n819), .A2(new_n740), .A3(KEYINPUT52), .A4(new_n822), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n813), .A2(new_n818), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT54), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n471), .A2(new_n764), .A3(new_n363), .A4(new_n735), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n547), .B1(new_n710), .B2(new_n711), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n779), .B(new_n832), .C1(new_n787), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n710), .A2(new_n711), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n745), .A2(new_n835), .A3(new_n547), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n693), .A2(new_n470), .A3(new_n356), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n682), .A3(new_n762), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n832), .A2(new_n629), .A3(new_n688), .A4(new_n712), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT50), .Z(new_n840));
  NAND2_X1  g654(.A1(new_n764), .A2(new_n471), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n836), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n803), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n834), .A2(new_n838), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT51), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n815), .A2(KEYINPUT53), .A3(new_n816), .A4(new_n817), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n825), .A2(new_n826), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n828), .B2(new_n829), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n832), .A2(new_n739), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n467), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n837), .B2(new_n649), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(KEYINPUT117), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(KEYINPUT117), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n743), .A2(new_n744), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n842), .ZN(new_n858));
  XNOR2_X1  g672(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n855), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n831), .A2(new_n845), .A3(new_n851), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(G952), .A2(G953), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n835), .B(KEYINPUT49), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n546), .A2(new_n629), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n763), .A2(new_n363), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n688), .A3(new_n866), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n862), .A2(new_n863), .B1(new_n693), .B2(new_n867), .ZN(G75));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n828), .A2(new_n829), .ZN(new_n871));
  INV_X1    g685(.A(new_n848), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(G902), .ZN(new_n874));
  INV_X1    g688(.A(G210), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n598), .A2(new_n597), .A3(new_n599), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n585), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n879), .B(new_n870), .C1(new_n874), .C2(new_n875), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n341), .A2(G952), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT120), .Z(new_n884));
  AND3_X1   g698(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(G51));
  XNOR2_X1  g699(.A(new_n849), .B(KEYINPUT54), .ZN(new_n886));
  XNOR2_X1  g700(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n543), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n534), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n874), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n773), .A2(G469), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT122), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n883), .B1(new_n889), .B2(new_n893), .ZN(G54));
  NAND2_X1  g708(.A1(KEYINPUT58), .A2(G475), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT123), .Z(new_n896));
  AND3_X1   g710(.A1(new_n890), .A2(new_n458), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n458), .B1(new_n890), .B2(new_n896), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n883), .ZN(G60));
  AND2_X1   g713(.A1(new_n637), .A2(new_n638), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n831), .A2(new_n851), .ZN(new_n901));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT59), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n900), .A2(new_n903), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n884), .B1(new_n886), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(G63));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT60), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n873), .A2(new_n664), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n347), .B(KEYINPUT125), .ZN(new_n911));
  INV_X1    g725(.A(new_n909), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n849), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n913), .A3(new_n884), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n914), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT61), .B1(new_n914), .B2(KEYINPUT124), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(G66));
  NAND2_X1  g731(.A1(G224), .A2(G953), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n799), .A2(G953), .B1(new_n472), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n578), .B(new_n584), .C1(G898), .C2(new_n341), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n919), .B(new_n920), .Z(G69));
  XNOR2_X1  g735(.A(new_n279), .B(KEYINPUT126), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n447), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(G227), .Z(new_n924));
  AND3_X1   g738(.A1(new_n924), .A2(G900), .A3(G953), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n819), .A2(new_n740), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n698), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT62), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n649), .A2(new_n657), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n365), .A2(new_n696), .A3(new_n745), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n790), .A2(new_n780), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n778), .A2(new_n857), .A3(new_n820), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n790), .A2(new_n780), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n757), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n926), .A2(new_n760), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  MUX2_X1   g753(.A(new_n933), .B(new_n939), .S(new_n923), .Z(new_n940));
  AOI21_X1  g754(.A(new_n925), .B1(new_n940), .B2(new_n341), .ZN(G72));
  NOR2_X1   g755(.A1(new_n282), .A2(new_n267), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n281), .A2(new_n268), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(G472), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT63), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n883), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n938), .A2(new_n942), .B1(new_n933), .B2(new_n943), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n799), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n944), .A2(new_n946), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n949), .B1(new_n830), .B2(new_n950), .ZN(G57));
endmodule


