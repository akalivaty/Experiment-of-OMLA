//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G29gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n202), .B1(new_n209), .B2(KEYINPUT15), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(KEYINPUT15), .B2(new_n209), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(KEYINPUT15), .A3(new_n202), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT17), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT87), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n215), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(G8gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n211), .A2(new_n212), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n214), .A2(new_n222), .B1(new_n220), .B2(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(KEYINPUT18), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(KEYINPUT18), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n219), .B(new_n220), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n224), .B(KEYINPUT13), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT88), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(G197gat), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT11), .B(G169gat), .Z(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n236), .B(KEYINPUT12), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n237), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n226), .A2(new_n231), .A3(new_n239), .A4(new_n227), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  NOR2_X1   g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(KEYINPUT23), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT23), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n243), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n246), .A2(new_n243), .A3(new_n249), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n253), .B1(new_n252), .B2(KEYINPUT64), .ZN(new_n257));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT24), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n251), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT65), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n257), .A2(new_n262), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n256), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI22_X1  g068(.A1(new_n252), .A2(KEYINPUT64), .B1(new_n265), .B2(KEYINPUT65), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n265), .A2(KEYINPUT65), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT66), .B1(new_n272), .B2(new_n257), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n255), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(KEYINPUT66), .A3(new_n257), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n267), .A2(new_n268), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n256), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(KEYINPUT67), .A3(new_n255), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n281));
  INV_X1    g080(.A(G183gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT27), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT27), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  AND4_X1   g085(.A1(KEYINPUT28), .A2(new_n283), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288));
  AOI21_X1  g087(.A(G190gat), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n245), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n294), .A2(KEYINPUT26), .A3(new_n244), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n244), .A2(KEYINPUT26), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n258), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n281), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT28), .B1(new_n302), .B2(new_n289), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT69), .B(new_n298), .C1(new_n303), .C2(new_n287), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n276), .A2(new_n280), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G226gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n298), .B1(new_n303), .B2(new_n287), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT29), .B1(new_n274), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT73), .B1(new_n311), .B2(new_n308), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n293), .A2(new_n299), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n255), .B2(new_n279), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n313), .B(new_n307), .C1(new_n315), .C2(KEYINPUT29), .ZN(new_n316));
  XOR2_X1   g115(.A(G211gat), .B(G218gat), .Z(new_n317));
  OR2_X1    g116(.A1(G197gat), .A2(G204gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(KEYINPUT72), .A3(new_n322), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n317), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n317), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n309), .A2(new_n312), .A3(new_n316), .A4(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n308), .A2(KEYINPUT29), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n308), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  AND3_X1   g138(.A1(new_n332), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n332), .B2(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n332), .A2(new_n336), .ZN(new_n344));
  INV_X1    g143(.A(new_n339), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n344), .A2(KEYINPUT30), .A3(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G134gat), .ZN(new_n350));
  INV_X1    g149(.A(G113gat), .ZN(new_n351));
  INV_X1    g150(.A(G120gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT1), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(G113gat), .A2(G120gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n350), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT1), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(G113gat), .B2(G120gat), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n358), .A2(new_n354), .A3(G134gat), .ZN(new_n359));
  OAI21_X1  g158(.A(G127gat), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n349), .B(G134gat), .C1(new_n358), .C2(new_n354), .ZN(new_n361));
  INV_X1    g160(.A(G127gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(new_n355), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n361), .B(new_n362), .C1(new_n363), .C2(G134gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G148gat), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n366), .A2(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(G141gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n367), .A2(new_n368), .B1(KEYINPUT2), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT75), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n376));
  INV_X1    g175(.A(G155gat), .ZN(new_n377));
  INV_X1    g176(.A(G162gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n371), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n369), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n370), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n378), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n370), .A2(new_n369), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n365), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n370), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n381), .B1(new_n380), .B2(new_n369), .ZN(new_n391));
  AND2_X1   g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392));
  AOI211_X1 g191(.A(KEYINPUT75), .B(new_n392), .C1(new_n379), .C2(new_n371), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n385), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT76), .A3(new_n365), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n383), .A2(new_n386), .ZN(new_n397));
  INV_X1    g196(.A(new_n365), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n389), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n348), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n404), .A3(new_n396), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(KEYINPUT3), .A3(new_n385), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n406), .A2(new_n398), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n394), .B2(new_n385), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n394), .A2(new_n385), .B1(new_n360), .B2(new_n364), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n402), .B1(new_n411), .B2(KEYINPUT4), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n405), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n403), .A2(new_n413), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n407), .A2(new_n409), .B1(new_n404), .B2(new_n387), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n395), .A2(KEYINPUT76), .A3(new_n365), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT76), .B1(new_n395), .B2(new_n365), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT4), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n415), .A2(new_n418), .A3(new_n348), .A4(new_n401), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT78), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n426), .A3(new_n419), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n347), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT35), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n306), .A2(new_n365), .ZN(new_n438));
  INV_X1    g237(.A(G227gat), .ZN(new_n439));
  INV_X1    g238(.A(G233gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n276), .A2(new_n305), .A3(new_n398), .A4(new_n280), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G71gat), .B(G99gat), .Z(new_n444));
  XNOR2_X1  g243(.A(G15gat), .B(G43gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT33), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(KEYINPUT32), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT71), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT71), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n443), .A2(new_n450), .A3(KEYINPUT32), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n443), .A2(KEYINPUT32), .ZN(new_n453));
  INV_X1    g252(.A(new_n443), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n453), .B(new_n446), .C1(new_n454), .C2(KEYINPUT33), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n441), .B1(new_n438), .B2(new_n442), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT34), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n452), .B2(new_n455), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT81), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n330), .B1(new_n408), .B2(KEYINPUT29), .ZN(new_n462));
  INV_X1    g261(.A(new_n317), .ZN(new_n463));
  AOI211_X1 g262(.A(new_n324), .B(new_n321), .C1(new_n318), .C2(new_n319), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT72), .B1(new_n320), .B2(new_n322), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT29), .B1(new_n466), .B2(new_n328), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n397), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g267(.A1(G228gat), .A2(G233gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n462), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT3), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n467), .B2(KEYINPUT79), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT29), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT79), .B(new_n475), .C1(new_n327), .C2(new_n329), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n397), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT80), .B(new_n330), .C1(new_n408), .C2(KEYINPUT29), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n472), .B1(new_n482), .B2(new_n469), .ZN(new_n483));
  INV_X1    g282(.A(G22gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n461), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G78gat), .B(G106gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G50gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n483), .A2(new_n484), .ZN(new_n490));
  AOI211_X1 g289(.A(G22gat), .B(new_n472), .C1(new_n482), .C2(new_n469), .ZN(new_n491));
  OAI22_X1  g290(.A1(new_n485), .A2(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n482), .A2(new_n469), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n471), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G22gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n483), .A2(new_n484), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n495), .A2(new_n461), .A3(new_n496), .A4(new_n488), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n437), .B1(new_n460), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n452), .A2(new_n455), .ZN(new_n500));
  INV_X1    g299(.A(new_n457), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n503));
  AND4_X1   g302(.A1(new_n437), .A2(new_n502), .A3(new_n498), .A4(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n436), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT39), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n404), .B1(new_n389), .B2(new_n396), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n406), .A2(new_n398), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n508), .A2(new_n408), .B1(KEYINPUT4), .B2(new_n411), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n506), .B(new_n402), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n401), .B1(new_n415), .B2(new_n418), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT39), .B1(new_n400), .B2(new_n402), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n426), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT40), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n426), .B1(new_n414), .B2(new_n419), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n343), .A2(new_n346), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n519), .A2(new_n520), .B1(new_n497), .B2(new_n492), .ZN(new_n521));
  INV_X1    g320(.A(new_n340), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n431), .A2(new_n432), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n345), .B1(new_n344), .B2(KEYINPUT37), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(new_n332), .B2(new_n336), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT38), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n344), .A2(new_n345), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n345), .A2(KEYINPUT37), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT38), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n309), .A2(new_n316), .A3(new_n312), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT83), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n531), .A2(new_n532), .A3(new_n330), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n531), .B2(new_n330), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n530), .B1(new_n536), .B2(new_n525), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n523), .A2(new_n527), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n458), .B2(new_n459), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n498), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n434), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n460), .A2(new_n498), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n435), .B1(new_n547), .B2(new_n434), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n505), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT85), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n505), .A2(new_n546), .A3(KEYINPUT85), .A4(new_n548), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n242), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  INV_X1    g357(.A(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G127gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n558), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n219), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n377), .ZN(new_n568));
  XOR2_X1   g367(.A(G183gat), .B(G211gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n570), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n575));
  OAI211_X1 g374(.A(G85gat), .B(G92gat), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n575), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(KEYINPUT90), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(KEYINPUT90), .B2(new_n580), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT91), .B(G92gat), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n578), .B(new_n582), .C1(G85gat), .C2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G99gat), .B(G106gat), .Z(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n589), .A2(new_n220), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n220), .A2(new_n221), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n214), .A2(new_n592), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT92), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n558), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n564), .A3(new_n587), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n606), .A2(new_n608), .ZN(new_n615));
  INV_X1    g414(.A(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G120gat), .B(G148gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT95), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n616), .B1(new_n609), .B2(new_n610), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n614), .A2(new_n617), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n613), .A2(new_n617), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n621), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n573), .A2(new_n605), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n553), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(new_n433), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(G1gat), .Z(G1324gat));
  OAI21_X1  g434(.A(G8gat), .B1(new_n633), .B2(new_n347), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT16), .B(G8gat), .Z(new_n639));
  NAND4_X1  g438(.A1(new_n553), .A2(new_n520), .A3(new_n632), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT42), .B1(new_n640), .B2(KEYINPUT96), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n640), .A2(KEYINPUT96), .A3(KEYINPUT42), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n637), .B(new_n638), .C1(new_n641), .C2(new_n642), .ZN(G1325gat));
  OAI21_X1  g442(.A(G15gat), .B1(new_n633), .B2(new_n543), .ZN(new_n644));
  INV_X1    g443(.A(new_n460), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n645), .A2(G15gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n633), .B2(new_n646), .ZN(G1326gat));
  NOR2_X1   g446(.A1(new_n633), .A2(new_n498), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT43), .B(G22gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(G1327gat));
  INV_X1    g449(.A(new_n605), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n573), .A2(new_n629), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n553), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n653), .A2(G29gat), .A3(new_n433), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT98), .B(KEYINPUT45), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(KEYINPUT44), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n551), .B2(new_n552), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n549), .B2(new_n651), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n573), .A2(new_n242), .A3(new_n629), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(G29gat), .B1(new_n662), .B2(new_n433), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n656), .A2(new_n663), .ZN(G1328gat));
  NOR3_X1   g463(.A1(new_n653), .A2(G36gat), .A3(new_n347), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT46), .ZN(new_n666));
  OAI21_X1  g465(.A(G36gat), .B1(new_n662), .B2(new_n347), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(G1329gat));
  OAI21_X1  g467(.A(G43gat), .B1(new_n662), .B2(new_n543), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT47), .B1(new_n669), .B2(KEYINPUT99), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n653), .A2(G43gat), .A3(new_n645), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n670), .B(new_n672), .ZN(G1330gat));
  NAND3_X1  g472(.A1(new_n660), .A2(new_n544), .A3(new_n661), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G50gat), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n498), .A2(G50gat), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n653), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT100), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g478(.A(new_n573), .ZN(new_n680));
  NOR4_X1   g479(.A1(new_n680), .A2(new_n651), .A3(new_n241), .A4(new_n630), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n549), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n433), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT101), .B(G57gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1332gat));
  AOI21_X1  g485(.A(new_n347), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT102), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1333gat));
  INV_X1    g490(.A(new_n543), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n682), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n645), .A2(G71gat), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n693), .A2(G71gat), .B1(new_n682), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g495(.A1(new_n682), .A2(new_n544), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT103), .B(G78gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1335gat));
  NOR2_X1   g498(.A1(new_n573), .A2(new_n241), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n549), .A2(KEYINPUT51), .A3(new_n651), .A4(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n549), .A2(new_n651), .A3(new_n700), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT51), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n703), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n433), .A2(G85gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n629), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n629), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n660), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G85gat), .B1(new_n712), .B2(new_n433), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(G1336gat));
  NOR4_X1   g513(.A1(new_n658), .A2(new_n347), .A3(new_n659), .A4(new_n710), .ZN(new_n715));
  INV_X1    g514(.A(new_n583), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n706), .A2(new_n701), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n347), .A2(G92gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n629), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT52), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n715), .B2(new_n716), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n707), .A2(KEYINPUT105), .A3(new_n629), .A4(new_n719), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n706), .A2(new_n702), .A3(new_n701), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n704), .A2(KEYINPUT104), .A3(new_n705), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n727), .A2(new_n629), .A3(new_n728), .A4(new_n719), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n723), .B(new_n725), .C1(new_n726), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n726), .A2(new_n731), .ZN(new_n733));
  INV_X1    g532(.A(new_n725), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT106), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n722), .B1(new_n732), .B2(new_n735), .ZN(G1337gat));
  NOR2_X1   g535(.A1(new_n645), .A2(G99gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n707), .A2(new_n629), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G99gat), .B1(new_n712), .B2(new_n543), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1338gat));
  NOR3_X1   g539(.A1(new_n630), .A2(new_n498), .A3(G106gat), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT53), .B1(new_n707), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n660), .A2(new_n544), .A3(new_n711), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G106gat), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(KEYINPUT107), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n706), .A2(new_n701), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n743), .A2(G106gat), .B1(new_n749), .B2(new_n741), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(G1339gat));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n632), .A2(new_n752), .A3(new_n242), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT108), .B1(new_n631), .B2(new_n241), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n223), .A2(new_n224), .B1(new_n228), .B2(new_n229), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n236), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n240), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n605), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n622), .B1(new_n623), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n614), .A2(KEYINPUT54), .A3(new_n625), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n609), .A2(new_n610), .A3(new_n616), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(KEYINPUT55), .B(new_n761), .C1(new_n762), .C2(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n766), .A2(new_n626), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n761), .B1(new_n762), .B2(new_n765), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n759), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n758), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n629), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n630), .A2(new_n758), .A3(KEYINPUT110), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n770), .A2(new_n241), .A3(new_n626), .A4(new_n766), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n771), .B1(new_n777), .B2(new_n605), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n755), .B1(new_n778), .B2(new_n573), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n498), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n780), .A2(KEYINPUT111), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n645), .B1(new_n780), .B2(KEYINPUT111), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n520), .A2(new_n433), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(G113gat), .A3(new_n241), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n779), .A2(new_n683), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n499), .A2(new_n504), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n347), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n351), .B1(new_n790), .B2(new_n242), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n786), .A2(new_n791), .ZN(G1340gat));
  NAND3_X1  g591(.A1(new_n785), .A2(G120gat), .A3(new_n629), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n352), .B1(new_n790), .B2(new_n630), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(G1341gat));
  XOR2_X1   g594(.A(KEYINPUT70), .B(G127gat), .Z(new_n796));
  NAND2_X1  g595(.A1(new_n783), .A2(new_n784), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n680), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n680), .A2(new_n796), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n790), .B2(new_n799), .ZN(G1342gat));
  NAND2_X1  g599(.A1(new_n787), .A2(new_n789), .ZN(new_n801));
  NOR4_X1   g600(.A1(new_n801), .A2(G134gat), .A3(new_n520), .A4(new_n605), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT56), .ZN(new_n803));
  OAI21_X1  g602(.A(G134gat), .B1(new_n797), .B2(new_n605), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1343gat));
  NOR2_X1   g604(.A1(new_n692), .A2(new_n498), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n520), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n242), .A2(G141gat), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n543), .A2(new_n784), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT112), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  INV_X1    g612(.A(new_n771), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n241), .A2(new_n626), .A3(new_n766), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n768), .A2(KEYINPUT113), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n817), .B(new_n761), .C1(new_n762), .C2(new_n765), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n769), .A3(new_n818), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n815), .A2(new_n819), .B1(new_n629), .B2(new_n772), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n820), .B2(new_n651), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n680), .ZN(new_n822));
  AOI211_X1 g621(.A(new_n813), .B(new_n498), .C1(new_n822), .C2(new_n755), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT57), .B1(new_n779), .B2(new_n544), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n241), .B(new_n812), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n808), .A2(new_n809), .B1(new_n825), .B2(G141gat), .ZN(new_n826));
  XOR2_X1   g625(.A(KEYINPUT114), .B(KEYINPUT58), .Z(new_n827));
  XNOR2_X1  g626(.A(new_n826), .B(new_n827), .ZN(G1344gat));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n812), .B1(new_n823), .B2(new_n824), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n829), .B(G148gat), .C1(new_n830), .C2(new_n630), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n779), .A2(new_n544), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n811), .A2(new_n630), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n573), .B1(new_n821), .B2(KEYINPUT115), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n814), .B(new_n837), .C1(new_n820), .C2(new_n651), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n836), .A2(new_n838), .B1(new_n242), .B2(new_n632), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n498), .A2(KEYINPUT57), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n834), .B(new_n835), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G148gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n832), .B1(new_n843), .B2(KEYINPUT59), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT116), .B(new_n829), .C1(new_n842), .C2(G148gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n831), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n808), .A2(new_n366), .A3(new_n629), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1345gat));
  OAI21_X1  g647(.A(G155gat), .B1(new_n830), .B2(new_n680), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n808), .A2(new_n377), .A3(new_n573), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1346gat));
  OAI21_X1  g650(.A(G162gat), .B1(new_n830), .B2(new_n605), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n651), .A2(new_n378), .A3(new_n347), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n807), .B2(new_n853), .ZN(G1347gat));
  NOR2_X1   g653(.A1(new_n347), .A2(new_n683), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n783), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n247), .A3(new_n242), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n779), .A2(new_n433), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n788), .A2(new_n347), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(G169gat), .B1(new_n860), .B2(new_n241), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n857), .A2(new_n861), .ZN(G1348gat));
  OAI21_X1  g661(.A(G176gat), .B1(new_n856), .B2(new_n630), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n860), .A2(new_n248), .A3(new_n629), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1349gat));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n680), .A2(new_n301), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n858), .A2(new_n859), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n859), .A4(new_n868), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n781), .A2(new_n782), .A3(new_n573), .A4(new_n855), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G183gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n873), .B2(new_n875), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1350gat));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n286), .A3(new_n651), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT119), .Z(new_n881));
  NAND4_X1  g680(.A1(new_n781), .A2(new_n782), .A3(new_n651), .A4(new_n855), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G190gat), .ZN(new_n883));
  XNOR2_X1  g682(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(G1351gat));
  AND3_X1   g686(.A1(new_n858), .A2(new_n520), .A3(new_n806), .ZN(new_n888));
  AOI21_X1  g687(.A(G197gat), .B1(new_n888), .B2(new_n241), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n543), .A2(new_n855), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT122), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n834), .B1(new_n839), .B2(new_n841), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT121), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n813), .B1(new_n779), .B2(new_n544), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n816), .A2(new_n769), .A3(new_n818), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n241), .A2(new_n626), .A3(new_n766), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n773), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n771), .B1(new_n897), .B2(new_n605), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n680), .B1(new_n898), .B2(new_n837), .ZN(new_n899));
  INV_X1    g698(.A(new_n838), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n899), .A2(new_n900), .B1(new_n241), .B2(new_n631), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n894), .B1(new_n901), .B2(new_n840), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n891), .B1(new_n893), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n241), .A2(G197gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n889), .B1(new_n905), .B2(new_n906), .ZN(G1352gat));
  NOR2_X1   g706(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n908));
  XOR2_X1   g707(.A(KEYINPUT123), .B(G204gat), .Z(new_n909));
  AND2_X1   g708(.A1(new_n629), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n888), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(new_n913));
  AOI211_X1 g712(.A(new_n630), .B(new_n891), .C1(new_n893), .C2(new_n904), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n909), .ZN(G1353gat));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916));
  INV_X1    g715(.A(G211gat), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n890), .A2(new_n680), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n902), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n919), .B2(KEYINPUT63), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n921), .A3(KEYINPUT63), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n834), .B(new_n918), .C1(new_n839), .C2(new_n841), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT125), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(G211gat), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(KEYINPUT126), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n920), .A2(new_n922), .A3(new_n925), .A4(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n888), .A2(new_n917), .A3(new_n573), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1354gat));
  AOI21_X1  g730(.A(G218gat), .B1(new_n888), .B2(new_n651), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n651), .A2(G218gat), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT127), .Z(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n905), .B2(new_n934), .ZN(G1355gat));
endmodule


