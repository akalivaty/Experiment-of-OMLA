//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G137), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n463), .A2(new_n466), .ZN(G160));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n460), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n459), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n459), .A2(G102), .A3(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n460), .B2(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n486), .B1(new_n489), .B2(new_n459), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(new_n469), .A3(new_n471), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n485), .B1(new_n490), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n486), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n487), .B1(new_n472), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT4), .B1(new_n460), .B2(new_n492), .ZN(new_n503));
  AND4_X1   g078(.A1(KEYINPUT4), .A2(new_n492), .A3(new_n469), .A4(new_n471), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(KEYINPUT68), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n498), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT70), .B(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(KEYINPUT70), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n512), .B(KEYINPUT5), .C1(new_n514), .C2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(G543), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n511), .A2(G62), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n508), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n511), .A2(new_n520), .A3(new_n517), .A4(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(G50), .A3(G543), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT69), .ZN(new_n529));
  NOR3_X1   g104(.A1(new_n523), .A2(new_n527), .A3(new_n529), .ZN(G166));
  NAND2_X1  g105(.A1(new_n524), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n511), .A2(new_n520), .A3(new_n517), .ZN(new_n534));
  NAND2_X1  g109(.A1(G63), .A2(G651), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n525), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT73), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n534), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n532), .A2(G52), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n525), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n534), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n556), .ZN(new_n558));
  NOR3_X1   g133(.A1(new_n557), .A2(new_n558), .A3(new_n508), .ZN(new_n559));
  INV_X1    g134(.A(new_n525), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G81), .B1(G43), .B2(new_n532), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT75), .Z(G188));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n534), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n560), .A2(G91), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n532), .A2(KEYINPUT9), .A3(G53), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n531), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n574), .A2(new_n575), .A3(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  INV_X1    g157(.A(G166), .ZN(G303));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n534), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n560), .A2(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n532), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND4_X1  g164(.A1(new_n511), .A2(G61), .A3(new_n517), .A4(new_n520), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n560), .A2(G86), .B1(G48), .B2(new_n532), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n592), .A2(KEYINPUT76), .A3(G651), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n532), .A2(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n525), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT77), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n534), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n525), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  INV_X1    g187(.A(G79), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n534), .A2(new_n612), .B1(new_n613), .B2(new_n515), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT78), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n616));
  OAI221_X1 g191(.A(new_n616), .B1(new_n613), .B2(new_n515), .C1(new_n534), .C2(new_n612), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n615), .A2(G651), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n532), .A2(G54), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n611), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n608), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n608), .B1(new_n621), .B2(G868), .ZN(G321));
  INV_X1    g198(.A(G299), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT79), .B1(new_n624), .B2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  MUX2_X1   g201(.A(KEYINPUT79), .B(new_n625), .S(new_n626), .Z(G297));
  MUX2_X1   g202(.A(KEYINPUT79), .B(new_n625), .S(new_n626), .Z(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n621), .B1(new_n629), .B2(G860), .ZN(G148));
  OR3_X1    g205(.A1(new_n557), .A2(new_n558), .A3(new_n508), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n561), .ZN(new_n632));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n620), .A2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n477), .A2(G123), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n479), .A2(G135), .ZN(new_n640));
  NOR2_X1   g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(new_n459), .B2(G111), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  INV_X1    g222(.A(G2100), .ZN(new_n648));
  OR3_X1    g223(.A1(new_n647), .A2(KEYINPUT81), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n647), .B1(KEYINPUT81), .B2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(KEYINPUT81), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n644), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2435), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2438), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(G14), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  XOR2_X1   g246(.A(new_n668), .B(KEYINPUT82), .Z(new_n672));
  OAI21_X1  g247(.A(KEYINPUT17), .B1(new_n672), .B2(new_n667), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(new_n669), .Z(new_n674));
  AND2_X1   g249(.A1(new_n672), .A2(new_n667), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT83), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(new_n648), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AOI21_X1  g258(.A(KEYINPUT84), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g259(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT84), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n686), .A2(new_n687), .B1(new_n681), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n682), .B(new_n683), .ZN(new_n690));
  OAI221_X1 g265(.A(new_n689), .B1(new_n687), .B2(new_n686), .C1(new_n681), .C2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT22), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  NAND4_X1  g272(.A1(new_n473), .A2(new_n475), .A3(G141), .A4(new_n459), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n473), .A2(new_n475), .A3(G129), .A4(G2105), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT26), .Z(new_n702));
  NAND4_X1  g277(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G32), .B(new_n703), .S(G29), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT27), .B(G1996), .Z(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  INV_X1    g281(.A(G34), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(KEYINPUT24), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(KEYINPUT24), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G160), .B2(new_n706), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G2084), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n704), .A2(new_n705), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G5), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G171), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT94), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n714), .B1(new_n718), .B2(G1961), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT95), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n715), .A2(KEYINPUT23), .A3(G20), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n722));
  INV_X1    g297(.A(G20), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G16), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n721), .B(new_n724), .C1(new_n624), .C2(new_n715), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1956), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G1961), .B2(new_n718), .ZN(new_n727));
  NOR2_X1   g302(.A1(G27), .A2(G29), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G164), .B2(G29), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT97), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT96), .B(G2078), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n706), .A2(G26), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n477), .A2(G128), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n479), .A2(G140), .ZN(new_n736));
  OR2_X1    g311(.A1(G104), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n733), .B(new_n734), .C1(new_n739), .C2(G29), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n733), .B2(new_n734), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT90), .B(G2067), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n720), .A2(new_n727), .A3(new_n732), .A4(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n563), .A2(new_n715), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n715), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(KEYINPUT89), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT89), .B2(new_n746), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1341), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n730), .A2(new_n731), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n715), .A2(G4), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n621), .B2(new_n715), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1348), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n744), .A2(new_n749), .A3(new_n750), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n715), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n715), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n759));
  NOR2_X1   g334(.A1(G6), .A2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G305), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT32), .B(G1981), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT87), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n762), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n715), .A2(G22), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G166), .B2(new_n715), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(G1971), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(G1971), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT88), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G23), .ZN(new_n771));
  OR3_X1    g346(.A1(new_n770), .A2(G16), .A3(G23), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n771), .B(new_n772), .C1(G288), .C2(new_n715), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT33), .B(G1976), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n765), .A2(new_n768), .A3(new_n769), .A4(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT34), .Z(new_n777));
  INV_X1    g352(.A(new_n479), .ZN(new_n778));
  INV_X1    g353(.A(G131), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n778), .A2(KEYINPUT86), .A3(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(G95), .A2(G2105), .ZN(new_n781));
  INV_X1    g356(.A(G107), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n468), .B1(new_n782), .B2(G2105), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n477), .A2(G119), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT86), .B1(new_n778), .B2(new_n779), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n780), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT85), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n706), .A2(G25), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n786), .A2(G29), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n787), .B2(new_n788), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT35), .B(G1991), .Z(new_n791));
  XOR2_X1   g366(.A(new_n790), .B(new_n791), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n715), .A2(G24), .ZN(new_n793));
  INV_X1    g368(.A(G290), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n715), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1986), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n759), .B1(new_n777), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n777), .A2(new_n759), .A3(new_n797), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n754), .B(new_n758), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n706), .A2(G35), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G162), .B2(new_n706), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT29), .Z(new_n803));
  NOR2_X1   g378(.A1(KEYINPUT98), .A2(G2090), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT98), .A2(G2090), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n805), .B(new_n806), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT30), .B(G28), .ZN(new_n808));
  OR2_X1    g383(.A1(KEYINPUT31), .A2(G11), .ZN(new_n809));
  NAND2_X1  g384(.A1(KEYINPUT31), .A2(G11), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n808), .A2(new_n706), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n643), .B2(new_n706), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT93), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT91), .B1(G29), .B2(G33), .ZN(new_n814));
  OR3_X1    g389(.A1(KEYINPUT91), .A2(G29), .A3(G33), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n479), .A2(G139), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(new_n459), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT25), .Z(new_n820));
  NAND3_X1  g395(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n814), .B(new_n815), .C1(new_n821), .C2(new_n706), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2072), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n823), .B1(new_n713), .B2(new_n712), .C1(new_n704), .C2(new_n705), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT92), .Z(new_n825));
  NOR4_X1   g400(.A1(new_n800), .A2(new_n807), .A3(new_n813), .A4(new_n825), .ZN(G311));
  NOR2_X1   g401(.A1(new_n800), .A2(new_n825), .ZN(new_n827));
  INV_X1    g402(.A(new_n807), .ZN(new_n828));
  INV_X1    g403(.A(new_n813), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G150));
  AOI22_X1  g405(.A1(new_n560), .A2(G93), .B1(G55), .B2(new_n532), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n534), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G651), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n831), .A2(new_n835), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT99), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(G860), .A3(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n632), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n559), .A2(new_n562), .A3(new_n836), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT39), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n621), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n848), .B(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n842), .B1(new_n851), .B2(G860), .ZN(G145));
  NAND2_X1  g427(.A1(new_n479), .A2(G142), .ZN(new_n853));
  NOR2_X1   g428(.A1(G106), .A2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G130), .B2(new_n477), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n646), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n786), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n495), .A2(new_n862), .A3(new_n496), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n495), .B2(new_n496), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n502), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n703), .ZN(new_n866));
  INV_X1    g441(.A(new_n739), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT100), .B1(new_n503), .B2(new_n504), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n495), .A2(new_n496), .A3(new_n862), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n490), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n703), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(new_n739), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT101), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n866), .A2(new_n867), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n739), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n821), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n868), .A2(new_n873), .A3(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n861), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n821), .B1(new_n874), .B2(new_n878), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(KEYINPUT102), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n860), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT102), .B1(new_n885), .B2(new_n882), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n888), .B(new_n859), .C1(KEYINPUT102), .C2(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n643), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(new_n894), .A3(new_n889), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n887), .A2(KEYINPUT103), .A3(new_n889), .A4(new_n894), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g475(.A(G290), .B(KEYINPUT106), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G288), .ZN(new_n903));
  NAND2_X1  g478(.A1(G303), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G166), .A2(G288), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n904), .A2(G305), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G305), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n620), .A2(new_n624), .A3(KEYINPUT104), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n620), .B2(new_n624), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n621), .A2(G299), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT41), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT105), .B1(new_n913), .B2(new_n914), .ZN(new_n918));
  INV_X1    g493(.A(new_n914), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n912), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n918), .A2(new_n921), .B1(G299), .B2(new_n621), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n922), .B2(KEYINPUT41), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n847), .A2(new_n635), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n847), .A2(new_n635), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n915), .A2(new_n916), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n928), .B2(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n911), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  INV_X1    g511(.A(new_n911), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n932), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G868), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n843), .A2(G868), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n633), .B1(new_n935), .B2(new_n938), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n945), .B2(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(G295));
  NAND2_X1  g522(.A1(new_n940), .A2(new_n943), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(G301), .A2(G168), .ZN(new_n950));
  NAND2_X1  g525(.A1(G171), .A2(G286), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n847), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n844), .A2(new_n846), .A3(new_n951), .A4(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n917), .B(new_n955), .C1(new_n922), .C2(KEYINPUT41), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n561), .A2(new_n631), .B1(new_n838), .B2(new_n840), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n957), .A2(new_n952), .A3(new_n845), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n844), .A2(new_n846), .B1(new_n951), .B2(new_n950), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n915), .A3(new_n916), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n911), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(G37), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n956), .A2(new_n911), .A3(new_n961), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT41), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n922), .A2(new_n960), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n953), .B2(new_n954), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n911), .B1(new_n971), .B2(new_n930), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n963), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n949), .B1(new_n968), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n967), .B1(new_n963), .B2(new_n964), .ZN(new_n978));
  NOR4_X1   g553(.A1(new_n962), .A2(new_n973), .A3(G37), .A4(new_n966), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n949), .B2(new_n980), .ZN(G397));
  INV_X1    g556(.A(KEYINPUT125), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n871), .B2(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n461), .A2(new_n462), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G2105), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n464), .A2(new_n465), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n459), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT109), .B(G40), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n786), .B(new_n791), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT110), .Z(new_n995));
  INV_X1    g570(.A(G2067), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n867), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n739), .A2(G2067), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n703), .A2(G1996), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n703), .A2(G1996), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(G290), .A2(G1986), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G290), .A2(G1986), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n993), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n871), .A2(new_n991), .A3(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT112), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n463), .A2(new_n466), .A3(new_n989), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n865), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G305), .A2(G1981), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n595), .A2(new_n1018), .A3(new_n596), .A4(new_n597), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1015), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1024), .A2(new_n903), .B1(new_n1018), .B2(new_n761), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1015), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(G303), .B2(G8), .ZN(new_n1028));
  NOR3_X1   g603(.A1(G166), .A2(KEYINPUT55), .A3(new_n1008), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n865), .A2(KEYINPUT45), .A3(new_n1010), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n869), .A2(new_n870), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n1034), .B2(new_n502), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n498), .A2(new_n506), .A3(new_n1010), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n991), .B1(new_n1038), .B2(new_n983), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1971), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n991), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(G2090), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1030), .B(G8), .C1(new_n1040), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n903), .A2(G1976), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1012), .A2(new_n1013), .A3(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1013), .B1(new_n1012), .B2(G8), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1047), .B(new_n1048), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G288), .A2(new_n1023), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1022), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1025), .A2(new_n1026), .B1(new_n1046), .B2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1056), .A2(new_n1022), .A3(new_n1046), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT50), .B1(new_n871), .B2(G1384), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n498), .A2(new_n506), .A3(new_n1041), .A4(new_n1010), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1011), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(G2090), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(new_n1040), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT111), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1066));
  NOR4_X1   g641(.A1(new_n871), .A2(new_n1032), .A3(new_n983), .A4(G1384), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1039), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1971), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1064), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(KEYINPUT113), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1065), .A2(new_n1072), .A3(G8), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1030), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n498), .A2(new_n506), .A3(KEYINPUT45), .A4(new_n1010), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n984), .A2(new_n1011), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n757), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1042), .A2(new_n713), .A3(new_n1043), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(G168), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1080), .A2(new_n1081), .A3(G8), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G286), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(G8), .A3(new_n1080), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1085), .B2(KEYINPUT51), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1059), .B(new_n1075), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1068), .B2(G2078), .ZN(new_n1090));
  INV_X1    g665(.A(G1961), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1044), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1089), .A2(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n984), .A2(new_n1076), .A3(new_n1011), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G171), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1080), .A2(G8), .ZN(new_n1098));
  AOI21_X1  g673(.A(G168), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT51), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1080), .A2(new_n1081), .A3(G8), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1097), .B1(new_n1102), .B2(KEYINPUT62), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT123), .B1(new_n1088), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1096), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1056), .A2(new_n1022), .A3(new_n1046), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1074), .B2(new_n1073), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1058), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1098), .A2(G286), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1059), .A2(new_n1075), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1059), .A2(new_n1075), .A3(KEYINPUT114), .A4(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1116), .B1(new_n1119), .B2(new_n1074), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1059), .A2(new_n1112), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1111), .A2(new_n1122), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1095), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n984), .A2(G40), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1037), .A2(G160), .A3(new_n1093), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1090), .B(new_n1092), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1128), .B2(G171), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT122), .B1(new_n1095), .B2(G171), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1124), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1096), .B1(new_n1128), .B2(G171), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1125), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(new_n1107), .A3(new_n1133), .A4(new_n1102), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT57), .B1(new_n580), .B2(KEYINPUT117), .ZN(new_n1136));
  XNOR2_X1  g711(.A(G299), .B(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT115), .B(G1956), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1063), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1063), .A2(KEYINPUT116), .A3(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT56), .B(G2072), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1037), .A2(new_n1039), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1137), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1063), .A2(KEYINPUT116), .A3(new_n1138), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT116), .B1(new_n1063), .B2(new_n1138), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1137), .B(new_n1145), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT61), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1137), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(new_n1149), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT58), .B(G1341), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n1012), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1068), .B2(G1996), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT120), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1163), .B(new_n1160), .C1(new_n1068), .C2(G1996), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n563), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1162), .A2(new_n1167), .A3(new_n563), .A4(new_n1164), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1157), .A2(new_n1158), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1158), .B1(new_n1157), .B2(new_n1169), .ZN(new_n1171));
  INV_X1    g746(.A(G1348), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1044), .A2(new_n1172), .B1(new_n996), .B2(new_n1007), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT118), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n621), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(KEYINPUT60), .A3(new_n620), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1170), .A2(new_n1171), .A3(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1175), .A2(KEYINPUT119), .A3(new_n620), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT119), .B1(new_n1175), .B2(new_n620), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1150), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1135), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1006), .B1(new_n1123), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1003), .A2(new_n993), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT48), .Z(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(new_n1002), .B2(new_n993), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT46), .ZN(new_n1191));
  OR3_X1    g766(.A1(new_n993), .A2(new_n1191), .A3(G1996), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n997), .A2(new_n998), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n992), .B1(new_n1193), .B2(new_n703), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1191), .B1(new_n993), .B2(G1996), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1192), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT47), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n780), .A2(new_n791), .A3(new_n784), .A4(new_n785), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n997), .B1(new_n1001), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n992), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1190), .A2(new_n1197), .A3(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT124), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n982), .B1(new_n1187), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1180), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1157), .A2(new_n1169), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(KEYINPUT121), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1157), .A2(new_n1169), .A3(new_n1158), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1149), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1134), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1111), .A2(new_n1122), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g789(.A(KEYINPUT125), .B(new_n1202), .C1(new_n1214), .C2(new_n1006), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1204), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1218));
  NAND3_X1  g792(.A1(new_n963), .A2(new_n974), .A3(new_n967), .ZN(new_n1219));
  OAI21_X1  g793(.A(new_n1219), .B1(new_n965), .B2(new_n967), .ZN(new_n1220));
  OAI21_X1  g794(.A(G319), .B1(new_n664), .B2(new_n665), .ZN(new_n1221));
  NOR3_X1   g795(.A1(G229), .A2(new_n1221), .A3(G227), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n899), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g797(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1218), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  NOR3_X1   g799(.A1(new_n980), .A2(KEYINPUT126), .A3(new_n1223), .ZN(new_n1226));
  NOR2_X1   g800(.A1(new_n1225), .A2(new_n1226), .ZN(G308));
  NAND3_X1  g801(.A1(new_n1220), .A2(new_n1224), .A3(new_n1218), .ZN(new_n1228));
  OAI21_X1  g802(.A(KEYINPUT126), .B1(new_n980), .B2(new_n1223), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1229), .ZN(G225));
endmodule


