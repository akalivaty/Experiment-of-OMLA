//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  INV_X1    g0043(.A(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT64), .B(G50), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n244), .A2(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT68), .A2(G58), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n254), .B(KEYINPUT8), .C1(KEYINPUT67), .C2(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n255), .A2(KEYINPUT8), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n253), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n216), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G13), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n266), .A2(new_n207), .A3(G1), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G50), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n264), .B1(new_n206), .B2(G20), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(G50), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT9), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT66), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n259), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT66), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G223), .A3(G1698), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n284), .B(new_n285), .C1(new_n226), .C2(new_n282), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(new_n288), .A3(G274), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT65), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n288), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n296), .B1(new_n288), .B2(new_n297), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n295), .B1(new_n301), .B2(G226), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n290), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G200), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n290), .A2(G190), .A3(new_n302), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n273), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n273), .A2(new_n304), .A3(new_n308), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n270), .A2(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT8), .B(G58), .ZN(new_n312));
  INV_X1    g0112(.A(new_n252), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n312), .A2(new_n313), .B1(new_n207), .B2(new_n226), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n315), .B(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n317), .B2(new_n260), .ZN(new_n318));
  INV_X1    g0118(.A(new_n264), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n311), .B1(G77), .B2(new_n268), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n294), .B1(new_n300), .B2(new_n227), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n282), .A2(KEYINPUT69), .A3(G232), .A4(new_n283), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n276), .A2(new_n281), .A3(G232), .A4(new_n283), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT69), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n276), .A2(new_n281), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G107), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n276), .A2(new_n281), .A3(G238), .A4(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n322), .A2(new_n325), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n321), .B1(new_n329), .B2(new_n289), .ZN(new_n330));
  OAI211_X1 g0130(.A(KEYINPUT71), .B(new_n320), .C1(new_n330), .C2(G169), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n320), .B1(new_n330), .B2(G169), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT71), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n320), .B1(G190), .B2(new_n330), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n272), .ZN(new_n343));
  INV_X1    g0143(.A(G169), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n343), .B1(new_n303), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G179), .B2(new_n303), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n310), .A2(new_n338), .A3(new_n342), .A4(new_n346), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT12), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n267), .B2(new_n220), .ZN(new_n350));
  INV_X1    g0150(.A(new_n270), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n348), .A2(new_n350), .B1(new_n351), .B2(new_n220), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n261), .B2(new_n226), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n354), .A2(KEYINPUT11), .A3(new_n264), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT11), .B1(new_n354), .B2(new_n264), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT13), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n221), .B1(new_n300), .B2(KEYINPUT72), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT72), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n298), .B2(new_n299), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n295), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n326), .A2(new_n365), .A3(G1698), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n276), .A2(new_n281), .A3(G232), .A4(G1698), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G97), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n289), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n360), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n299), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n288), .A2(new_n296), .A3(new_n297), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(KEYINPUT72), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(new_n363), .A3(G238), .ZN(new_n375));
  AND4_X1   g0175(.A1(new_n360), .A2(new_n370), .A3(new_n375), .A4(new_n294), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n359), .B(G169), .C1(new_n371), .C2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n370), .A2(new_n375), .A3(new_n294), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT13), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n364), .A2(new_n360), .A3(new_n370), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n359), .B1(new_n383), .B2(G169), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n358), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n379), .A2(new_n380), .A3(G190), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n371), .A2(new_n376), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n357), .B(new_n386), .C1(new_n387), .C2(new_n339), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G159), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n313), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT67), .B(G58), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n213), .B1(new_n392), .B2(new_n220), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n391), .B1(new_n393), .B2(G20), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n280), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n274), .A2(new_n275), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n398), .B2(new_n207), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n278), .A2(new_n207), .A3(new_n280), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(KEYINPUT73), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G68), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT16), .B(new_n394), .C1(new_n400), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT67), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G58), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n254), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n201), .B1(new_n408), .B2(G68), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n409), .A2(new_n207), .B1(new_n390), .B2(new_n313), .ZN(new_n410));
  AOI21_X1  g0210(.A(G20), .B1(new_n276), .B2(new_n281), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n395), .B1(new_n411), .B2(KEYINPUT7), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n410), .B1(new_n412), .B2(G68), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n264), .B(new_n405), .C1(new_n413), .C2(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n258), .A2(new_n268), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n270), .B2(new_n258), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n365), .A2(G1698), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n417), .B1(G223), .B2(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n288), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n288), .A2(G232), .A3(new_n297), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n294), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G190), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n420), .A2(new_n422), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(G200), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n414), .A2(KEYINPUT74), .A3(new_n416), .A4(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n412), .A2(G68), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT16), .B1(new_n430), .B2(new_n394), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n405), .A2(new_n264), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n416), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n420), .A2(new_n422), .A3(new_n332), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(G169), .B2(new_n425), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n427), .A2(new_n428), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n433), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n429), .A2(new_n438), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n347), .A2(new_n389), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n268), .A2(G97), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n206), .A2(G33), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n268), .A2(new_n319), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n447), .B2(G97), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n412), .A2(G107), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n252), .A2(G77), .ZN(new_n451));
  AND2_X1   g0251(.A1(G97), .A2(G107), .ZN(new_n452));
  NOR2_X1   g0252(.A1(G97), .A2(G107), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(KEYINPUT75), .B2(KEYINPUT6), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(KEYINPUT6), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(G97), .B(G107), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n451), .B1(new_n459), .B2(new_n207), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n450), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n449), .B1(new_n462), .B2(new_n264), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n206), .A2(G45), .ZN(new_n464));
  OR2_X1    g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  NAND2_X1  g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G274), .ZN(new_n468));
  AND2_X1   g0268(.A1(G1), .A2(G13), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n287), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n292), .A2(G1), .ZN(new_n472));
  INV_X1    g0272(.A(new_n466), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n288), .ZN(new_n476));
  INV_X1    g0276(.A(G257), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G250), .A2(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n283), .A2(G244), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n276), .A3(new_n281), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n398), .B2(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT76), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n288), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT76), .A4(new_n485), .ZN(new_n489));
  AOI211_X1 g0289(.A(G190), .B(new_n478), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n487), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n289), .A3(new_n489), .ZN(new_n492));
  INV_X1    g0292(.A(new_n478), .ZN(new_n493));
  AOI21_X1  g0293(.A(G200), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n463), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n460), .B1(new_n412), .B2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n448), .B1(new_n496), .B2(new_n319), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(new_n332), .A3(new_n493), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(G169), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n221), .A2(new_n283), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n227), .A2(G1698), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n502), .C1(new_n274), .C2(new_n275), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G116), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n288), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n288), .A2(G274), .A3(new_n472), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n223), .B1(new_n206), .B2(G45), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n288), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT78), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(G190), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n470), .A2(new_n472), .B1(new_n288), .B2(new_n507), .ZN(new_n513));
  INV_X1    g0313(.A(new_n504), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G238), .A2(G1698), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n227), .B2(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n278), .A2(new_n280), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n513), .B(G190), .C1(new_n518), .C2(new_n288), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT78), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n513), .B1(new_n518), .B2(new_n288), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n512), .A2(new_n520), .B1(G200), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n517), .A2(new_n207), .A3(G68), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT77), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT77), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n517), .A2(new_n525), .A3(new_n207), .A4(G68), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n260), .A2(new_n527), .A3(G97), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n453), .A2(new_n222), .B1(new_n368), .B2(new_n207), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(new_n527), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n524), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n264), .ZN(new_n532));
  INV_X1    g0332(.A(new_n317), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n267), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n447), .A2(G87), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n510), .A2(G169), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n521), .A2(G179), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n447), .A2(new_n317), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n532), .A2(new_n534), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n522), .A2(new_n536), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n495), .A2(new_n500), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G303), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n276), .B2(new_n281), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n477), .A2(new_n283), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n229), .A2(G1698), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n546), .B(new_n547), .C1(new_n274), .C2(new_n275), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n289), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n475), .A2(G270), .A3(new_n288), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n551), .A2(new_n471), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n268), .A2(G116), .A3(new_n319), .A4(new_n445), .ZN(new_n554));
  INV_X1    g0354(.A(G116), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n267), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n263), .A2(new_n216), .B1(G20), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n485), .B(new_n207), .C1(G33), .C2(new_n456), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n557), .A2(KEYINPUT20), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT20), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n554), .B(new_n556), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n553), .A2(KEYINPUT21), .A3(G169), .A4(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n561), .A2(G179), .A3(new_n550), .A4(new_n552), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n344), .B1(new_n550), .B2(new_n552), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT21), .B1(new_n565), .B2(new_n561), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n475), .A2(G264), .A3(new_n288), .ZN(new_n568));
  INV_X1    g0368(.A(G294), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n259), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G250), .A2(G1698), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n477), .B2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n570), .B1(new_n572), .B2(new_n517), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n471), .B(new_n568), .C1(new_n573), .C2(new_n288), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(G179), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n344), .B2(new_n574), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(new_n228), .A3(G20), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT79), .ZN(new_n580));
  OAI221_X1 g0380(.A(new_n578), .B1(G20), .B2(new_n504), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n207), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT22), .ZN(new_n585));
  OR3_X1    g0385(.A1(new_n222), .A2(KEYINPUT22), .A3(G20), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n326), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT24), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n583), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n319), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT25), .B1(new_n267), .B2(new_n228), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n267), .A2(KEYINPUT25), .A3(new_n228), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n447), .A2(G107), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n576), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n591), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n590), .B1(new_n583), .B2(new_n587), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n264), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n574), .A2(new_n339), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G190), .B2(new_n574), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n561), .B1(new_n553), .B2(G200), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n423), .B2(new_n553), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n567), .A2(new_n598), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n443), .A2(new_n543), .A3(new_n608), .ZN(G372));
  NAND3_X1  g0409(.A1(new_n388), .A2(new_n337), .A3(new_n334), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT83), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n385), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n611), .B1(new_n385), .B2(new_n610), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n427), .B(KEYINPUT17), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n438), .A2(KEYINPUT82), .A3(new_n441), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT82), .ZN(new_n618));
  AOI211_X1 g0418(.A(KEYINPUT18), .B(new_n435), .C1(new_n414), .C2(new_n416), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n440), .B1(new_n433), .B2(new_n436), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n310), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n495), .A2(new_n500), .A3(new_n542), .A4(new_n604), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n598), .B(KEYINPUT80), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n567), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n522), .A2(new_n536), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n539), .A2(new_n541), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n500), .ZN(new_n630));
  XNOR2_X1  g0430(.A(KEYINPUT81), .B(KEYINPUT26), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n632), .B(new_n628), .C1(new_n630), .C2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n443), .B1(new_n626), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n623), .A2(new_n346), .A3(new_n635), .ZN(G369));
  NAND3_X1  g0436(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n637), .A2(KEYINPUT84), .A3(KEYINPUT27), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT84), .B1(new_n637), .B2(KEYINPUT27), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(G213), .B1(new_n637), .B2(KEYINPUT27), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G343), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n592), .B2(new_n597), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n598), .A2(new_n645), .A3(new_n604), .ZN(new_n646));
  XOR2_X1   g0446(.A(new_n646), .B(KEYINPUT86), .Z(new_n647));
  INV_X1    g0447(.A(new_n598), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n644), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n561), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n567), .A2(new_n606), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n567), .B2(new_n650), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n567), .A2(new_n644), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n625), .B2(new_n644), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n655), .A2(new_n658), .ZN(G399));
  INV_X1    g0459(.A(new_n210), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G41), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n453), .A2(new_n222), .A3(new_n555), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n661), .A2(new_n206), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n215), .B2(new_n661), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n664), .B(KEYINPUT28), .Z(new_n665));
  INV_X1    g0465(.A(KEYINPUT31), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT87), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n505), .B2(new_n509), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n513), .B(KEYINPUT87), .C1(new_n518), .C2(new_n288), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n574), .A3(new_n669), .A4(new_n332), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n551), .A2(new_n471), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT66), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n673));
  OAI21_X1  g0473(.A(G303), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n548), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n671), .B1(new_n675), .B2(new_n289), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT30), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n492), .A2(new_n493), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n568), .B1(new_n573), .B2(new_n288), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n521), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n681), .A2(new_n676), .A3(new_n682), .A4(G179), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n550), .A2(new_n552), .A3(G179), .ZN(new_n684));
  INV_X1    g0484(.A(new_n505), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n477), .A2(G1698), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(G250), .B2(G1698), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n687), .A2(new_n398), .B1(new_n259), .B2(new_n569), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n289), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n685), .A2(new_n689), .A3(new_n513), .A4(new_n568), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT30), .B1(new_n684), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n683), .A2(new_n691), .A3(new_n499), .ZN(new_n692));
  AOI211_X1 g0492(.A(new_n666), .B(new_n643), .C1(new_n679), .C2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n495), .A2(new_n500), .A3(new_n542), .A4(new_n643), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n693), .A2(KEYINPUT88), .B1(new_n694), .B2(new_n607), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n679), .A2(new_n692), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(KEYINPUT88), .A3(KEYINPUT31), .A4(new_n644), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n643), .B1(new_n679), .B2(new_n692), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(KEYINPUT31), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(G330), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT89), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n702), .B(G330), .C1(new_n695), .C2(new_n699), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n643), .B1(new_n634), .B2(new_n626), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n630), .A2(new_n633), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n709), .B(new_n628), .C1(new_n630), .C2(new_n631), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n624), .B1(new_n598), .B2(new_n567), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT29), .B(new_n643), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n665), .B1(new_n715), .B2(G1), .ZN(G364));
  AOI21_X1  g0516(.A(new_n216), .B1(G20), .B2(new_n344), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR4_X1   g0518(.A1(new_n207), .A2(new_n332), .A3(new_n339), .A4(G190), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n282), .B1(new_n720), .B2(new_n220), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n207), .A2(new_n423), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n332), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n207), .A2(G190), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n723), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n408), .A2(new_n725), .B1(new_n728), .B2(G77), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n339), .A2(G179), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n729), .B1(new_n222), .B2(new_n731), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n207), .A2(KEYINPUT93), .A3(G190), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT93), .B1(new_n207), .B2(G190), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n730), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n721), .B(new_n732), .C1(G107), .C2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT94), .B(G159), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT95), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT32), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT32), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n207), .B1(new_n738), .B2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT96), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT96), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(G20), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT92), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n750), .A2(G97), .B1(new_n756), .B2(G50), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n737), .A2(new_n743), .A3(new_n744), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(G326), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G322), .A2(new_n725), .B1(new_n728), .B2(G311), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT33), .B(G317), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n719), .A2(new_n761), .B1(new_n746), .B2(G294), .ZN(new_n762));
  AND4_X1   g0562(.A1(new_n326), .A2(new_n759), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n731), .B(KEYINPUT97), .ZN(new_n764));
  INV_X1    g0564(.A(new_n739), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n764), .A2(G303), .B1(G329), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n763), .B(new_n766), .C1(new_n767), .C2(new_n735), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n718), .B1(new_n758), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n266), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n206), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n661), .A2(KEYINPUT90), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT90), .B1(new_n661), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n660), .A2(new_n326), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G355), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G116), .B2(new_n210), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n247), .A2(new_n292), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n660), .A2(new_n517), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n292), .B2(new_n215), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n779), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT91), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n717), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n776), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n769), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n787), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n652), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n654), .A2(new_n775), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n653), .A2(G330), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(G396));
  AND2_X1   g0596(.A1(new_n320), .A2(new_n644), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n340), .B2(new_n341), .ZN(new_n798));
  INV_X1    g0598(.A(new_n337), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n331), .A2(new_n333), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT99), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n338), .A2(new_n803), .A3(new_n798), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n337), .A2(new_n333), .A3(new_n331), .A4(new_n797), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT100), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n334), .A2(KEYINPUT100), .A3(new_n337), .A4(new_n797), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n802), .A2(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n706), .B(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n776), .B1(new_n810), .B2(new_n705), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n705), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n717), .A2(new_n785), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n775), .B1(new_n226), .B2(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n326), .B1(new_n555), .B2(new_n727), .C1(new_n720), .C2(new_n767), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n764), .A2(G107), .B1(G87), .B2(new_n736), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n739), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n815), .B(new_n818), .C1(G303), .C2(new_n756), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n749), .A2(new_n456), .B1(new_n569), .B2(new_n724), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT98), .ZN(new_n821));
  INV_X1    g0621(.A(new_n740), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G143), .A2(new_n725), .B1(new_n728), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G150), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n720), .C1(new_n755), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT34), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n735), .A2(new_n220), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n830), .B(new_n517), .C1(new_n392), .C2(new_n745), .ZN(new_n831));
  INV_X1    g0631(.A(new_n764), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n832), .A2(new_n202), .B1(new_n833), .B2(new_n739), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n831), .B(new_n834), .C1(new_n826), .C2(new_n827), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n819), .A2(new_n821), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n807), .A2(new_n808), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n803), .B1(new_n338), .B2(new_n798), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n814), .B1(new_n718), .B2(new_n836), .C1(new_n840), .C2(new_n786), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n812), .A2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(KEYINPUT35), .ZN(new_n843));
  OAI211_X1 g0643(.A(G116), .B(new_n217), .C1(new_n459), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n843), .B2(new_n459), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT36), .Z(new_n846));
  AOI211_X1 g0646(.A(new_n226), .B(new_n214), .C1(new_n408), .C2(G68), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n220), .A2(G50), .ZN(new_n848));
  OAI211_X1 g0648(.A(G1), .B(new_n266), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT101), .Z(new_n851));
  NAND2_X1  g0651(.A1(new_n433), .A2(new_n642), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n414), .A2(new_n416), .A3(new_n426), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n437), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  INV_X1    g0655(.A(new_n416), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n394), .B1(new_n400), .B2(new_n404), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT103), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT16), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(KEYINPUT103), .B(new_n394), .C1(new_n400), .C2(new_n404), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n432), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n853), .B1(new_n863), .B2(new_n435), .ZN(new_n864));
  INV_X1    g0664(.A(new_n642), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n855), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n442), .A2(new_n866), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT38), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n614), .A2(new_n617), .A3(new_n621), .ZN(new_n871));
  INV_X1    g0671(.A(new_n852), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n871), .A2(new_n872), .B1(new_n855), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n874), .B2(KEYINPUT38), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT39), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n868), .B2(new_n869), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n870), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT14), .B1(new_n387), .B2(new_n344), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n381), .A3(new_n377), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n358), .A3(new_n643), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT104), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n334), .A2(new_n337), .A3(new_n643), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n706), .B2(new_n809), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n385), .A2(KEYINPUT102), .A3(new_n388), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n357), .A2(new_n643), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT102), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n385), .A2(new_n894), .A3(new_n388), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n388), .A2(new_n891), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n883), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n879), .A2(new_n870), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n622), .A2(new_n865), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n887), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n708), .A2(new_n443), .A3(new_n712), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n623), .A2(new_n346), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n905), .B(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(G330), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT105), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n871), .A2(new_n872), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n855), .A2(new_n873), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n869), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT40), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n696), .A2(new_n644), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n666), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n698), .A2(KEYINPUT31), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n917), .B(new_n918), .C1(new_n607), .C2(new_n694), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n840), .A2(new_n893), .A3(new_n898), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n910), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  AND4_X1   g0721(.A1(new_n840), .A2(new_n893), .A3(new_n898), .A4(new_n919), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n922), .A2(KEYINPUT105), .A3(KEYINPUT40), .A4(new_n875), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n902), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n921), .A2(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n443), .A2(new_n919), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n909), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n908), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n206), .B2(new_n770), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n908), .A2(new_n929), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n851), .B1(new_n931), .B2(new_n932), .ZN(G367));
  INV_X1    g0733(.A(new_n655), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n495), .B(new_n500), .C1(new_n463), .C2(new_n643), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n500), .A2(new_n643), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n937), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n647), .A2(new_n939), .A3(new_n656), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n935), .A2(new_n598), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n644), .B1(new_n944), .B2(new_n500), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n536), .A2(new_n643), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n541), .A3(new_n539), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n629), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT106), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(KEYINPUT106), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n954), .B1(new_n947), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT108), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n938), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n938), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n661), .B(KEYINPUT41), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n658), .A2(new_n937), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT44), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n658), .A2(new_n937), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT45), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n934), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n649), .B1(new_n567), .B2(new_n644), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n657), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n654), .A2(KEYINPUT109), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n654), .A2(KEYINPUT109), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n973), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n973), .B2(new_n976), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n967), .A2(new_n934), .A3(new_n969), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n971), .A2(new_n715), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n965), .B1(new_n981), .B2(new_n715), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n963), .B(new_n964), .C1(new_n772), .C2(new_n982), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n788), .B1(new_n210), .B2(new_n533), .C1(new_n782), .C2(new_n241), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n776), .A2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G150), .A2(new_n725), .B1(new_n728), .B2(G50), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n392), .B2(new_n731), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n326), .B(new_n987), .C1(new_n719), .C2(new_n822), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n735), .A2(new_n226), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G137), .B2(new_n765), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n749), .A2(new_n220), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G143), .B2(new_n756), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n764), .A2(KEYINPUT46), .A3(G116), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT110), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n735), .A2(new_n456), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n398), .B1(new_n727), .B2(new_n767), .C1(new_n544), .C2(new_n724), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(G317), .C2(new_n765), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n731), .B2(new_n555), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n228), .B2(new_n745), .C1(new_n720), .C2(new_n569), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G311), .B2(new_n756), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n995), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT47), .Z(new_n1005));
  OAI221_X1 g0805(.A(new_n985), .B1(new_n792), .B2(new_n950), .C1(new_n1005), .C2(new_n718), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n983), .A2(new_n1006), .ZN(G387));
  AOI22_X1  g0807(.A1(G317), .A2(new_n725), .B1(new_n728), .B2(G303), .ZN(new_n1008));
  INV_X1    g0808(.A(G322), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1008), .B1(new_n817), .B2(new_n720), .C1(new_n755), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n731), .A2(new_n569), .B1(new_n745), .B2(new_n767), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n735), .A2(new_n555), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n517), .B(new_n1019), .C1(G326), .C2(new_n765), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n749), .A2(new_n533), .B1(new_n755), .B2(new_n390), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n398), .B1(new_n725), .B2(G50), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n220), .B2(new_n727), .C1(new_n226), .C2(new_n731), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n258), .A2(new_n720), .B1(new_n824), .B2(new_n739), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1022), .A2(new_n1024), .A3(new_n996), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n718), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n781), .B1(new_n238), .B2(new_n292), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n777), .A2(new_n662), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(G45), .B(new_n662), .C1(G68), .C2(G77), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n312), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT50), .B1(new_n312), .B2(G50), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1031), .A2(new_n1035), .B1(new_n228), .B2(new_n660), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n776), .B1(new_n1036), .B2(new_n789), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1028), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT111), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n649), .A2(new_n787), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT112), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1039), .A2(new_n1043), .A3(new_n1040), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n979), .A2(new_n772), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n979), .A2(new_n715), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n661), .B(KEYINPUT113), .Z(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n978), .B2(new_n714), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n1046), .B2(new_n1048), .ZN(G393));
  INV_X1    g0849(.A(new_n980), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1050), .A2(new_n970), .B1(new_n714), .B2(new_n978), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n981), .A2(new_n1051), .A3(new_n1047), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n788), .B1(new_n456), .B2(new_n210), .C1(new_n782), .C2(new_n250), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n776), .A2(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n326), .B1(new_n767), .B2(new_n731), .C1(new_n569), .C2(new_n727), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n720), .A2(new_n544), .B1(new_n745), .B2(new_n555), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n228), .B2(new_n735), .C1(new_n1009), .C2(new_n739), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n756), .A2(G317), .B1(G311), .B2(new_n725), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n750), .A2(G77), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n517), .B1(new_n727), .B2(new_n312), .C1(new_n220), .C2(new_n731), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G50), .B2(new_n719), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G87), .A2(new_n736), .B1(new_n765), .B2(G143), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n755), .A2(new_n824), .B1(new_n390), .B2(new_n724), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n1058), .A2(new_n1060), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1054), .B1(new_n1068), .B2(new_n717), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n939), .B2(new_n792), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1050), .A2(KEYINPUT114), .A3(new_n970), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT114), .B1(new_n1050), .B2(new_n970), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n772), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1052), .B(new_n1070), .C1(new_n1071), .C2(new_n1073), .ZN(G390));
  AOI21_X1  g0874(.A(new_n809), .B1(new_n701), .B2(new_n703), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n899), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n643), .B1(new_n710), .B2(new_n711), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n888), .B1(new_n1077), .B2(new_n809), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n899), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n885), .A3(new_n875), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n901), .A2(new_n886), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1076), .B(new_n1080), .C1(new_n1081), .C2(new_n881), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n920), .A2(new_n909), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1080), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n885), .A2(new_n900), .B1(new_n877), .B2(new_n880), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n919), .A2(KEYINPUT115), .A3(G330), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT115), .B1(new_n919), .B2(G330), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1088), .A2(new_n1089), .A3(new_n809), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT116), .B1(new_n1090), .B2(new_n899), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1078), .B1(new_n1075), .B2(new_n899), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT116), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n893), .A2(new_n898), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n919), .A2(G330), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n840), .B1(new_n1095), .B2(KEYINPUT115), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1093), .B(new_n1094), .C1(new_n1096), .C2(new_n1088), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1091), .A2(new_n1092), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n899), .B1(new_n704), .B2(new_n840), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n889), .B1(new_n1099), .B2(new_n1083), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n443), .A2(new_n1095), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n623), .A2(new_n906), .A3(new_n346), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT117), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1101), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1087), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1047), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1107), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1112));
  AOI211_X1 g0912(.A(KEYINPUT117), .B(new_n1103), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1087), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1082), .A2(new_n1086), .A3(new_n772), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n724), .A2(new_n833), .B1(new_n727), .B2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n326), .B(new_n1119), .C1(G137), .C2(new_n719), .ZN(new_n1120));
  INV_X1    g0920(.A(G128), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n755), .C1(new_n390), .C2(new_n749), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n731), .A2(new_n824), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1124), .B1(new_n202), .B2(new_n735), .C1(new_n1125), .C2(new_n739), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n724), .A2(new_n555), .B1(new_n727), .B2(new_n456), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n282), .B(new_n1127), .C1(G107), .C2(new_n719), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1061), .B(new_n1128), .C1(new_n767), .C2(new_n755), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n830), .B1(new_n569), .B2(new_n739), .C1(new_n832), .C2(new_n222), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1122), .A2(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n717), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n775), .B1(new_n258), .B2(new_n813), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n881), .C2(new_n786), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1117), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1116), .A2(new_n1136), .ZN(G378));
  NAND2_X1  g0937(.A1(new_n921), .A2(new_n923), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n909), .B1(new_n925), .B2(new_n924), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT119), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT119), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n310), .A2(new_n346), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n343), .A2(new_n865), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1140), .A2(new_n1141), .A3(new_n1150), .ZN(new_n1151));
  AND4_X1   g0951(.A1(KEYINPUT119), .A2(new_n1138), .A3(new_n1139), .A4(new_n1150), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n905), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n905), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1141), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1150), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT119), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1152), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1154), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1153), .A2(new_n1160), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1156), .A2(new_n786), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n813), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n776), .B1(G50), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n517), .A2(G41), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(G33), .A2(G41), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1165), .A2(G50), .A3(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1165), .B1(new_n226), .B2(new_n731), .C1(new_n228), .C2(new_n724), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1168), .B(new_n991), .C1(G97), .C2(new_n719), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n735), .A2(new_n392), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n739), .A2(new_n767), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n317), .C2(new_n728), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1169), .B(new_n1172), .C1(new_n555), .C2(new_n755), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1167), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n727), .A2(new_n825), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1121), .A2(new_n724), .B1(new_n731), .B2(new_n1118), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G132), .C2(new_n719), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n1125), .B2(new_n755), .C1(new_n824), .C2(new_n749), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1166), .B1(new_n735), .B2(new_n740), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G124), .B2(new_n765), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT118), .Z(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1175), .B1(new_n1174), .B2(new_n1173), .C1(new_n1180), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1164), .B1(new_n1186), .B2(new_n717), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1161), .A2(new_n772), .B1(new_n1162), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1103), .B(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1114), .B2(new_n1087), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1161), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT57), .B1(new_n1109), .B2(new_n1190), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n905), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1158), .A2(new_n1159), .A3(new_n1154), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1047), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1188), .B1(new_n1193), .B2(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G375));
  AOI21_X1  g1003(.A(new_n771), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n739), .A2(new_n1121), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1170), .B(new_n1205), .C1(G159), .C2(new_n764), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n755), .A2(new_n833), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n398), .B1(new_n725), .B2(G137), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n824), .B2(new_n727), .C1(new_n720), .C2(new_n1118), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1207), .B(new_n1209), .C1(G50), .C2(new_n750), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n755), .A2(new_n569), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G283), .A2(new_n725), .B1(new_n728), .B2(G107), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(new_n326), .C1(new_n555), .C2(new_n720), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(new_n317), .C2(new_n750), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n739), .A2(new_n544), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n989), .B(new_n1215), .C1(G97), .C2(new_n764), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1206), .A2(new_n1210), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n776), .B1(G68), .B2(new_n1163), .C1(new_n1217), .C2(new_n718), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1094), .B2(new_n785), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1204), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1114), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1098), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(new_n965), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1220), .B1(new_n1221), .B2(new_n1224), .ZN(G381));
  AOI21_X1  g1025(.A(new_n1135), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1226));
  OR2_X1    g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  OR3_X1    g1027(.A1(G390), .A2(G384), .A3(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1228), .A2(G387), .A3(G381), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1202), .A2(new_n1226), .A3(new_n1229), .ZN(G407));
  INV_X1    g1030(.A(G213), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(G343), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1202), .A2(new_n1226), .A3(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT122), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(G213), .A3(G407), .ZN(G409));
  OAI211_X1 g1035(.A(G378), .B(new_n1188), .C1(new_n1193), .C2(new_n1198), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1109), .A2(new_n1190), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1197), .A2(new_n1237), .A3(new_n965), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1162), .A2(new_n1187), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1197), .B2(new_n771), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1226), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1232), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1047), .B1(new_n1223), .B2(KEYINPUT60), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1106), .A2(new_n1108), .A3(new_n1222), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(KEYINPUT60), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1220), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1243), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT60), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1114), .B2(new_n1222), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G384), .B(new_n1220), .C1(new_n1250), .C2(new_n1244), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1242), .A2(KEYINPUT63), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n983), .A2(new_n1255), .A3(new_n1006), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1227), .A2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(G390), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1254), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1258), .B(G390), .Z(new_n1261));
  INV_X1    g1061(.A(new_n1256), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1255), .B1(new_n983), .B2(new_n1006), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1253), .A2(new_n1260), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1232), .ZN(new_n1266));
  INV_X1    g1066(.A(G2897), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT124), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1268), .B1(new_n1252), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1268), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(KEYINPUT124), .A3(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1270), .A2(new_n1273), .B1(new_n1269), .B2(new_n1252), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1266), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1242), .A2(new_n1252), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1278), .A2(KEYINPUT123), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT123), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1265), .B(new_n1277), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1264), .A2(KEYINPUT127), .A3(new_n1260), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT127), .B1(new_n1264), .B2(new_n1260), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1252), .A2(new_n1269), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1272), .B1(new_n1271), .B2(KEYINPUT124), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1269), .B(new_n1268), .C1(new_n1248), .C2(new_n1251), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1286), .B1(new_n1290), .B2(new_n1242), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1278), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1242), .A2(KEYINPUT62), .A3(new_n1252), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1291), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1285), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT62), .B1(new_n1242), .B2(new_n1252), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1242), .A2(KEYINPUT62), .A3(new_n1252), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1277), .B(new_n1296), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1282), .B1(new_n1297), .B2(new_n1301), .ZN(G405));
  NAND3_X1  g1102(.A1(new_n1200), .A2(new_n1226), .A3(new_n1201), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1271), .B1(new_n1303), .B2(new_n1236), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1271), .A3(new_n1236), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1285), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1303), .A2(new_n1271), .A3(new_n1236), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n1308), .A2(new_n1304), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1307), .A2(new_n1309), .ZN(G402));
endmodule


