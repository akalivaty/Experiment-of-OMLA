//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n640, new_n642, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n460), .A2(new_n462), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT65), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT66), .ZN(G160));
  NAND2_X1  g050(.A1(new_n464), .A2(G136), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n463), .A2(G112), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n469), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI221_X1 g055(.A(new_n476), .B1(new_n477), .B2(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT67), .Z(G162));
  NAND3_X1  g057(.A1(new_n469), .A2(G126), .A3(G2105), .ZN(new_n483));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n463), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n487), .A2(KEYINPUT68), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n490), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(new_n486), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(G164));
  XNOR2_X1  g071(.A(KEYINPUT69), .B(G651), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT70), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(G651), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n501), .B(KEYINPUT6), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n499), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT71), .B(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n512), .B(KEYINPUT5), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n510), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n507), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n510), .A2(new_n511), .A3(new_n516), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT73), .B1(new_n506), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT74), .B(G88), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n499), .A2(new_n505), .A3(G543), .A4(new_n500), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n497), .B1(new_n528), .B2(G50), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n523), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  AOI21_X1  g106(.A(new_n518), .B1(new_n507), .B2(new_n517), .ZN(new_n532));
  NOR3_X1   g107(.A1(new_n506), .A2(new_n520), .A3(KEYINPUT73), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n528), .A2(G51), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT76), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n535), .A2(new_n538), .A3(new_n539), .A4(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n534), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n520), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(new_n497), .B1(new_n528), .B2(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR3_X1    g127(.A1(new_n552), .A2(new_n503), .A3(new_n504), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n534), .A2(G81), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n528), .A2(G43), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n553), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n567), .B1(new_n532), .B2(new_n533), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n519), .A2(KEYINPUT78), .A3(new_n521), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(G91), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n510), .A2(new_n516), .A3(new_n572), .A4(new_n511), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(G65), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n527), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n528), .A2(new_n579), .A3(G53), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n576), .A2(G651), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n570), .A2(new_n581), .A3(KEYINPUT80), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT80), .B1(new_n570), .B2(new_n581), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G299));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n550), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n545), .A2(KEYINPUT81), .A3(new_n549), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G301));
  NAND3_X1  g164(.A1(new_n568), .A2(G87), .A3(new_n569), .ZN(new_n590));
  INV_X1    g165(.A(G74), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n502), .B1(new_n520), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n528), .B2(G49), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(G288));
  NAND3_X1  g169(.A1(new_n568), .A2(G86), .A3(new_n569), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n520), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(new_n497), .B1(new_n528), .B2(G48), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n520), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n497), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n603), .A2(KEYINPUT82), .A3(new_n497), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT84), .B(G85), .Z(new_n609));
  NAND3_X1  g184(.A1(new_n519), .A2(new_n521), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT83), .B(G47), .Z(new_n611));
  NOR2_X1   g186(.A1(new_n527), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(G290));
  INV_X1    g189(.A(G301), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n571), .A2(new_n573), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g199(.A(KEYINPUT86), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(G651), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n568), .A2(G92), .A3(new_n569), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n528), .A2(G54), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n568), .A2(new_n630), .A3(G92), .A4(new_n569), .ZN(new_n631));
  AND4_X1   g206(.A1(new_n626), .A2(new_n628), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n618), .B1(G868), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT85), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(KEYINPUT85), .B2(new_n617), .ZN(G284));
  OAI21_X1  g210(.A(new_n634), .B1(KEYINPUT85), .B2(new_n617), .ZN(G321));
  NAND2_X1  g211(.A1(G286), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n584), .B2(G868), .ZN(G297));
  OAI21_X1  g213(.A(new_n637), .B1(new_n584), .B2(G868), .ZN(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n632), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n559), .A2(new_n616), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n628), .A2(new_n626), .A3(new_n629), .A4(new_n631), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n643), .A2(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n642), .B1(new_n644), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(KEYINPUT88), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(KEYINPUT88), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n648), .B(new_n649), .C1(G111), .C2(new_n463), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n464), .A2(G135), .ZN(new_n651));
  INV_X1    g226(.A(G123), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n479), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G2096), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(KEYINPUT87), .B2(G2100), .ZN(new_n655));
  INV_X1    g230(.A(new_n467), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n469), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT12), .Z(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT13), .Z(new_n659));
  NAND2_X1  g234(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI221_X1 g236(.A(new_n661), .B1(G2096), .B2(new_n653), .C1(new_n660), .C2(new_n659), .ZN(G156));
  XOR2_X1   g237(.A(KEYINPUT15), .B(G2435), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2438), .ZN(new_n664));
  XOR2_X1   g239(.A(G2427), .B(G2430), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT89), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT14), .ZN(new_n668));
  XOR2_X1   g243(.A(G2443), .B(G2446), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1341), .B(G1348), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2451), .B(G2454), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  AND2_X1   g250(.A1(new_n675), .A2(G14), .ZN(G401));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT18), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(KEYINPUT90), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(new_n677), .ZN(new_n684));
  INV_X1    g259(.A(new_n680), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n677), .B(KEYINPUT17), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n684), .B(new_n685), .C1(new_n683), .C2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n683), .A3(new_n680), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2096), .B(G2100), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  INV_X1    g281(.A(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n705), .B(new_n708), .Z(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  INV_X1    g285(.A(G1981), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT92), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n709), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(G229));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NOR2_X1   g291(.A1(G162), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(G35), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT103), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(KEYINPUT103), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT29), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G2090), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT104), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n722), .A2(new_n723), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n716), .A2(G26), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n464), .A2(G140), .ZN(new_n728));
  OR2_X1    g303(.A1(G104), .A2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n729), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n730));
  INV_X1    g305(.A(G128), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n730), .C1(new_n731), .C2(new_n479), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n727), .B1(new_n732), .B2(G29), .ZN(new_n733));
  MUX2_X1   g308(.A(new_n727), .B(new_n733), .S(KEYINPUT28), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2067), .ZN(new_n735));
  OR2_X1    g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  NAND2_X1  g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n736), .A2(new_n716), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G160), .B2(new_n716), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G2084), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G11), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT30), .B(G28), .Z(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n735), .A2(new_n740), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n656), .A2(G103), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT99), .B(KEYINPUT25), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n464), .A2(G139), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n747), .B(new_n748), .C1(new_n463), .C2(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(G33), .B(new_n750), .S(G29), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2072), .ZN(new_n752));
  INV_X1    g327(.A(G27), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT102), .B1(new_n753), .B2(G29), .ZN(new_n754));
  OR3_X1    g329(.A1(new_n753), .A2(KEYINPUT102), .A3(G29), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n754), .B(new_n755), .C1(G164), .C2(new_n716), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2078), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n726), .A2(new_n744), .A3(new_n752), .A4(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G16), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n759), .A2(KEYINPUT23), .A3(G20), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT23), .ZN(new_n761));
  INV_X1    g336(.A(G20), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G16), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n760), .B(new_n763), .C1(new_n584), .C2(new_n759), .ZN(new_n764));
  INV_X1    g339(.A(G1956), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n759), .A2(G21), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G168), .B2(new_n759), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n725), .A2(new_n758), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(G171), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G5), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(G1961), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n739), .A2(G2084), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT101), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n716), .A2(G32), .ZN(new_n780));
  INV_X1    g355(.A(new_n479), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G129), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n656), .A2(G105), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n464), .A2(G141), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND4_X1  g361(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n780), .B1(new_n788), .B2(new_n716), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT100), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT27), .B(G1996), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  NOR4_X1   g368(.A1(new_n771), .A2(new_n775), .A3(new_n777), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G19), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n560), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT98), .B(G1341), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT36), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n590), .A2(new_n802), .A3(new_n593), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n590), .B2(new_n593), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n801), .B1(new_n805), .B2(new_n759), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G1976), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n808));
  INV_X1    g383(.A(G1976), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n809), .B(new_n801), .C1(new_n805), .C2(new_n759), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n808), .B1(new_n807), .B2(new_n810), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n759), .A2(G22), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G166), .B2(new_n759), .ZN(new_n816));
  INV_X1    g391(.A(G1971), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n759), .A2(G6), .ZN(new_n819));
  INV_X1    g394(.A(G305), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n759), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT32), .B(G1981), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n814), .A2(KEYINPUT34), .A3(new_n818), .A4(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n813), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n825), .A2(new_n818), .A3(new_n811), .A4(new_n823), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G290), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G16), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G16), .B2(G24), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(new_n707), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n716), .A2(G25), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n464), .A2(G131), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT93), .ZN(new_n836));
  OR2_X1    g411(.A1(G95), .A2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n837), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT94), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n781), .A2(G119), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n834), .B1(new_n846), .B2(new_n716), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT35), .B(G1991), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n847), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n832), .A2(new_n707), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n833), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n799), .B1(new_n829), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g429(.A(KEYINPUT36), .B(new_n852), .C1(new_n824), .C2(new_n828), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n794), .B(new_n798), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n759), .A2(G4), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n632), .B2(new_n759), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G1348), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n653), .A2(new_n716), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n856), .A2(new_n859), .A3(new_n860), .ZN(G311));
  AND4_X1   g436(.A1(new_n758), .A2(new_n725), .A3(new_n766), .A4(new_n770), .ZN(new_n862));
  INV_X1    g437(.A(new_n775), .ZN(new_n863));
  INV_X1    g438(.A(new_n793), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n776), .A4(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n854), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n829), .A2(new_n799), .A3(new_n853), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n859), .ZN(new_n869));
  INV_X1    g444(.A(new_n860), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n798), .ZN(G150));
  NAND2_X1  g446(.A1(new_n534), .A2(G93), .ZN(new_n872));
  NAND2_X1  g447(.A1(G80), .A2(G543), .ZN(new_n873));
  INV_X1    g448(.A(G67), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n520), .B2(new_n874), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n875), .A2(new_n497), .B1(new_n528), .B2(G55), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND3_X1  g454(.A1(new_n559), .A2(new_n872), .A3(new_n876), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n553), .B(new_n877), .C1(new_n557), .C2(new_n558), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n632), .A2(G559), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT38), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n883), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n879), .B1(new_n886), .B2(G860), .ZN(G145));
  XNOR2_X1  g462(.A(new_n750), .B(new_n787), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n494), .A2(new_n486), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n732), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n888), .B(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n781), .A2(G130), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n464), .A2(G142), .ZN(new_n893));
  OR2_X1    g468(.A1(G106), .A2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n894), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n843), .A2(new_n844), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n843), .B2(new_n844), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT105), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n658), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n903), .A3(new_n658), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n891), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(G160), .B(new_n653), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G162), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n891), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n906), .A2(KEYINPUT106), .A3(new_n907), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n908), .A2(new_n914), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n906), .A2(new_n907), .A3(new_n891), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n912), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g497(.A1(G290), .A2(G303), .ZN(new_n923));
  NAND4_X1  g498(.A1(G166), .A2(new_n610), .A3(new_n608), .A4(new_n613), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n923), .A2(G305), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G305), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  OAI22_X1  g501(.A1(new_n925), .A2(new_n926), .B1(new_n804), .B2(new_n803), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n924), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n820), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(G305), .A3(new_n924), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n805), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n927), .A2(new_n931), .A3(KEYINPUT109), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT109), .B1(new_n927), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT110), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n927), .A2(new_n931), .A3(new_n935), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n927), .A2(new_n931), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n927), .A2(new_n931), .A3(KEYINPUT109), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT42), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n936), .A2(new_n937), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n582), .B2(new_n583), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n570), .A2(new_n581), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT80), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n570), .A2(new_n581), .A3(KEYINPUT80), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n946), .A2(new_n952), .A3(new_n632), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n643), .B(KEYINPUT107), .C1(new_n583), .C2(new_n582), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT41), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT41), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n957), .A3(new_n954), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(KEYINPUT108), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n880), .A2(new_n644), .A3(new_n881), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n882), .B1(G559), .B2(new_n643), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n959), .A2(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n962), .A2(new_n955), .A3(new_n961), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n945), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n936), .A2(new_n937), .A3(new_n944), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n967), .A2(new_n964), .A3(new_n963), .ZN(new_n968));
  OAI21_X1  g543(.A(G868), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n877), .A2(new_n616), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(G295));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n972), .A3(new_n970), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n945), .A2(new_n965), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n967), .B1(new_n964), .B2(new_n963), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n616), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n970), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT111), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(G331));
  NOR2_X1   g554(.A1(G168), .A2(new_n550), .ZN(new_n980));
  AOI21_X1  g555(.A(G286), .B1(new_n587), .B2(new_n588), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n534), .A2(G81), .B1(new_n528), .B2(G43), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(new_n555), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n877), .B1(new_n984), .B2(new_n553), .ZN(new_n985));
  INV_X1    g560(.A(new_n881), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n880), .B(new_n881), .C1(new_n981), .C2(new_n980), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n959), .A2(new_n960), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n954), .A3(new_n953), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n992), .A3(new_n942), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n958), .B2(new_n956), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n989), .A2(new_n955), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n934), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n996), .A3(new_n917), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n990), .A2(new_n992), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n934), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(KEYINPUT43), .A3(new_n917), .A4(new_n993), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n997), .A2(new_n998), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1001), .A2(new_n917), .A3(new_n993), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n998), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1004), .B1(new_n1007), .B2(new_n1003), .ZN(G397));
  INV_X1    g583(.A(G40), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n468), .A2(new_n473), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n494), .B2(new_n486), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1011), .A2(new_n1014), .A3(KEYINPUT45), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1015), .A2(G1996), .A3(new_n787), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  INV_X1    g594(.A(G2067), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n732), .B(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(G1996), .B2(new_n787), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n1018), .B(new_n1019), .C1(new_n1015), .C2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n846), .A2(new_n849), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n845), .A2(new_n848), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1015), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(G290), .B(G1986), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1015), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT63), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n595), .A2(new_n711), .A3(new_n599), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT115), .B(G86), .Z(new_n1032));
  NAND2_X1  g607(.A1(new_n534), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1033), .A2(new_n599), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1031), .B1(new_n1034), .B2(new_n711), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1014), .A2(new_n1010), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1035), .A2(new_n1036), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n805), .B2(new_n809), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n809), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1042), .B(new_n1048), .C1(new_n805), .C2(new_n809), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n492), .A2(new_n495), .A3(new_n1012), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(KEYINPUT113), .A3(new_n1052), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1013), .A2(new_n1052), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(new_n1010), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n817), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(new_n1012), .C1(new_n494), .C2(new_n486), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1010), .A2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g638(.A(G2090), .B(new_n1063), .C1(KEYINPUT50), .C2(new_n1051), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT114), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1060), .A2(new_n1068), .A3(new_n1065), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(G8), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G303), .A2(G8), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT55), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1050), .A2(KEYINPUT119), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1072), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1068), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1077));
  AOI211_X1 g652(.A(KEYINPUT114), .B(new_n1064), .C1(new_n1059), .C2(new_n817), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1079), .B2(G8), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1030), .B1(new_n1074), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(G8), .A3(new_n1076), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1063), .B1(new_n1051), .B2(KEYINPUT50), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1087), .A2(G2084), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1011), .B1(new_n1013), .B2(new_n1052), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n769), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1041), .B(G286), .C1(new_n1088), .C2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1083), .A2(new_n1084), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1084), .B1(new_n1083), .B2(new_n1094), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1097));
  NAND2_X1  g672(.A1(new_n1050), .A2(new_n1085), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1011), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(KEYINPUT50), .B2(new_n1051), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1060), .B1(G2090), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1076), .B1(new_n1101), .B2(G8), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1103), .B2(new_n1093), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1095), .A2(new_n1096), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1106));
  XOR2_X1   g681(.A(new_n1031), .B(KEYINPUT117), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1045), .A2(new_n809), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(G288), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1106), .B1(new_n1042), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1087), .B2(new_n774), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1086), .A2(KEYINPUT124), .A3(G1961), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1059), .B2(G2078), .ZN(new_n1116));
  INV_X1    g691(.A(G2078), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1090), .A2(KEYINPUT53), .A3(new_n1117), .A4(new_n1058), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1089), .A2(new_n1090), .A3(KEYINPUT53), .A4(new_n1117), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1116), .B(new_n1120), .C1(G1961), .C2(new_n1086), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1119), .A2(new_n550), .B1(new_n1121), .B2(new_n615), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT54), .B1(new_n1119), .B2(G301), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n615), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1122), .A2(KEYINPUT54), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1039), .A2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n1127), .B(KEYINPUT121), .Z(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(G1996), .B2(new_n1059), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1129), .A2(new_n560), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1130), .A2(KEYINPUT59), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1040), .A2(new_n1020), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1132), .B(KEYINPUT60), .C1(new_n1086), .C2(G1348), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(new_n643), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1132), .B1(new_n1086), .B2(G1348), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1136), .A2(new_n1137), .B1(KEYINPUT60), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1011), .B(new_n1057), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(new_n1056), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1100), .A2(new_n765), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n947), .B(KEYINPUT57), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1146), .A2(KEYINPUT61), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1129), .A2(KEYINPUT59), .A3(new_n560), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1131), .A2(new_n1140), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1146), .A2(new_n1148), .B1(new_n643), .B2(new_n1139), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1147), .B2(new_n1145), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1125), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1158));
  OAI21_X1  g733(.A(G8), .B1(new_n1158), .B2(G286), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT51), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT51), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1158), .B2(G286), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1124), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1163), .B(new_n1165), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1157), .A2(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1103), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1110), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1029), .B1(new_n1105), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(G1996), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1015), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1172), .B(new_n1173), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n1021), .A2(new_n788), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1015), .A2(new_n1175), .B1(KEYINPUT126), .B2(KEYINPUT46), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT47), .Z(new_n1178));
  NAND3_X1  g753(.A1(new_n830), .A2(new_n707), .A3(new_n1015), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT48), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1023), .A2(new_n1026), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1025), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1023), .B1(KEYINPUT125), .B2(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1182), .A2(KEYINPUT125), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1183), .A2(new_n1184), .B1(G2067), .B2(new_n732), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1178), .B(new_n1181), .C1(new_n1185), .C2(new_n1015), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1170), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(G319), .ZN(new_n1189));
  NOR2_X1   g763(.A1(G401), .A2(new_n1189), .ZN(new_n1190));
  AND4_X1   g764(.A1(new_n691), .A2(new_n921), .A3(new_n1190), .A4(new_n714), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n999), .A2(new_n1002), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1192), .A2(KEYINPUT127), .ZN(new_n1193));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  NAND4_X1  g768(.A1(new_n999), .A2(new_n1002), .A3(new_n1191), .A4(new_n1194), .ZN(new_n1195));
  AND2_X1   g769(.A1(new_n1193), .A2(new_n1195), .ZN(G308));
  NAND2_X1  g770(.A1(new_n1193), .A2(new_n1195), .ZN(G225));
endmodule


