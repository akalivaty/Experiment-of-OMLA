//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NOR2_X1   g0012(.A1(G58), .A2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n207), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  INV_X1    g0029(.A(G238), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n209), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n212), .B(new_n219), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  INV_X1    g0044(.A(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n227), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  XNOR2_X1  g0051(.A(KEYINPUT79), .B(KEYINPUT21), .ZN(new_n252));
  AND2_X1   g0052(.A1(G264), .A2(G1698), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT77), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n254), .A2(new_n255), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G303), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  OAI211_X1 g0061(.A(G257), .B(new_n261), .C1(new_n254), .C2(new_n255), .ZN(new_n262));
  OAI211_X1 g0062(.A(KEYINPUT77), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n258), .A2(new_n260), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n206), .A2(G45), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  AND2_X1   g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n273), .ZN(new_n277));
  INV_X1    g0077(.A(new_n275), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n206), .B(G45), .C1(new_n267), .C2(KEYINPUT5), .ZN(new_n279));
  OAI211_X1 g0079(.A(G270), .B(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n266), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G283), .ZN(new_n285));
  INV_X1    g0085(.A(G97), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n207), .C1(G33), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n217), .ZN(new_n289));
  INV_X1    g0089(.A(G116), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n287), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n287), .A2(KEYINPUT20), .A3(new_n289), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G116), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n206), .A2(G33), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n297), .A2(new_n299), .A3(new_n217), .A4(new_n288), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n298), .B1(new_n301), .B2(G116), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n284), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n283), .A2(new_n303), .A3(KEYINPUT78), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT78), .B1(new_n283), .B2(new_n303), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n252), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n281), .B1(new_n264), .B2(new_n265), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n296), .A2(new_n302), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G179), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n283), .A2(new_n303), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT21), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n283), .B2(G200), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n283), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n307), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n297), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n289), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n206), .A2(G20), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(G50), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G50), .B2(new_n297), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT8), .B(G58), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n207), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(G20), .A2(G33), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n327), .B1(G150), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n202), .A2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n324), .B1(new_n331), .B2(new_n289), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT9), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n332), .B(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT3), .A2(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n261), .A2(G222), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G223), .A2(G1698), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n340), .B(new_n265), .C1(G77), .C2(new_n337), .ZN(new_n341));
  INV_X1    g0141(.A(G45), .ZN(new_n342));
  AOI21_X1  g0142(.A(G1), .B1(new_n267), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n277), .A2(G274), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G226), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n277), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n341), .B(new_n344), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n316), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(G200), .B2(new_n348), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n334), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT10), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n348), .A2(G179), .ZN(new_n353));
  AOI211_X1 g0153(.A(new_n332), .B(new_n353), .C1(new_n284), .C2(new_n348), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(G232), .A2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n254), .B2(new_n255), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT69), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  OAI211_X1 g0160(.A(G226), .B(new_n261), .C1(new_n254), .C2(new_n255), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT69), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n357), .C1(new_n254), .C2(new_n255), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n265), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n344), .A2(KEYINPUT70), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT70), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n274), .A2(new_n367), .A3(new_n343), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n265), .A2(new_n343), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n366), .A2(new_n368), .B1(G238), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n365), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n365), .B2(new_n370), .ZN(new_n374));
  OAI21_X1  g0174(.A(G200), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n328), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n376), .A2(new_n245), .B1(new_n207), .B2(G68), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n326), .A2(new_n221), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n289), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT11), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n320), .A2(new_n229), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT12), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT71), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n384), .A3(KEYINPUT12), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n383), .B(new_n385), .C1(KEYINPUT12), .C2(new_n381), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n321), .A2(G68), .A3(new_n322), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n365), .A2(new_n370), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(G190), .A3(new_n372), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n375), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n373), .A2(new_n374), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT14), .B1(new_n395), .B2(new_n284), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n391), .A2(G179), .A3(new_n372), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT14), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(G169), .C1(new_n373), .C2(new_n374), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n394), .B1(new_n400), .B2(new_n388), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n335), .A2(new_n207), .A3(new_n336), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n336), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n229), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n227), .A2(new_n229), .ZN(new_n409));
  OAI21_X1  g0209(.A(G20), .B1(new_n409), .B2(new_n213), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n328), .A2(G159), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n403), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT7), .B1(new_n259), .B2(new_n207), .ZN(new_n414));
  NOR4_X1   g0214(.A1(new_n254), .A2(new_n255), .A3(new_n405), .A4(G20), .ZN(new_n415));
  OAI21_X1  g0215(.A(G68), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n412), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(KEYINPUT16), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n413), .A2(new_n418), .A3(new_n289), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n325), .B1(new_n206), .B2(G20), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n321), .B1(new_n320), .B2(new_n325), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n345), .A2(G1698), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n422), .B1(G223), .B2(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n265), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n369), .A2(G232), .B1(new_n274), .B2(new_n343), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n316), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n277), .B1(new_n423), .B2(new_n424), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n344), .B1(new_n347), .B2(new_n228), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n419), .A2(new_n421), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT72), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT72), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n419), .A2(new_n433), .A3(new_n436), .A4(new_n421), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(KEYINPUT17), .A3(new_n437), .ZN(new_n438));
  XOR2_X1   g0238(.A(KEYINPUT73), .B(KEYINPUT17), .Z(new_n439));
  NAND4_X1  g0239(.A1(new_n419), .A2(new_n433), .A3(new_n421), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G179), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n426), .A2(new_n442), .A3(new_n427), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n284), .B1(new_n430), .B2(new_n431), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n419), .B2(new_n421), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT18), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n369), .A2(G244), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n344), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT67), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT67), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n452), .A3(new_n344), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G238), .A2(G1698), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n337), .B(new_n454), .C1(new_n228), .C2(G1698), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n265), .C1(G107), .C2(new_n337), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT68), .ZN(new_n458));
  OR3_X1    g0258(.A1(new_n457), .A2(new_n458), .A3(new_n316), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n457), .B2(new_n316), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT15), .B(G87), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n461), .A2(new_n326), .B1(new_n207), .B2(new_n221), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n325), .A2(new_n376), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n289), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n321), .A2(G77), .A3(new_n322), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(G77), .C2(new_n297), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n457), .B2(G200), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n460), .A3(new_n467), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n457), .A2(G179), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n457), .A2(new_n284), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n466), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR4_X1   g0272(.A1(new_n356), .A2(new_n402), .A3(new_n448), .A4(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(G257), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n474));
  OAI211_X1 g0274(.A(G250), .B(new_n261), .C1(new_n254), .C2(new_n255), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G294), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n265), .B1(new_n270), .B2(new_n275), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n265), .A2(new_n477), .B1(new_n478), .B2(G264), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n276), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n429), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n477), .A2(new_n265), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(G264), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n482), .A2(new_n483), .A3(new_n276), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n316), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n320), .A2(KEYINPUT25), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT25), .B1(new_n320), .B2(new_n487), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n489), .A2(new_n490), .B1(new_n487), .B2(new_n300), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n207), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT22), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n337), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n497));
  OAI211_X1 g0297(.A(KEYINPUT80), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT23), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(new_n487), .A3(G20), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n496), .A2(new_n497), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT24), .ZN(new_n507));
  AND4_X1   g0307(.A1(new_n505), .A2(new_n498), .A3(new_n499), .A4(new_n501), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n497), .A4(new_n496), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n493), .B1(new_n511), .B2(new_n289), .ZN(new_n512));
  INV_X1    g0312(.A(new_n289), .ZN(new_n513));
  AOI211_X1 g0313(.A(KEYINPUT81), .B(new_n513), .C1(new_n507), .C2(new_n510), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n486), .B(new_n492), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n320), .A2(new_n286), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n300), .B2(new_n286), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n286), .A2(new_n487), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n487), .A2(KEYINPUT6), .A3(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(G20), .B1(G77), .B2(new_n328), .ZN(new_n524));
  OAI21_X1  g0324(.A(G107), .B1(new_n414), .B2(new_n415), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n517), .B1(new_n526), .B2(new_n289), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(G257), .B(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n276), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n224), .B1(new_n335), .B2(new_n336), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT74), .ZN(new_n533));
  OAI211_X1 g0333(.A(G244), .B(new_n261), .C1(new_n254), .C2(new_n255), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(G1698), .B1(new_n335), .B2(new_n336), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n537), .A2(KEYINPUT74), .A3(KEYINPUT4), .A4(G244), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n532), .A2(new_n536), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n530), .B1(new_n540), .B2(new_n265), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n442), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n528), .B(new_n542), .C1(G169), .C2(new_n541), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(G190), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(new_n527), .C1(new_n429), .C2(new_n541), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n515), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n207), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT75), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n551), .A3(new_n207), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n223), .A2(new_n286), .A3(new_n487), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT76), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n326), .C2(new_n286), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n337), .A2(new_n207), .A3(G68), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n326), .B2(new_n286), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n554), .A2(new_n557), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n289), .ZN(new_n562));
  INV_X1    g0362(.A(new_n461), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n301), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n461), .A2(new_n320), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n206), .A2(new_n271), .A3(G45), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n224), .B1(new_n342), .B2(G1), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n277), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n230), .A2(new_n261), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n222), .A2(G1698), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n571), .C1(new_n254), .C2(new_n255), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G179), .B(new_n569), .C1(new_n574), .C2(new_n277), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n277), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  INV_X1    g0376(.A(new_n569), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n575), .B1(new_n284), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n566), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n301), .A2(G87), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n562), .A2(new_n565), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(G190), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n429), .B2(new_n578), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n492), .B1(new_n512), .B2(new_n514), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT82), .B1(new_n480), .B2(new_n442), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT82), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n484), .A2(new_n588), .A3(G179), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n587), .B(new_n589), .C1(new_n284), .C2(new_n484), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n585), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n319), .A2(new_n473), .A3(new_n547), .A4(new_n591), .ZN(G372));
  NAND2_X1  g0392(.A1(new_n579), .A2(KEYINPUT83), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT83), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n575), .B(new_n594), .C1(new_n578), .C2(new_n284), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n566), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n582), .A2(KEYINPUT84), .ZN(new_n598));
  INV_X1    g0398(.A(new_n584), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT84), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n562), .A2(new_n600), .A3(new_n565), .A4(new_n581), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n515), .A2(new_n543), .A3(new_n545), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n252), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT78), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n309), .A2(G169), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(new_n308), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n607), .B2(new_n304), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n313), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n586), .A2(new_n590), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n597), .B1(new_n603), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n540), .A2(new_n265), .ZN(new_n613));
  INV_X1    g0413(.A(new_n530), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n527), .B1(new_n284), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n602), .A2(new_n616), .A3(new_n596), .A4(new_n542), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n543), .A2(new_n585), .ZN(new_n618));
  MUX2_X1   g0418(.A(new_n617), .B(new_n618), .S(KEYINPUT26), .Z(new_n619));
  NAND2_X1  g0419(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n473), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n399), .A2(new_n397), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n391), .A2(new_n372), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n398), .B1(new_n623), .B2(G169), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n388), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n471), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n393), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n441), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n447), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n354), .B1(new_n630), .B2(new_n352), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n621), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g0432(.A(new_n632), .B(KEYINPUT85), .Z(G369));
  INV_X1    g0433(.A(new_n309), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n609), .A2(new_n317), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n608), .B2(new_n313), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT86), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n586), .A2(new_n640), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n515), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n610), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT87), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n586), .A2(new_n590), .A3(new_n641), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n648), .A2(new_n515), .B1(new_n586), .B2(new_n590), .ZN(new_n654));
  INV_X1    g0454(.A(new_n652), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT87), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n647), .A2(new_n657), .A3(G330), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n609), .A2(new_n640), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n653), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n652), .A3(new_n660), .ZN(G399));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  INV_X1    g0462(.A(new_n210), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(G41), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n210), .A2(KEYINPUT88), .A3(new_n267), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n553), .A2(G116), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n215), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n640), .B1(new_n612), .B2(new_n619), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT29), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n603), .A2(new_n611), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n543), .B2(new_n585), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n617), .B2(new_n674), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n596), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(KEYINPUT29), .A3(new_n641), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G330), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n576), .A2(new_n577), .A3(new_n442), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n479), .A2(new_n681), .A3(new_n266), .A4(new_n282), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT30), .B1(new_n615), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n479), .A2(new_n681), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n541), .A3(new_n685), .A4(new_n308), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n442), .B1(new_n576), .B2(new_n577), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n484), .A2(new_n308), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n615), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n641), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n690), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n641), .A2(new_n693), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n547), .A2(new_n319), .A3(new_n591), .A4(new_n641), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n680), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n679), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n670), .B1(new_n701), .B2(G1), .ZN(G364));
  INV_X1    g0502(.A(new_n666), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n207), .A2(G13), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n206), .B1(new_n704), .B2(G45), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n647), .B2(G330), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(G330), .B2(new_n647), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n210), .A2(new_n337), .ZN(new_n710));
  INV_X1    g0510(.A(G355), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n710), .A2(new_n711), .B1(G116), .B2(new_n210), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n210), .A2(new_n259), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT89), .Z(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n342), .B2(new_n216), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n247), .A2(G45), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n272), .B1(new_n207), .B2(G169), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n207), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT90), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT92), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n707), .B1(new_n718), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n442), .A2(new_n429), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n207), .B1(new_n732), .B2(G190), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n207), .A2(G190), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n442), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n734), .A2(G294), .B1(G311), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G326), .ZN(new_n740));
  NAND3_X1  g0540(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n316), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT95), .Z(new_n743));
  OAI21_X1  g0543(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT96), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n741), .A2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(KEYINPUT33), .A2(G317), .ZN(new_n748));
  NAND2_X1  g0548(.A1(KEYINPUT33), .A2(G317), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n207), .A2(new_n316), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n736), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n337), .B1(new_n753), .B2(G322), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n429), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n735), .ZN(new_n757));
  INV_X1    g0557(.A(G303), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n751), .A2(new_n756), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n754), .B1(new_n755), .B2(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n732), .A2(new_n735), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n750), .B(new_n760), .C1(G329), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n745), .A2(new_n763), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n337), .B1(new_n752), .B2(new_n227), .C1(new_n229), .C2(new_n747), .ZN(new_n765));
  INV_X1    g0565(.A(new_n757), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G77), .A2(new_n738), .B1(new_n766), .B2(G107), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(new_n223), .B2(new_n759), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n765), .B(new_n768), .C1(G50), .C2(new_n742), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n761), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n769), .B(new_n773), .C1(new_n286), .C2(new_n733), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n764), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n729), .B1(new_n775), .B2(new_n722), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n647), .B2(new_n726), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n709), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n466), .A2(new_n640), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n468), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n471), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n627), .A2(new_n641), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n671), .B(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n707), .B1(new_n785), .B2(new_n699), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n699), .B2(new_n785), .ZN(new_n787));
  INV_X1    g0587(.A(new_n707), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n722), .A2(new_n724), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(new_n221), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n337), .B1(new_n738), .B2(G116), .ZN(new_n791));
  INV_X1    g0591(.A(new_n742), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n791), .B1(new_n792), .B2(new_n758), .C1(new_n755), .C2(new_n747), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n753), .A2(G294), .ZN(new_n794));
  INV_X1    g0594(.A(new_n759), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G107), .A2(new_n795), .B1(new_n766), .B2(G87), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n794), .B(new_n796), .C1(new_n761), .C2(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n793), .B(new_n798), .C1(G97), .C2(new_n734), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n259), .B1(new_n766), .B2(G68), .ZN(new_n800));
  INV_X1    g0600(.A(G132), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n800), .B1(new_n245), .B2(new_n759), .C1(new_n761), .C2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT97), .B(G143), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n753), .A2(new_n804), .B1(new_n738), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  INV_X1    g0606(.A(G150), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n792), .B2(new_n806), .C1(new_n807), .C2(new_n747), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT34), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n802), .B(new_n810), .C1(G58), .C2(new_n734), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n799), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n724), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n790), .B1(new_n723), .B2(new_n813), .C1(new_n784), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n787), .A2(new_n815), .ZN(G384));
  OR2_X1    g0616(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n817), .A2(G116), .A3(new_n218), .A4(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT36), .Z(new_n820));
  OR3_X1    g0620(.A1(new_n215), .A2(new_n221), .A3(new_n409), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n245), .A2(G68), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n206), .B(G13), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT103), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n694), .A2(new_n825), .A3(new_n695), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n683), .A2(new_n686), .B1(new_n615), .B2(new_n689), .ZN(new_n827));
  INV_X1    g0627(.A(new_n695), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT103), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT102), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n691), .B2(KEYINPUT31), .ZN(new_n832));
  OAI211_X1 g0632(.A(KEYINPUT102), .B(new_n693), .C1(new_n827), .C2(new_n641), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n585), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n610), .A2(new_n835), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n836), .A2(new_n546), .A3(new_n318), .A4(new_n640), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n784), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT98), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n388), .A2(new_n640), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n401), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n625), .A2(new_n393), .A3(new_n840), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT98), .ZN(new_n843));
  INV_X1    g0643(.A(new_n840), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n841), .A2(new_n843), .B1(new_n400), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n413), .A2(new_n418), .A3(new_n289), .ZN(new_n847));
  INV_X1    g0647(.A(new_n421), .ZN(new_n848));
  AOI21_X1  g0648(.A(G169), .B1(new_n426), .B2(new_n427), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n430), .A2(new_n431), .A3(G179), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n638), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n847), .A2(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n435), .A2(new_n853), .A3(new_n854), .A4(new_n437), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT99), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n419), .A2(new_n421), .B1(new_n445), .B2(new_n638), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n859), .A2(KEYINPUT99), .A3(new_n435), .A4(new_n437), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n435), .A2(new_n853), .A3(new_n437), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n857), .A2(new_n860), .B1(KEYINPUT37), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n419), .A2(new_n421), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n852), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n441), .B2(new_n447), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n857), .A2(new_n860), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n854), .B1(new_n853), .B2(new_n434), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT100), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n869), .B1(new_n857), .B2(new_n860), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n865), .B1(new_n874), .B2(KEYINPUT100), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n846), .B(KEYINPUT40), .C1(new_n867), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n400), .A2(new_n844), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n839), .B1(new_n401), .B2(new_n840), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n842), .A2(KEYINPUT98), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n697), .A2(new_n832), .A3(new_n830), .A4(new_n833), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n784), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n868), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n864), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n448), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(new_n867), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n878), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n877), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT104), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n473), .A2(new_n883), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n896), .A2(new_n897), .A3(new_n680), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n671), .A2(new_n784), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n783), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n882), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n901), .A2(new_n890), .B1(new_n447), .B2(new_n852), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT101), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n876), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n866), .B1(new_n862), .B2(new_n865), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n905), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n903), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT39), .B1(new_n889), .B2(new_n867), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(KEYINPUT101), .C1(new_n876), .C2(new_n906), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n626), .A2(new_n641), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n902), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n672), .A2(new_n473), .A3(new_n678), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n631), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n898), .A2(new_n919), .B1(new_n206), .B2(new_n704), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n898), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n824), .B1(new_n920), .B2(new_n921), .ZN(G367));
  NOR2_X1   g0722(.A1(new_n238), .A2(new_n715), .ZN(new_n923));
  INV_X1    g0723(.A(new_n728), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n210), .B2(new_n461), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n707), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT107), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n641), .B1(new_n598), .B2(new_n601), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n597), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n602), .A2(new_n596), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n928), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n337), .B1(new_n752), .B2(new_n807), .C1(new_n770), .C2(new_n747), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n766), .A2(G77), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n227), .B2(new_n759), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n932), .B(new_n934), .C1(G50), .C2(new_n738), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n734), .A2(G68), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n762), .A2(G137), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n743), .A2(new_n803), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n766), .A2(G97), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n758), .B2(new_n752), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n746), .A2(G294), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n259), .B1(new_n737), .B2(new_n755), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT46), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n759), .A2(new_n944), .A3(new_n290), .ZN(new_n945));
  NOR4_X1   g0745(.A1(new_n941), .A2(new_n942), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n487), .B2(new_n733), .C1(new_n797), .C2(new_n743), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n944), .B1(new_n759), .B2(new_n290), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n762), .A2(G317), .B1(KEYINPUT108), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(KEYINPUT108), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n939), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT47), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n722), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n927), .B1(new_n726), .B2(new_n931), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT109), .Z(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n660), .A2(new_n652), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n543), .B(new_n545), .C1(new_n527), .C2(new_n641), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n616), .A2(new_n542), .A3(new_n640), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n958), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n660), .A2(KEYINPUT45), .A3(new_n652), .A4(new_n962), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n962), .B1(new_n660), .B2(new_n652), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n966), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n658), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n653), .A2(new_n656), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT86), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n646), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n974), .B1(new_n976), .B2(new_n680), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n977), .A2(new_n658), .A3(new_n659), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n659), .B1(new_n977), .B2(new_n658), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n978), .A2(new_n700), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n967), .B(KEYINPUT44), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n658), .A3(new_n966), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n973), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n701), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n666), .B(KEYINPUT41), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n706), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT42), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n653), .A2(new_n656), .A3(new_n659), .A4(new_n962), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n992), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(KEYINPUT42), .A3(new_n990), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n543), .B1(new_n960), .B2(new_n610), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n641), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT105), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n931), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n996), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n996), .B2(new_n998), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1004), .A2(new_n1007), .B1(new_n658), .B2(new_n963), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n658), .A2(new_n963), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n996), .A2(new_n998), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1003), .C1(new_n1010), .C2(new_n1006), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n957), .B1(new_n987), .B2(new_n1012), .ZN(G387));
  NOR2_X1   g0813(.A1(new_n980), .A2(new_n666), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n978), .A2(new_n979), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n701), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n325), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n245), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n667), .B(new_n342), .C1(new_n229), .C2(new_n221), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n714), .B1(new_n1019), .B2(new_n1020), .C1(new_n242), .C2(new_n342), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(G107), .B2(new_n210), .C1(new_n667), .C2(new_n710), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n788), .B1(new_n1022), .B2(new_n924), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n734), .A2(new_n563), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n245), .B2(new_n752), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT110), .Z(new_n1026));
  AOI22_X1  g0826(.A1(new_n738), .A2(G68), .B1(new_n1017), .B2(new_n746), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT111), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n795), .A2(G77), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1029), .A2(new_n940), .A3(new_n337), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n807), .B2(new_n761), .C1(new_n770), .C2(new_n792), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1026), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n761), .A2(new_n740), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n259), .B1(new_n757), .B2(new_n290), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G317), .A2(new_n753), .B1(new_n738), .B2(G303), .ZN(new_n1035));
  XOR2_X1   g0835(.A(KEYINPUT112), .B(G322), .Z(new_n1036));
  OAI221_X1 g0836(.A(new_n1035), .B1(new_n797), .B2(new_n747), .C1(new_n743), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT48), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n734), .A2(G283), .B1(G294), .B2(new_n795), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1033), .B(new_n1034), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1032), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1023), .B1(new_n1047), .B2(new_n723), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n726), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1048), .B1(new_n974), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1015), .B2(new_n706), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1016), .A2(new_n1051), .ZN(G393));
  INV_X1    g0852(.A(new_n982), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n658), .B1(new_n981), .B2(new_n966), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n963), .A2(new_n1049), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n924), .B1(new_n286), .B2(new_n210), .C1(new_n250), .C2(new_n715), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT114), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n788), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n742), .A2(G317), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n797), .B2(new_n752), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT52), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n734), .A2(G116), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n759), .A2(new_n755), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n259), .B1(new_n757), .B2(new_n487), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(G294), .C2(new_n738), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n758), .B2(new_n747), .C1(new_n761), .C2(new_n1036), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n734), .A2(G77), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n337), .B1(new_n757), .B2(new_n223), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n759), .A2(new_n229), .B1(new_n737), .B2(new_n325), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G50), .C2(new_n746), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1070), .B(new_n1073), .C1(new_n761), .C2(new_n803), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n753), .A2(G159), .B1(G150), .B2(new_n742), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT51), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1065), .A2(new_n1069), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT115), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n723), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1060), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1055), .A2(new_n706), .B1(new_n1056), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n980), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1084), .A2(new_n703), .A3(new_n983), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1082), .A2(new_n1085), .ZN(G390));
  NAND2_X1  g0886(.A1(new_n901), .A2(new_n914), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n910), .A2(new_n912), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n882), .A2(new_n698), .A3(new_n784), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n677), .A2(new_n641), .A3(new_n782), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1090), .A2(new_n783), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n914), .B1(new_n876), .B2(new_n867), .C1(new_n1091), .C2(new_n845), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n883), .A2(G330), .A3(new_n784), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n845), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n917), .B(new_n631), .C1(new_n680), .C2(new_n894), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1090), .A2(new_n783), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n698), .A2(new_n784), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n882), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1094), .A2(new_n845), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(KEYINPUT116), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n1091), .A3(new_n1089), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1101), .A2(new_n882), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n900), .B1(new_n1109), .B2(new_n1095), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1099), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n666), .B1(new_n1098), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1095), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1088), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT116), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1117));
  AND4_X1   g0917(.A1(KEYINPUT116), .A2(new_n1103), .A3(new_n1091), .A4(new_n1089), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1099), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT117), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(KEYINPUT117), .B(new_n1121), .C1(new_n1093), .C2(new_n1097), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1112), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n913), .A2(new_n814), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n259), .B1(new_n759), .B2(new_n223), .C1(new_n755), .C2(new_n792), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G107), .B2(new_n746), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n762), .A2(G294), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n752), .A2(new_n290), .B1(new_n757), .B2(new_n229), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G97), .B2(new_n738), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1070), .A2(new_n1128), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT53), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n759), .B2(new_n807), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n795), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n762), .A2(G125), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1137), .A2(new_n737), .B1(new_n757), .B2(new_n245), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n259), .B(new_n1138), .C1(G132), .C2(new_n753), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G128), .A2(new_n742), .B1(new_n746), .B2(G137), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n733), .A2(new_n770), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1132), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n722), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n789), .A2(new_n325), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n707), .A3(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1116), .A2(new_n705), .B1(new_n1126), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1125), .A2(new_n1148), .ZN(G378));
  NAND3_X1  g0949(.A1(new_n1114), .A2(new_n1115), .A3(new_n1111), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1120), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n332), .A2(new_n638), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n356), .B(new_n1154), .Z(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n356), .B(new_n1154), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1156), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1161), .A2(new_n877), .A3(G330), .A4(new_n891), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n877), .A2(G330), .A3(new_n891), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n916), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1162), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n912), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n868), .A2(KEYINPUT100), .A3(new_n870), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n888), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n874), .A2(KEYINPUT100), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n866), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT101), .B1(new_n1174), .B2(new_n911), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n915), .B1(new_n1168), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n902), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1167), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1152), .B1(new_n1166), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1151), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n703), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(KEYINPUT119), .A3(new_n1162), .A4(new_n1165), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n914), .B1(new_n910), .B2(new_n912), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT119), .B1(new_n1184), .B2(new_n902), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1167), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1151), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1183), .A2(new_n1186), .A3(new_n706), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1164), .A2(new_n724), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G50), .B1(new_n336), .B2(new_n267), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n757), .A2(new_n227), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n752), .A2(new_n487), .B1(new_n737), .B2(new_n461), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n762), .C2(G283), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n742), .A2(G116), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1029), .A2(new_n267), .A3(new_n259), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G97), .B2(new_n746), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n936), .A3(new_n1195), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT58), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1191), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(G128), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1201), .A2(new_n752), .B1(new_n759), .B2(new_n1137), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G137), .B2(new_n738), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G125), .A2(new_n742), .B1(new_n746), .B2(G132), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n733), .C2(new_n807), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n762), .A2(G124), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n766), .C2(G159), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1200), .B1(new_n1199), .B2(new_n1198), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n722), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n789), .A2(new_n245), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1190), .A2(new_n707), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1189), .A2(KEYINPUT120), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT120), .B1(new_n1189), .B2(new_n1214), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1182), .A2(new_n1188), .B1(new_n1215), .B2(new_n1216), .ZN(G375));
  OAI211_X1 g1017(.A(new_n1099), .B(new_n1110), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1121), .A2(new_n986), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n845), .A2(new_n724), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT121), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n337), .B1(new_n757), .B2(new_n227), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n762), .A2(G128), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n752), .A2(new_n806), .B1(new_n737), .B2(new_n807), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G159), .B2(new_n795), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1137), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1227), .A2(new_n746), .B1(G132), .B2(new_n742), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(new_n733), .C2(new_n245), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1224), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n742), .A2(G294), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n933), .A2(new_n259), .A3(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G97), .A2(new_n795), .B1(new_n753), .B2(G283), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n487), .B2(new_n737), .C1(new_n761), .C2(new_n758), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(G116), .C2(new_n746), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1230), .B1(new_n1235), .B2(new_n1024), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(new_n723), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n788), .B(new_n1237), .C1(new_n229), .C2(new_n789), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1119), .A2(new_n706), .B1(new_n1220), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1219), .A2(new_n1239), .ZN(G381));
  NAND3_X1  g1040(.A1(new_n1016), .A2(new_n778), .A3(new_n1051), .ZN(new_n1241));
  OR4_X1    g1041(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1241), .ZN(new_n1242));
  OR4_X1    g1042(.A1(G387), .A2(new_n1242), .A3(G375), .A4(G378), .ZN(G407));
  AND2_X1   g1043(.A1(new_n1125), .A2(new_n1148), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n639), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G375), .C2(new_n1247), .ZN(G409));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT124), .B1(G387), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1241), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n985), .B1(new_n983), .B2(new_n701), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1008), .B(new_n1011), .C1(new_n1253), .C2(new_n706), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n957), .A3(G390), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G390), .B1(new_n1254), .B2(new_n957), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1250), .A2(new_n1252), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1257), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1252), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1259), .A2(KEYINPUT124), .A3(new_n1260), .A4(new_n1255), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1258), .A2(new_n1261), .A3(KEYINPUT125), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1099), .B1(new_n1098), .B2(new_n1111), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1267), .A2(new_n985), .A3(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1166), .A2(new_n1179), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1214), .B1(new_n1270), .B2(new_n705), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1125), .B(new_n1148), .C1(new_n1269), .C2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(G375), .B2(new_n1244), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT122), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1218), .A2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n1110), .A4(new_n1099), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(new_n1121), .A3(new_n703), .A4(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1278), .A2(G384), .A3(new_n1239), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1278), .B2(new_n1239), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1239), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1278), .A2(G384), .A3(new_n1239), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(KEYINPUT122), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1281), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1273), .A2(new_n1245), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1216), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1189), .A2(KEYINPUT120), .A3(new_n1214), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1152), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n666), .B1(new_n1151), .B2(new_n1180), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(G378), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1246), .B1(new_n1297), .B2(new_n1272), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1288), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1290), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1246), .A2(G2897), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1281), .A2(new_n1286), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT123), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT123), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1281), .A2(new_n1286), .A3(new_n1306), .A4(new_n1303), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(G2897), .A3(new_n1246), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1305), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1302), .B1(new_n1310), .B2(new_n1298), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1266), .B1(new_n1301), .B2(new_n1311), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1313), .B(new_n1302), .C1(new_n1310), .C2(new_n1298), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1289), .A2(KEYINPUT63), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1298), .A2(new_n1317), .A3(new_n1288), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1315), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1312), .A2(new_n1320), .ZN(G405));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1265), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT125), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1264), .A2(KEYINPUT127), .A3(new_n1265), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G375), .A2(new_n1244), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(new_n1297), .A3(new_n1308), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1287), .B1(new_n1327), .B2(new_n1297), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1328), .B1(new_n1329), .B2(KEYINPUT126), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(KEYINPUT126), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1325), .B(new_n1326), .C1(new_n1330), .C2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(G375), .A2(new_n1244), .ZN(new_n1334));
  AOI21_X1  g1134(.A(G378), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1288), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1338));
  AOI22_X1  g1138(.A1(new_n1336), .A2(new_n1337), .B1(new_n1338), .B2(new_n1308), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(KEYINPUT127), .A4(new_n1331), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1333), .A2(new_n1341), .ZN(G402));
endmodule


