

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G651), .A2(n600), .ZN(n816) );
  NOR2_X2 U555 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XOR2_X1 U556 ( .A(G651), .B(KEYINPUT68), .Z(n522) );
  NOR2_X1 U557 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U558 ( .A1(n682), .A2(n796), .ZN(n684) );
  XNOR2_X1 U559 ( .A(n681), .B(KEYINPUT76), .ZN(n796) );
  INV_X1 U560 ( .A(n665), .ZN(n723) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n651) );
  BUF_X1 U562 ( .A(n685), .Z(n548) );
  AND2_X1 U563 ( .A1(n665), .A2(G1996), .ZN(n667) );
  AND2_X1 U564 ( .A1(n755), .A2(n743), .ZN(n744) );
  NAND2_X1 U565 ( .A1(G160), .A2(G40), .ZN(n653) );
  XNOR2_X1 U566 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n526) );
  XNOR2_X1 U567 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n523) );
  AND2_X1 U568 ( .A1(n690), .A2(n689), .ZN(n524) );
  INV_X1 U569 ( .A(KEYINPUT26), .ZN(n666) );
  INV_X1 U570 ( .A(KEYINPUT97), .ZN(n701) );
  AND2_X1 U571 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U572 ( .A(n523), .B(KEYINPUT32), .ZN(n731) );
  XNOR2_X1 U573 ( .A(n732), .B(n731), .ZN(n757) );
  INV_X1 U574 ( .A(KEYINPUT103), .ZN(n765) );
  XNOR2_X1 U575 ( .A(n688), .B(KEYINPUT77), .ZN(n691) );
  AND2_X1 U576 ( .A1(n691), .A2(n524), .ZN(n692) );
  XNOR2_X1 U577 ( .A(n527), .B(n526), .ZN(n530) );
  XNOR2_X1 U578 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n773) );
  BUF_X1 U579 ( .A(n796), .Z(n984) );
  NOR2_X2 U580 ( .A1(n536), .A2(n535), .ZN(G160) );
  INV_X1 U581 ( .A(G2105), .ZN(n525) );
  AND2_X2 U582 ( .A1(n525), .A2(G2104), .ZN(n537) );
  NAND2_X1 U583 ( .A1(G101), .A2(n537), .ZN(n527) );
  XOR2_X1 U584 ( .A(KEYINPUT17), .B(n528), .Z(n538) );
  BUF_X2 U585 ( .A(n538), .Z(n912) );
  NAND2_X1 U586 ( .A1(G137), .A2(n912), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n536) );
  INV_X1 U588 ( .A(G2104), .ZN(n531) );
  AND2_X1 U589 ( .A1(n531), .A2(G2105), .ZN(n908) );
  NAND2_X1 U590 ( .A1(G125), .A2(n908), .ZN(n534) );
  NAND2_X1 U591 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  XOR2_X1 U592 ( .A(n532), .B(KEYINPUT66), .Z(n541) );
  BUF_X2 U593 ( .A(n541), .Z(n906) );
  NAND2_X1 U594 ( .A1(G113), .A2(n906), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U596 ( .A1(G102), .A2(n537), .ZN(n540) );
  NAND2_X1 U597 ( .A1(G138), .A2(n538), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G126), .A2(n908), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G114), .A2(n541), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U602 ( .A1(n545), .A2(n544), .ZN(G164) );
  XNOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n546), .B(KEYINPUT67), .ZN(n600) );
  NAND2_X1 U605 ( .A1(n816), .A2(G47), .ZN(n550) );
  NOR2_X1 U606 ( .A1(G543), .A2(n522), .ZN(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT1), .B(n547), .Z(n685) );
  NAND2_X1 U608 ( .A1(G60), .A2(n548), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U610 ( .A(n551), .B(KEYINPUT71), .ZN(n557) );
  NOR2_X2 U611 ( .A1(n600), .A2(n522), .ZN(n810) );
  NAND2_X1 U612 ( .A1(G72), .A2(n810), .ZN(n552) );
  XOR2_X1 U613 ( .A(KEYINPUT69), .B(n552), .Z(n554) );
  NOR2_X1 U614 ( .A1(G651), .A2(G543), .ZN(n809) );
  NAND2_X1 U615 ( .A1(n809), .A2(G85), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT70), .B(n555), .Z(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n558), .B(KEYINPUT72), .ZN(G290) );
  XOR2_X1 U620 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n560) );
  NAND2_X1 U621 ( .A1(G73), .A2(n810), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n560), .B(n559), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n809), .A2(G86), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G61), .A2(n548), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G48), .A2(n816), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT85), .B(n565), .Z(n566) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(G305) );
  NAND2_X1 U630 ( .A1(n816), .A2(G52), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G64), .A2(n548), .ZN(n568) );
  NAND2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G90), .A2(n809), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G77), .A2(n810), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n572), .Z(n573) );
  NOR2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT73), .B(n575), .Z(G171) );
  NAND2_X1 U639 ( .A1(n816), .A2(G51), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G63), .A2(n548), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT6), .B(n578), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n809), .A2(G89), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT4), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G76), .A2(n810), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n582), .B(KEYINPUT5), .Z(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT7), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(KEYINPUT78), .B(n586), .ZN(G168) );
  NAND2_X1 U651 ( .A1(n816), .A2(G53), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G78), .A2(n810), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n809), .A2(G91), .ZN(n589) );
  XOR2_X1 U655 ( .A(KEYINPUT74), .B(n589), .Z(n590) );
  NOR2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G65), .A2(n548), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(G299) );
  XOR2_X1 U659 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U660 ( .A1(G88), .A2(n809), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G75), .A2(n810), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n816), .A2(G50), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G62), .A2(n548), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U666 ( .A1(n599), .A2(n598), .ZN(G166) );
  INV_X1 U667 ( .A(G166), .ZN(G303) );
  NAND2_X1 U668 ( .A1(G87), .A2(n600), .ZN(n602) );
  NAND2_X1 U669 ( .A1(G74), .A2(G651), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U671 ( .A1(n548), .A2(n603), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n816), .A2(G49), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(G288) );
  NOR2_X1 U674 ( .A1(n653), .A2(n651), .ZN(n606) );
  XNOR2_X1 U675 ( .A(KEYINPUT88), .B(n606), .ZN(n648) );
  INV_X1 U676 ( .A(n648), .ZN(n643) );
  NAND2_X1 U677 ( .A1(G128), .A2(n908), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G116), .A2(n906), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT35), .ZN(n615) );
  NAND2_X1 U681 ( .A1(n912), .A2(G140), .ZN(n610) );
  XOR2_X1 U682 ( .A(KEYINPUT89), .B(n610), .Z(n612) );
  NAND2_X1 U683 ( .A1(n537), .A2(G104), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U685 ( .A(KEYINPUT34), .B(n613), .Z(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n616), .B(KEYINPUT36), .ZN(n922) );
  XOR2_X1 U688 ( .A(G2067), .B(KEYINPUT37), .Z(n639) );
  NOR2_X1 U689 ( .A1(n922), .A2(n639), .ZN(n936) );
  NAND2_X1 U690 ( .A1(n908), .A2(G129), .ZN(n617) );
  XOR2_X1 U691 ( .A(KEYINPUT91), .B(n617), .Z(n619) );
  NAND2_X1 U692 ( .A1(G117), .A2(n906), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U694 ( .A(KEYINPUT92), .B(n620), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n537), .A2(G105), .ZN(n621) );
  XOR2_X1 U696 ( .A(KEYINPUT38), .B(n621), .Z(n622) );
  NOR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n912), .A2(G141), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n902) );
  NOR2_X1 U700 ( .A1(G1996), .A2(n902), .ZN(n933) );
  NAND2_X1 U701 ( .A1(G95), .A2(n537), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G131), .A2(n912), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U704 ( .A(KEYINPUT90), .B(n628), .Z(n632) );
  NAND2_X1 U705 ( .A1(n906), .A2(G107), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G119), .A2(n908), .ZN(n629) );
  AND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n918) );
  AND2_X1 U709 ( .A1(n918), .A2(G1991), .ZN(n634) );
  AND2_X1 U710 ( .A1(n902), .A2(G1996), .ZN(n633) );
  NOR2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n941) );
  NOR2_X1 U712 ( .A1(n643), .A2(n941), .ZN(n646) );
  NOR2_X1 U713 ( .A1(G1986), .A2(G290), .ZN(n635) );
  NOR2_X1 U714 ( .A1(G1991), .A2(n918), .ZN(n937) );
  NOR2_X1 U715 ( .A1(n635), .A2(n937), .ZN(n636) );
  NOR2_X1 U716 ( .A1(n646), .A2(n636), .ZN(n637) );
  NOR2_X1 U717 ( .A1(n933), .A2(n637), .ZN(n638) );
  XOR2_X1 U718 ( .A(KEYINPUT39), .B(n638), .Z(n640) );
  NAND2_X1 U719 ( .A1(n922), .A2(n639), .ZN(n951) );
  NOR2_X1 U720 ( .A1(n643), .A2(n951), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n640), .A2(n645), .ZN(n641) );
  NOR2_X1 U722 ( .A1(n936), .A2(n641), .ZN(n642) );
  NOR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(KEYINPUT104), .ZN(n772) );
  OR2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U726 ( .A(n647), .B(KEYINPUT93), .ZN(n650) );
  XNOR2_X1 U727 ( .A(G1986), .B(G290), .ZN(n992) );
  NAND2_X1 U728 ( .A1(n648), .A2(n992), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n770) );
  INV_X1 U730 ( .A(n651), .ZN(n652) );
  NOR2_X2 U731 ( .A1(n653), .A2(n652), .ZN(n665) );
  NAND2_X1 U732 ( .A1(G8), .A2(n723), .ZN(n754) );
  NOR2_X1 U733 ( .A1(G1981), .A2(G305), .ZN(n654) );
  XOR2_X1 U734 ( .A(n654), .B(KEYINPUT24), .Z(n655) );
  NOR2_X1 U735 ( .A1(n754), .A2(n655), .ZN(n768) );
  INV_X1 U736 ( .A(G1961), .ZN(n986) );
  NAND2_X1 U737 ( .A1(n723), .A2(n986), .ZN(n658) );
  BUF_X1 U738 ( .A(n665), .Z(n656) );
  XNOR2_X1 U739 ( .A(G2078), .B(KEYINPUT25), .ZN(n961) );
  NAND2_X1 U740 ( .A1(n656), .A2(n961), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n658), .A2(n657), .ZN(n715) );
  NOR2_X1 U742 ( .A1(G171), .A2(n715), .ZN(n663) );
  NOR2_X1 U743 ( .A1(G1966), .A2(n754), .ZN(n735) );
  NOR2_X1 U744 ( .A1(G2084), .A2(n723), .ZN(n733) );
  NOR2_X1 U745 ( .A1(n735), .A2(n733), .ZN(n659) );
  NAND2_X1 U746 ( .A1(G8), .A2(n659), .ZN(n660) );
  XNOR2_X1 U747 ( .A(KEYINPUT30), .B(n660), .ZN(n661) );
  NOR2_X1 U748 ( .A1(n661), .A2(G168), .ZN(n662) );
  NOR2_X1 U749 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U750 ( .A(KEYINPUT31), .B(n664), .ZN(n720) );
  XNOR2_X1 U751 ( .A(n667), .B(n666), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n723), .A2(G1341), .ZN(n668) );
  NAND2_X1 U753 ( .A1(n669), .A2(n668), .ZN(n682) );
  NAND2_X1 U754 ( .A1(n685), .A2(G56), .ZN(n670) );
  XNOR2_X1 U755 ( .A(n670), .B(KEYINPUT14), .ZN(n672) );
  INV_X1 U756 ( .A(KEYINPUT75), .ZN(n671) );
  XNOR2_X1 U757 ( .A(n672), .B(n671), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n809), .A2(G81), .ZN(n673) );
  XNOR2_X1 U759 ( .A(n673), .B(KEYINPUT12), .ZN(n675) );
  NAND2_X1 U760 ( .A1(G68), .A2(n810), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n676), .B(KEYINPUT13), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G43), .A2(n816), .ZN(n677) );
  AND2_X1 U764 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n680), .A2(n679), .ZN(n681) );
  INV_X1 U766 ( .A(KEYINPUT64), .ZN(n683) );
  XNOR2_X1 U767 ( .A(n684), .B(n683), .ZN(n698) );
  NAND2_X1 U768 ( .A1(n809), .A2(G92), .ZN(n687) );
  NAND2_X1 U769 ( .A1(G66), .A2(n685), .ZN(n686) );
  NAND2_X1 U770 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U771 ( .A1(n816), .A2(G54), .ZN(n690) );
  NAND2_X1 U772 ( .A1(G79), .A2(n810), .ZN(n689) );
  XNOR2_X1 U773 ( .A(KEYINPUT15), .B(n692), .ZN(n1000) );
  OR2_X1 U774 ( .A1(n698), .A2(n1000), .ZN(n697) );
  AND2_X1 U775 ( .A1(n656), .A2(G2067), .ZN(n693) );
  XOR2_X1 U776 ( .A(n693), .B(KEYINPUT96), .Z(n695) );
  NAND2_X1 U777 ( .A1(n723), .A2(G1348), .ZN(n694) );
  NAND2_X1 U778 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U779 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U780 ( .A1(n698), .A2(n1000), .ZN(n699) );
  NAND2_X1 U781 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U782 ( .A(n702), .B(n701), .ZN(n707) );
  NAND2_X1 U783 ( .A1(n656), .A2(G2072), .ZN(n703) );
  XNOR2_X1 U784 ( .A(n703), .B(KEYINPUT27), .ZN(n705) );
  AND2_X1 U785 ( .A1(G1956), .A2(n723), .ZN(n704) );
  NOR2_X1 U786 ( .A1(n705), .A2(n704), .ZN(n708) );
  INV_X1 U787 ( .A(G299), .ZN(n824) );
  NAND2_X1 U788 ( .A1(n708), .A2(n824), .ZN(n706) );
  NAND2_X1 U789 ( .A1(n707), .A2(n706), .ZN(n713) );
  NOR2_X1 U790 ( .A1(n708), .A2(n824), .ZN(n711) );
  XNOR2_X1 U791 ( .A(KEYINPUT28), .B(KEYINPUT95), .ZN(n709) );
  XNOR2_X1 U792 ( .A(n709), .B(KEYINPUT94), .ZN(n710) );
  XNOR2_X1 U793 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U795 ( .A(n714), .B(KEYINPUT29), .ZN(n717) );
  AND2_X1 U796 ( .A1(G171), .A2(n715), .ZN(n716) );
  NOR2_X1 U797 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U798 ( .A(KEYINPUT98), .B(n718), .ZN(n719) );
  XNOR2_X1 U799 ( .A(n721), .B(KEYINPUT99), .ZN(n737) );
  AND2_X1 U800 ( .A1(G286), .A2(G8), .ZN(n722) );
  NAND2_X1 U801 ( .A1(n737), .A2(n722), .ZN(n730) );
  INV_X1 U802 ( .A(G8), .ZN(n728) );
  NOR2_X1 U803 ( .A1(G1971), .A2(n754), .ZN(n725) );
  NOR2_X1 U804 ( .A1(G2090), .A2(n723), .ZN(n724) );
  NOR2_X1 U805 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U806 ( .A1(n726), .A2(G303), .ZN(n727) );
  OR2_X1 U807 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U808 ( .A1(n730), .A2(n729), .ZN(n732) );
  AND2_X1 U809 ( .A1(G8), .A2(n733), .ZN(n734) );
  NOR2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U811 ( .A1(n737), .A2(n736), .ZN(n739) );
  INV_X1 U812 ( .A(KEYINPUT100), .ZN(n738) );
  XNOR2_X1 U813 ( .A(n739), .B(n738), .ZN(n755) );
  NAND2_X1 U814 ( .A1(G1976), .A2(G288), .ZN(n995) );
  INV_X1 U815 ( .A(n754), .ZN(n760) );
  NAND2_X1 U816 ( .A1(n995), .A2(n760), .ZN(n747) );
  INV_X1 U817 ( .A(n747), .ZN(n742) );
  NOR2_X1 U818 ( .A1(G1976), .A2(G288), .ZN(n746) );
  NAND2_X1 U819 ( .A1(n746), .A2(KEYINPUT33), .ZN(n740) );
  NOR2_X1 U820 ( .A1(n740), .A2(n754), .ZN(n750) );
  INV_X1 U821 ( .A(n750), .ZN(n741) );
  NAND2_X1 U822 ( .A1(n757), .A2(n744), .ZN(n752) );
  NOR2_X1 U823 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U824 ( .A1(n746), .A2(n745), .ZN(n996) );
  NOR2_X1 U825 ( .A1(n747), .A2(n996), .ZN(n748) );
  NOR2_X1 U826 ( .A1(n748), .A2(KEYINPUT33), .ZN(n749) );
  OR2_X1 U827 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U829 ( .A(G1981), .B(G305), .Z(n981) );
  NAND2_X1 U830 ( .A1(n753), .A2(n981), .ZN(n764) );
  AND2_X1 U831 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n762) );
  NOR2_X1 U833 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U834 ( .A1(G8), .A2(n758), .ZN(n759) );
  OR2_X1 U835 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n764), .A2(n763), .ZN(n766) );
  XNOR2_X1 U838 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U839 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U840 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U841 ( .A1(n772), .A2(n771), .ZN(n774) );
  XNOR2_X1 U842 ( .A(n774), .B(n773), .ZN(G329) );
  INV_X1 U843 ( .A(G171), .ZN(G301) );
  XOR2_X1 U844 ( .A(G2438), .B(G2454), .Z(n776) );
  XNOR2_X1 U845 ( .A(G2435), .B(G2430), .ZN(n775) );
  XNOR2_X1 U846 ( .A(n776), .B(n775), .ZN(n777) );
  XOR2_X1 U847 ( .A(n777), .B(KEYINPUT106), .Z(n779) );
  XNOR2_X1 U848 ( .A(G1341), .B(G1348), .ZN(n778) );
  XNOR2_X1 U849 ( .A(n779), .B(n778), .ZN(n783) );
  XOR2_X1 U850 ( .A(G2446), .B(G2451), .Z(n781) );
  XNOR2_X1 U851 ( .A(G2443), .B(G2427), .ZN(n780) );
  XNOR2_X1 U852 ( .A(n781), .B(n780), .ZN(n782) );
  XOR2_X1 U853 ( .A(n783), .B(n782), .Z(n784) );
  AND2_X1 U854 ( .A1(G14), .A2(n784), .ZN(G401) );
  AND2_X1 U855 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U856 ( .A1(G123), .A2(n908), .ZN(n785) );
  XNOR2_X1 U857 ( .A(n785), .B(KEYINPUT18), .ZN(n787) );
  NAND2_X1 U858 ( .A1(n537), .A2(G99), .ZN(n786) );
  NAND2_X1 U859 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U860 ( .A1(G135), .A2(n912), .ZN(n789) );
  NAND2_X1 U861 ( .A1(G111), .A2(n906), .ZN(n788) );
  NAND2_X1 U862 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U863 ( .A1(n791), .A2(n790), .ZN(n938) );
  XNOR2_X1 U864 ( .A(n938), .B(G2096), .ZN(n792) );
  XNOR2_X1 U865 ( .A(n792), .B(KEYINPUT81), .ZN(n793) );
  OR2_X1 U866 ( .A1(G2100), .A2(n793), .ZN(G156) );
  INV_X1 U867 ( .A(G57), .ZN(G237) );
  NAND2_X1 U868 ( .A1(G7), .A2(G661), .ZN(n794) );
  XOR2_X1 U869 ( .A(n794), .B(KEYINPUT10), .Z(n848) );
  NAND2_X1 U870 ( .A1(n848), .A2(G567), .ZN(n795) );
  XOR2_X1 U871 ( .A(KEYINPUT11), .B(n795), .Z(G234) );
  INV_X1 U872 ( .A(G860), .ZN(n802) );
  OR2_X1 U873 ( .A1(n802), .A2(n984), .ZN(G153) );
  NAND2_X1 U874 ( .A1(G868), .A2(G301), .ZN(n798) );
  INV_X1 U875 ( .A(G868), .ZN(n832) );
  NAND2_X1 U876 ( .A1(n1000), .A2(n832), .ZN(n797) );
  NAND2_X1 U877 ( .A1(n798), .A2(n797), .ZN(G284) );
  NOR2_X1 U878 ( .A1(G286), .A2(n832), .ZN(n799) );
  XOR2_X1 U879 ( .A(KEYINPUT79), .B(n799), .Z(n801) );
  NOR2_X1 U880 ( .A1(G868), .A2(G299), .ZN(n800) );
  NOR2_X1 U881 ( .A1(n801), .A2(n800), .ZN(G297) );
  NAND2_X1 U882 ( .A1(n802), .A2(G559), .ZN(n803) );
  INV_X1 U883 ( .A(n1000), .ZN(n855) );
  NAND2_X1 U884 ( .A1(n803), .A2(n855), .ZN(n804) );
  XNOR2_X1 U885 ( .A(n804), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U886 ( .A1(n984), .A2(G868), .ZN(n807) );
  NAND2_X1 U887 ( .A1(G868), .A2(n855), .ZN(n805) );
  NOR2_X1 U888 ( .A1(G559), .A2(n805), .ZN(n806) );
  NOR2_X1 U889 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U890 ( .A(KEYINPUT80), .B(n808), .ZN(G282) );
  NAND2_X1 U891 ( .A1(G93), .A2(n809), .ZN(n812) );
  NAND2_X1 U892 ( .A1(G80), .A2(n810), .ZN(n811) );
  NAND2_X1 U893 ( .A1(n812), .A2(n811), .ZN(n815) );
  NAND2_X1 U894 ( .A1(n548), .A2(G67), .ZN(n813) );
  XOR2_X1 U895 ( .A(KEYINPUT82), .B(n813), .Z(n814) );
  NOR2_X1 U896 ( .A1(n815), .A2(n814), .ZN(n818) );
  NAND2_X1 U897 ( .A1(n816), .A2(G55), .ZN(n817) );
  NAND2_X1 U898 ( .A1(n818), .A2(n817), .ZN(n831) );
  NAND2_X1 U899 ( .A1(G559), .A2(n855), .ZN(n819) );
  XNOR2_X1 U900 ( .A(n819), .B(n984), .ZN(n828) );
  NOR2_X1 U901 ( .A1(G860), .A2(n828), .ZN(n820) );
  XNOR2_X1 U902 ( .A(n820), .B(KEYINPUT83), .ZN(n821) );
  XNOR2_X1 U903 ( .A(n831), .B(n821), .ZN(G145) );
  XNOR2_X1 U904 ( .A(KEYINPUT19), .B(G288), .ZN(n822) );
  XNOR2_X1 U905 ( .A(n822), .B(n831), .ZN(n823) );
  XOR2_X1 U906 ( .A(n823), .B(G290), .Z(n826) );
  XOR2_X1 U907 ( .A(G303), .B(n824), .Z(n825) );
  XNOR2_X1 U908 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U909 ( .A(n827), .B(G305), .ZN(n854) );
  XNOR2_X1 U910 ( .A(n854), .B(n828), .ZN(n829) );
  NAND2_X1 U911 ( .A1(n829), .A2(G868), .ZN(n830) );
  XNOR2_X1 U912 ( .A(n830), .B(KEYINPUT86), .ZN(n834) );
  NAND2_X1 U913 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U914 ( .A1(n834), .A2(n833), .ZN(G295) );
  NAND2_X1 U915 ( .A1(G2084), .A2(G2078), .ZN(n835) );
  XOR2_X1 U916 ( .A(KEYINPUT20), .B(n835), .Z(n836) );
  NAND2_X1 U917 ( .A1(G2090), .A2(n836), .ZN(n837) );
  XNOR2_X1 U918 ( .A(KEYINPUT21), .B(n837), .ZN(n838) );
  NAND2_X1 U919 ( .A1(n838), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U920 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U921 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n840) );
  NAND2_X1 U922 ( .A1(G132), .A2(G82), .ZN(n839) );
  XNOR2_X1 U923 ( .A(n840), .B(n839), .ZN(n841) );
  NOR2_X1 U924 ( .A1(n841), .A2(G218), .ZN(n842) );
  NAND2_X1 U925 ( .A1(G96), .A2(n842), .ZN(n852) );
  NAND2_X1 U926 ( .A1(n852), .A2(G2106), .ZN(n846) );
  NAND2_X1 U927 ( .A1(G69), .A2(G120), .ZN(n843) );
  NOR2_X1 U928 ( .A1(G237), .A2(n843), .ZN(n844) );
  NAND2_X1 U929 ( .A1(G108), .A2(n844), .ZN(n853) );
  NAND2_X1 U930 ( .A1(n853), .A2(G567), .ZN(n845) );
  NAND2_X1 U931 ( .A1(n846), .A2(n845), .ZN(n930) );
  NAND2_X1 U932 ( .A1(G483), .A2(G661), .ZN(n847) );
  NOR2_X1 U933 ( .A1(n930), .A2(n847), .ZN(n851) );
  NAND2_X1 U934 ( .A1(n851), .A2(G36), .ZN(G176) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n848), .ZN(G217) );
  INV_X1 U936 ( .A(n848), .ZN(G223) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n849) );
  NAND2_X1 U938 ( .A1(G661), .A2(n849), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U940 ( .A1(n851), .A2(n850), .ZN(G188) );
  INV_X1 U942 ( .A(G132), .ZN(G219) );
  INV_X1 U943 ( .A(G120), .ZN(G236) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  INV_X1 U945 ( .A(G82), .ZN(G220) );
  INV_X1 U946 ( .A(G69), .ZN(G235) );
  NOR2_X1 U947 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  XOR2_X1 U949 ( .A(n854), .B(n984), .Z(n857) );
  XOR2_X1 U950 ( .A(G301), .B(n855), .Z(n856) );
  XNOR2_X1 U951 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U952 ( .A(n858), .B(G286), .ZN(n859) );
  NOR2_X1 U953 ( .A1(G37), .A2(n859), .ZN(G397) );
  XOR2_X1 U954 ( .A(KEYINPUT111), .B(G1991), .Z(n862) );
  INV_X1 U955 ( .A(G1996), .ZN(n860) );
  XOR2_X1 U956 ( .A(n860), .B(G1986), .Z(n861) );
  XNOR2_X1 U957 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U958 ( .A(n863), .B(KEYINPUT41), .Z(n865) );
  XNOR2_X1 U959 ( .A(G1971), .B(G1976), .ZN(n864) );
  XNOR2_X1 U960 ( .A(n865), .B(n864), .ZN(n869) );
  XNOR2_X1 U961 ( .A(G1956), .B(n986), .ZN(n867) );
  XNOR2_X1 U962 ( .A(G1981), .B(G1966), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U964 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U965 ( .A(KEYINPUT110), .B(G2474), .ZN(n870) );
  XNOR2_X1 U966 ( .A(n871), .B(n870), .ZN(G229) );
  XNOR2_X1 U967 ( .A(G2072), .B(G2067), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n872), .B(KEYINPUT42), .ZN(n882) );
  XOR2_X1 U969 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n874) );
  XNOR2_X1 U970 ( .A(KEYINPUT108), .B(G2096), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U972 ( .A(G2100), .B(G2078), .Z(n876) );
  XNOR2_X1 U973 ( .A(G2090), .B(G2084), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U975 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U976 ( .A(KEYINPUT109), .B(G2678), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(G227) );
  NAND2_X1 U979 ( .A1(G124), .A2(n908), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n883), .B(KEYINPUT44), .ZN(n885) );
  NAND2_X1 U981 ( .A1(n537), .A2(G100), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G136), .A2(n912), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G112), .A2(n906), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n888) );
  NOR2_X1 U986 ( .A1(n889), .A2(n888), .ZN(G162) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n891) );
  XNOR2_X1 U988 ( .A(G164), .B(KEYINPUT114), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(n892), .B(n938), .Z(n894) );
  XNOR2_X1 U991 ( .A(G160), .B(G162), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n905) );
  NAND2_X1 U993 ( .A1(G130), .A2(n908), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G118), .A2(n906), .ZN(n895) );
  NAND2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n901) );
  NAND2_X1 U996 ( .A1(G106), .A2(n537), .ZN(n898) );
  NAND2_X1 U997 ( .A1(G142), .A2(n912), .ZN(n897) );
  NAND2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U999 ( .A(n899), .B(KEYINPUT45), .Z(n900) );
  NOR2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1002 ( .A(n905), .B(n904), .Z(n920) );
  NAND2_X1 U1003 ( .A1(G115), .A2(n906), .ZN(n907) );
  XOR2_X1 U1004 ( .A(KEYINPUT113), .B(n907), .Z(n910) );
  NAND2_X1 U1005 ( .A1(n908), .A2(G127), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n911), .B(KEYINPUT47), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(G139), .A2(n912), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n917) );
  NAND2_X1 U1010 ( .A1(n537), .A2(G103), .ZN(n915) );
  XOR2_X1 U1011 ( .A(KEYINPUT112), .B(n915), .Z(n916) );
  NOR2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n947) );
  XOR2_X1 U1013 ( .A(n918), .B(n947), .Z(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1015 ( .A(n922), .B(n921), .Z(n923) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n923), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G229), .A2(G227), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n924), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G397), .A2(n925), .ZN(n929) );
  NOR2_X1 U1020 ( .A1(G401), .A2(n930), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(KEYINPUT115), .B(n926), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(G395), .A2(n927), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(n930), .ZN(G319) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n931) );
  XNOR2_X1 U1028 ( .A(KEYINPUT118), .B(n931), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(KEYINPUT51), .B(n934), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n946) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT117), .B(n939), .Z(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n944) );
  XOR2_X1 U1035 ( .A(G2084), .B(G160), .Z(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT116), .B(n942), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n954) );
  XOR2_X1 U1039 ( .A(G2072), .B(n947), .Z(n949) );
  XOR2_X1 U1040 ( .A(G164), .B(G2078), .Z(n948) );
  NOR2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(n950), .B(KEYINPUT50), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(n955), .ZN(n956) );
  INV_X1 U1046 ( .A(KEYINPUT55), .ZN(n1030) );
  NAND2_X1 U1047 ( .A1(n956), .A2(n1030), .ZN(n957) );
  NAND2_X1 U1048 ( .A1(n957), .A2(G29), .ZN(n1039) );
  XNOR2_X1 U1049 ( .A(KEYINPUT119), .B(G2090), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(n958), .B(G35), .ZN(n977) );
  XOR2_X1 U1051 ( .A(G1991), .B(G25), .Z(n959) );
  NAND2_X1 U1052 ( .A1(n959), .A2(G28), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(KEYINPUT120), .ZN(n970) );
  XOR2_X1 U1054 ( .A(G32), .B(G1996), .Z(n968) );
  XOR2_X1 U1055 ( .A(n961), .B(G27), .Z(n966) );
  XNOR2_X1 U1056 ( .A(G2072), .B(G33), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT121), .B(n964), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(KEYINPUT122), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n972), .B(n971), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(G2084), .B(G34), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n973), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n1031) );
  NOR2_X1 U1069 ( .A1(G29), .A2(KEYINPUT55), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n1031), .A2(n978), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n979), .ZN(n1037) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .ZN(n1006) );
  XOR2_X1 U1073 ( .A(G1966), .B(KEYINPUT123), .Z(n980) );
  XNOR2_X1 U1074 ( .A(G168), .B(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT57), .ZN(n990) );
  XOR2_X1 U1077 ( .A(n984), .B(G1341), .Z(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT125), .B(n985), .ZN(n988) );
  XOR2_X1 U1079 ( .A(n986), .B(G301), .Z(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n1004) );
  XOR2_X1 U1083 ( .A(G1956), .B(G299), .Z(n994) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT124), .B(n999), .Z(n1002) );
  XNOR2_X1 U1089 ( .A(G1348), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(KEYINPUT126), .B(n1007), .ZN(n1035) );
  XOR2_X1 U1094 ( .A(G5), .B(G1961), .Z(n1020) );
  XNOR2_X1 U1095 ( .A(G1348), .B(KEYINPUT59), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1008), .B(G4), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1981), .B(G6), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G20), .B(G1956), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(G19), .B(G1341), .Z(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1016), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G21), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XNOR2_X1 U1108 ( .A(G1971), .B(G22), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(G24), .B(G1986), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1111 ( .A(G1976), .B(G23), .Z(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1028), .Z(n1029) );
  NOR2_X1 U1116 ( .A1(G16), .A2(n1029), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1121 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1040), .ZN(G150) );
  INV_X1 U1123 ( .A(G150), .ZN(G311) );
endmodule

