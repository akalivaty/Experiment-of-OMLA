//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G221), .A2(G220), .A3(G219), .A4(G218), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n466), .A2(new_n469), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT68), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G113), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(new_n463), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n476), .A2(KEYINPUT68), .A3(new_n477), .ZN(new_n481));
  OAI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND3_X1  g059(.A1(new_n467), .A2(G2105), .A3(new_n471), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT70), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT71), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(G136), .B2(new_n473), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n467), .A2(new_n471), .ZN(new_n496));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n466), .A2(new_n469), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n468), .A2(G138), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n497), .A2(new_n495), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n502), .B1(KEYINPUT73), .B2(new_n506), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(new_n504), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n498), .B(new_n507), .C1(new_n510), .C2(new_n496), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT5), .B(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n519), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n515), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(new_n518), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n522), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n521), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n518), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n523), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n515), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n540), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(new_n518), .A2(G43), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n521), .A2(new_n522), .A3(G81), .ZN(new_n546));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n522), .B2(G56), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n545), .B(new_n546), .C1(new_n548), .C2(new_n515), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  XNOR2_X1  g130(.A(new_n522), .B(KEYINPUT74), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(G78), .A2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OR3_X1    g136(.A1(new_n530), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n530), .B2(new_n561), .ZN(new_n563));
  AND2_X1   g138(.A1(KEYINPUT5), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(KEYINPUT5), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n565), .A2(new_n567), .B1(new_n516), .B2(new_n517), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n562), .A2(new_n563), .B1(G91), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n560), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  OAI21_X1  g147(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n573));
  INV_X1    g148(.A(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n530), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n568), .A2(G87), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT75), .ZN(G288));
  NAND2_X1  g153(.A1(new_n522), .A2(G61), .ZN(new_n579));
  INV_X1    g154(.A(G73), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n580), .B2(new_n513), .ZN(new_n581));
  OR3_X1    g156(.A1(new_n580), .A2(new_n513), .A3(KEYINPUT76), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(G48), .B2(new_n518), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n523), .ZN(G305));
  NAND2_X1  g161(.A1(new_n518), .A2(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(new_n523), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n515), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n556), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g171(.A1(G79), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n523), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n568), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n601), .A2(new_n602), .B1(G54), .B2(new_n518), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n594), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n594), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n608), .B2(G168), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n608), .B2(G168), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n502), .A2(new_n474), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT13), .B(G2100), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n486), .A2(G123), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(G111), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G2105), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n473), .B2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n622), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT83), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(KEYINPUT17), .ZN(new_n661));
  INV_X1    g236(.A(new_n655), .ZN(new_n662));
  INV_X1    g237(.A(new_n656), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n658), .A3(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(new_n657), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n671), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n671), .B2(new_n677), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT84), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  MUX2_X1   g262(.A(G6), .B(G305), .S(G16), .Z(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT32), .B(G1981), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1971), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(G23), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n577), .B2(new_n691), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT33), .B(G1976), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n690), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  OR2_X1    g279(.A1(G95), .A2(G2105), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n705), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n706));
  INV_X1    g281(.A(G119), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n485), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G131), .B2(new_n473), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  AOI21_X1  g287(.A(new_n691), .B1(G290), .B2(KEYINPUT86), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(KEYINPUT86), .B2(G290), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n691), .A2(G24), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT85), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n712), .B(new_n718), .C1(new_n699), .C2(new_n700), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n702), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT89), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n691), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n691), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G1966), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT96), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n691), .A2(G5), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G171), .B2(new_n691), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G1961), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G1966), .B2(new_n725), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT30), .B(G28), .Z(new_n733));
  OAI221_X1 g308(.A(new_n732), .B1(G29), .B2(new_n733), .C1(new_n729), .C2(G1961), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G19), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n550), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1341), .ZN(new_n737));
  OR3_X1    g312(.A1(new_n731), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2078), .ZN(new_n739));
  NOR2_X1   g314(.A1(G164), .A2(new_n703), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G27), .B2(new_n703), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n727), .B(new_n738), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n691), .A2(G20), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G299), .B2(G16), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT99), .B(G1956), .Z(new_n746));
  XOR2_X1   g321(.A(new_n745), .B(new_n746), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n703), .A2(G32), .ZN(new_n748));
  INV_X1    g323(.A(G141), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n472), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT94), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT95), .B(KEYINPUT26), .Z(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n474), .A2(G105), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G129), .B2(new_n486), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n751), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n748), .B1(new_n759), .B2(new_n703), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT27), .B(G1996), .Z(new_n761));
  XOR2_X1   g336(.A(new_n760), .B(new_n761), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n631), .A2(G29), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G4), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n605), .B2(G16), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n741), .A2(new_n739), .B1(new_n767), .B2(G1348), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n765), .B(new_n768), .C1(G1348), .C2(new_n767), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n742), .A2(new_n747), .A3(new_n762), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n703), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n703), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G2090), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT98), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n703), .A2(G33), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT25), .Z(new_n778));
  INV_X1    g353(.A(G139), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n502), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n778), .B1(new_n472), .B2(new_n779), .C1(new_n468), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT92), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(new_n703), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT93), .B(G2072), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(G34), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n703), .B1(new_n786), .B2(G34), .ZN(new_n788));
  OAI22_X1  g363(.A1(new_n483), .A2(new_n703), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2084), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n764), .B2(new_n763), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n703), .A2(G26), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT28), .ZN(new_n794));
  INV_X1    g369(.A(G128), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n468), .A2(G116), .ZN(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n485), .A2(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G140), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n472), .A2(KEYINPUT90), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(KEYINPUT90), .B1(new_n472), .B2(new_n799), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n794), .B1(new_n802), .B2(new_n703), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT91), .B(G2067), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n785), .A2(new_n792), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n773), .A2(G2090), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n770), .A2(new_n775), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n723), .A2(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  NAND3_X1  g385(.A1(new_n521), .A2(G55), .A3(G543), .ZN(new_n811));
  INV_X1    g386(.A(G93), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n523), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT100), .ZN(new_n814));
  NAND2_X1  g389(.A1(G80), .A2(G543), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n522), .B2(G67), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n814), .B1(new_n817), .B2(new_n515), .ZN(new_n818));
  OAI21_X1  g393(.A(G67), .B1(new_n564), .B2(new_n566), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n815), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n820), .A2(KEYINPUT100), .A3(G651), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n813), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT103), .B(G860), .Z(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT37), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n605), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n822), .B2(new_n549), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n568), .A2(G93), .B1(new_n518), .B2(G55), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT100), .B1(new_n820), .B2(G651), .ZN(new_n831));
  AOI211_X1 g406(.A(new_n814), .B(new_n515), .C1(new_n819), .C2(new_n815), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(KEYINPUT101), .A3(new_n550), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n549), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT102), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n822), .A2(new_n838), .A3(new_n549), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n827), .B(new_n841), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n823), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n825), .B1(new_n844), .B2(new_n846), .ZN(G145));
  INV_X1    g422(.A(KEYINPUT106), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n782), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT92), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n781), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT106), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n798), .ZN(new_n854));
  INV_X1    g429(.A(new_n801), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n472), .A2(KEYINPUT90), .A3(new_n799), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n511), .ZN(new_n858));
  NAND2_X1  g433(.A1(G164), .A2(new_n802), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n758), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n758), .A2(new_n859), .A3(new_n858), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n853), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n864));
  OR2_X1    g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n866));
  INV_X1    g441(.A(G142), .ZN(new_n867));
  INV_X1    g442(.A(G130), .ZN(new_n868));
  OAI221_X1 g443(.A(new_n866), .B1(new_n472), .B2(new_n867), .C1(new_n868), .C2(new_n485), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n709), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n485), .B2(new_n868), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(G142), .B2(new_n473), .ZN(new_n872));
  INV_X1    g447(.A(G131), .ZN(new_n873));
  OAI221_X1 g448(.A(new_n706), .B1(new_n472), .B2(new_n873), .C1(new_n707), .C2(new_n485), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n870), .A2(new_n875), .A3(new_n620), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n620), .B1(new_n870), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n864), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(new_n875), .ZN(new_n879));
  INV_X1    g454(.A(new_n620), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n870), .A2(new_n875), .A3(new_n620), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(KEYINPUT107), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n862), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n852), .B1(new_n885), .B2(new_n860), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n863), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT108), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n863), .A2(new_n886), .ZN(new_n889));
  INV_X1    g464(.A(new_n884), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(KEYINPUT108), .A3(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n493), .A2(new_n630), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n488), .A2(new_n625), .A3(new_n492), .A4(new_n629), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n483), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n483), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n895), .A3(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n894), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n881), .A2(new_n882), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n889), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n909), .A3(new_n887), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(KEYINPUT109), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n905), .B1(new_n892), .B2(new_n893), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n911), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g494(.A(new_n614), .B(new_n841), .Z(new_n920));
  AOI22_X1  g495(.A1(new_n560), .A2(new_n569), .B1(new_n598), .B2(new_n603), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n560), .A2(new_n598), .A3(new_n569), .A4(new_n603), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT41), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  INV_X1    g500(.A(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n920), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n920), .B1(new_n921), .B2(new_n926), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  XNOR2_X1  g509(.A(G305), .B(new_n592), .ZN(new_n935));
  XOR2_X1   g510(.A(G166), .B(new_n577), .Z(new_n936));
  XOR2_X1   g511(.A(new_n935), .B(new_n936), .Z(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n933), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n930), .A2(new_n932), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(G868), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n822), .A2(G868), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(G295));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n944), .B2(new_n946), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n938), .B1(new_n933), .B2(new_n934), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n941), .A2(new_n937), .A3(new_n942), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n608), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n952), .A2(KEYINPUT110), .A3(new_n945), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n949), .A2(new_n953), .ZN(G331));
  NAND2_X1  g529(.A1(new_n841), .A2(G171), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n835), .A2(new_n840), .A3(G301), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(G168), .A3(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n835), .A2(new_n840), .A3(G301), .ZN(new_n958));
  AOI21_X1  g533(.A(G301), .B1(new_n835), .B2(new_n840), .ZN(new_n959));
  OAI21_X1  g534(.A(G286), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n928), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n926), .A2(new_n921), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n957), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n937), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n960), .A2(new_n957), .A3(KEYINPUT111), .A4(new_n963), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND4_X1   g545(.A1(KEYINPUT112), .A2(new_n970), .A3(new_n938), .A4(new_n962), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n961), .B1(new_n968), .B2(new_n969), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT112), .B1(new_n972), .B2(new_n938), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT43), .B(new_n966), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n911), .B1(new_n972), .B2(new_n938), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n970), .A2(new_n938), .A3(new_n962), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(KEYINPUT112), .A3(new_n938), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n974), .B1(new_n980), .B2(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT44), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(new_n966), .C1(new_n971), .C2(new_n973), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n987), .ZN(G397));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n758), .B(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n802), .B(G2067), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n709), .B(new_n711), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n592), .B(G1986), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n511), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n475), .A2(new_n482), .A3(G40), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(G171), .B2(KEYINPUT127), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1001), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1000), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n739), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n1011));
  INV_X1    g586(.A(G1961), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n511), .A2(new_n1014), .A3(new_n997), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1007), .A3(new_n1015), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1010), .A2(new_n1011), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1009), .A2(KEYINPUT53), .A3(new_n739), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(G301), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(G301), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1006), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n998), .A2(new_n1001), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n577), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1025), .B(new_n1027), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G305), .A2(G1981), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT115), .B(G86), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n568), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n584), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT116), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT116), .B(new_n1037), .C1(new_n1030), .C2(new_n1034), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1025), .A3(new_n1038), .ZN(new_n1039));
  OAI221_X1 g614(.A(G8), .B1(new_n1026), .B2(new_n1028), .C1(new_n998), .C2(new_n1001), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1029), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G166), .A2(new_n1024), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT55), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(KEYINPUT114), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(KEYINPUT114), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1043), .A2(KEYINPUT55), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1009), .A2(G1971), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT113), .B(G2090), .Z(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1016), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(G8), .B(new_n1048), .C1(new_n1049), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1049), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1015), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1013), .A2(new_n1056), .A3(new_n1007), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1014), .B1(new_n511), .B2(new_n997), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT118), .B1(new_n1058), .B2(new_n1001), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1050), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1024), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1042), .B(new_n1053), .C1(new_n1062), .C2(new_n1048), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G171), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(new_n1005), .A3(new_n1019), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G168), .A2(new_n1024), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT51), .B1(new_n1068), .B2(KEYINPUT126), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1016), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1000), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1072));
  INV_X1    g647(.A(G1966), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1071), .A2(new_n790), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1069), .B(new_n1070), .C1(new_n1074), .C2(new_n1024), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1070), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1013), .A2(new_n790), .A3(new_n1007), .A4(new_n1015), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1024), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1079), .B2(new_n1068), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1074), .A2(new_n1069), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1022), .A2(new_n1064), .A3(new_n1067), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  INV_X1    g660(.A(G2067), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1016), .A2(new_n1085), .B1(new_n1086), .B2(new_n1023), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(new_n604), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n998), .A2(new_n1001), .A3(G2067), .ZN(new_n1089));
  AOI211_X1 g664(.A(new_n605), .B(new_n1089), .C1(new_n1016), .C2(new_n1085), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT58), .B(G1341), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1072), .A2(G1996), .B1(new_n1023), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n550), .ZN(new_n1094));
  NOR2_X1   g669(.A1(KEYINPUT124), .A2(KEYINPUT59), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1094), .A2(new_n1095), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1091), .B(new_n1097), .C1(new_n1094), .C2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT120), .B(G1956), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT56), .B(G2072), .Z(new_n1101));
  OAI22_X1  g676(.A1(new_n1060), .A2(new_n1100), .B1(new_n1072), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G299), .A2(KEYINPUT121), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  OAI221_X1 g682(.A(new_n1105), .B1(new_n1072), .B2(new_n1101), .C1(new_n1060), .C2(new_n1100), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT61), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1099), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1072), .A2(new_n1101), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1056), .B1(new_n1013), .B2(new_n1007), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1058), .A2(KEYINPUT118), .A3(new_n1001), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1015), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1100), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1111), .B1(new_n1117), .B2(new_n1105), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1102), .A2(KEYINPUT123), .A3(new_n1106), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1108), .A2(KEYINPUT61), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT125), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1121), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1110), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1108), .B1(new_n1120), .B2(new_n1088), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1084), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1081), .A2(new_n1130), .A3(new_n1082), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1129), .A2(new_n1021), .A3(new_n1064), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1079), .A2(KEYINPUT119), .A3(G168), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT119), .B1(new_n1079), .B2(G168), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1063), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1042), .A2(new_n1053), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(G8), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1048), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1133), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1139), .B(new_n1142), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1053), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G288), .A2(G1976), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1039), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1030), .B(KEYINPUT117), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1145), .A2(new_n1042), .B1(new_n1149), .B2(new_n1025), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1132), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1003), .B1(new_n1128), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1002), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1153), .A2(G1986), .A3(G290), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT48), .Z(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1153), .B2(new_n994), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n709), .A2(new_n711), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n992), .A2(new_n1157), .B1(G2067), .B2(new_n857), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1002), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT47), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1153), .B1(new_n991), .B2(new_n759), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1002), .A2(KEYINPUT46), .A3(new_n989), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT46), .B1(new_n1002), .B2(new_n989), .ZN(new_n1163));
  OR3_X1    g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1156), .B(new_n1159), .C1(new_n1160), .C2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1152), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g742(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n985), .A2(new_n918), .A3(new_n1169), .ZN(G225));
  INV_X1    g744(.A(G225), .ZN(G308));
endmodule


