//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT79), .Z(new_n189));
  INV_X1    g003(.A(KEYINPUT81), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(new_n195), .A3(new_n191), .A4(G104), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n191), .A2(G104), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n193), .A2(new_n194), .A3(new_n196), .A4(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G107), .ZN(new_n201));
  OAI21_X1  g015(.A(G101), .B1(new_n201), .B2(new_n197), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n208), .A2(KEYINPUT66), .A3(new_n210), .A4(new_n212), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(G146), .B1(new_n205), .B2(new_n207), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g033(.A(G128), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n208), .A2(new_n210), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n203), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g037(.A1(new_n223), .A2(KEYINPUT10), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n193), .A2(new_n196), .A3(new_n198), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n209), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT64), .B(G143), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G146), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n204), .A2(G146), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n230), .B2(G146), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n231), .A2(new_n234), .B1(new_n236), .B2(new_n232), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n225), .A2(new_n238), .A3(G101), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n227), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT11), .B1(new_n241), .B2(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OR2_X1    g058(.A1(KEYINPUT65), .A2(G137), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT65), .A2(G137), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT11), .A2(G134), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n244), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n244), .B2(new_n248), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(G128), .B1(new_n235), .B2(new_n219), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(KEYINPUT67), .C1(new_n218), .C2(new_n228), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT67), .B1(new_n231), .B2(new_n253), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT66), .B1(new_n236), .B2(new_n212), .ZN(new_n257));
  INV_X1    g071(.A(new_n216), .ZN(new_n258));
  OAI22_X1  g072(.A1(new_n255), .A2(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n203), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(KEYINPUT10), .A3(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n224), .A2(new_n240), .A3(new_n252), .A4(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G110), .B(G140), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n264), .A2(G227), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n263), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n224), .A2(new_n240), .A3(new_n261), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G137), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(G137), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(KEYINPUT11), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT65), .A2(G137), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT65), .A2(G137), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT11), .A2(G134), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G131), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n244), .A2(new_n248), .A3(new_n249), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n222), .B1(new_n257), .B2(new_n258), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n260), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n205), .A2(new_n207), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n228), .B1(new_n287), .B2(new_n209), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n211), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n254), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n217), .A3(new_n203), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n293), .A2(KEYINPUT82), .A3(KEYINPUT12), .A4(new_n280), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n252), .B1(new_n285), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(KEYINPUT12), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT82), .B1(new_n295), .B2(KEYINPUT12), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n262), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(KEYINPUT12), .A3(new_n280), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT12), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n290), .A2(new_n254), .B1(new_n215), .B2(new_n216), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n223), .B1(new_n305), .B2(new_n203), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n306), .B2(new_n252), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n307), .A3(new_n294), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT83), .A3(new_n262), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n266), .B(KEYINPUT80), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n283), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G469), .B1(new_n312), .B2(G902), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n267), .B1(new_n281), .B2(new_n262), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n303), .A2(KEYINPUT84), .A3(new_n307), .A4(new_n294), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n268), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n315), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G469), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n189), .B1(new_n313), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n325));
  OR2_X1    g139(.A1(KEYINPUT68), .A2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT68), .A2(G119), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(G116), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G116), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G119), .ZN(new_n330));
  INV_X1    g144(.A(G113), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT2), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G113), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n328), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n328), .B2(new_n330), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n325), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n328), .A2(new_n330), .ZN(new_n339));
  INV_X1    g153(.A(new_n335), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n328), .A2(new_n330), .A3(new_n335), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT69), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n227), .A2(new_n338), .A3(new_n343), .A4(new_n239), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n326), .A2(new_n345), .A3(G116), .A4(new_n327), .ZN(new_n346));
  OAI211_X1 g160(.A(G113), .B(new_n346), .C1(new_n339), .C2(new_n345), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n260), .A2(new_n347), .A3(new_n342), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G122), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n344), .A2(new_n348), .A3(new_n350), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(KEYINPUT6), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n291), .A2(new_n355), .A3(new_n217), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n208), .A2(new_n210), .A3(new_n232), .ZN(new_n357));
  INV_X1    g171(.A(new_n234), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n288), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G125), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G224), .A3(new_n264), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n264), .A2(G224), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n356), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n349), .A2(new_n366), .A3(new_n351), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n354), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n356), .A2(KEYINPUT7), .A3(new_n360), .A4(new_n363), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n350), .B(KEYINPUT8), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n328), .A2(KEYINPUT5), .A3(new_n330), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n346), .A2(G113), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n342), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(new_n203), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n347), .A2(new_n342), .B1(new_n199), .B2(new_n202), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n369), .A2(new_n353), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n360), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(new_n356), .B2(KEYINPUT85), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n305), .A2(new_n380), .A3(new_n355), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n379), .A2(new_n381), .B1(KEYINPUT7), .B2(new_n363), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n377), .B1(new_n382), .B2(KEYINPUT86), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n356), .A2(KEYINPUT85), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n360), .A3(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n363), .A2(KEYINPUT7), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n385), .A2(KEYINPUT86), .A3(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n322), .B(new_n368), .C1(new_n383), .C2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G210), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n386), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n382), .A2(KEYINPUT86), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n377), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(new_n322), .A3(new_n389), .A4(new_n368), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G214), .B1(G237), .B2(G902), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT87), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n401));
  INV_X1    g215(.A(new_n399), .ZN(new_n402));
  AOI211_X1 g216(.A(new_n401), .B(new_n402), .C1(new_n391), .C2(new_n397), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT96), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n187), .A2(new_n405), .A3(G953), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT13), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT93), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT93), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT13), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n409), .A2(new_n411), .B1(new_n211), .B2(G143), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT94), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT95), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT95), .B1(new_n418), .B2(new_n414), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT94), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n204), .A2(G128), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n418), .B(new_n420), .C1(new_n414), .C2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n413), .A2(new_n417), .A3(new_n419), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G134), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n329), .A2(G122), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n329), .A2(G122), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n191), .ZN(new_n428));
  INV_X1    g242(.A(new_n421), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n418), .A2(new_n270), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(new_n426), .A3(G107), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G134), .B1(new_n407), .B2(new_n421), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n430), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n191), .B1(new_n425), .B2(KEYINPUT14), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n437), .A2(new_n427), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n427), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n406), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n432), .B1(new_n423), .B2(G134), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n443));
  INV_X1    g257(.A(new_n406), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n404), .B(new_n322), .C1(new_n441), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G478), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n434), .A2(new_n440), .A3(new_n406), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n444), .B1(new_n442), .B2(new_n443), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n448), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n404), .A3(new_n322), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(G234), .A2(G237), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n455), .A2(G952), .A3(new_n264), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(G898), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT97), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n455), .A2(G902), .A3(G953), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n449), .A2(new_n454), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT19), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n355), .A2(G140), .ZN(new_n466));
  INV_X1    g280(.A(G140), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G125), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(G125), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n355), .A2(G140), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT19), .ZN(new_n472));
  AOI21_X1  g286(.A(G146), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT16), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT16), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n466), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n474), .A2(G146), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n464), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G237), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(new_n264), .A3(G143), .A4(G214), .ZN(new_n480));
  INV_X1    g294(.A(G214), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n481), .A2(G237), .A3(G953), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n287), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G131), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n249), .B(new_n480), .C1(new_n287), .C2(new_n482), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT19), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT19), .B1(new_n470), .B2(new_n471), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n209), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n474), .A2(new_n476), .A3(G146), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(KEYINPUT90), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n478), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n493));
  OAI211_X1 g307(.A(KEYINPUT18), .B(G131), .C1(new_n483), .C2(new_n493), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n287), .A2(new_n482), .ZN(new_n495));
  NAND2_X1  g309(.A1(KEYINPUT18), .A2(G131), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(KEYINPUT89), .A3(new_n496), .A4(new_n480), .ZN(new_n497));
  OAI21_X1  g311(.A(G146), .B1(new_n466), .B2(new_n468), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n470), .A2(new_n471), .A3(new_n209), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n498), .B2(new_n499), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n494), .B(new_n497), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n492), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n200), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n483), .A2(KEYINPUT17), .A3(G131), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n484), .A2(new_n510), .A3(new_n485), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n514));
  AOI21_X1  g328(.A(G146), .B1(new_n474), .B2(new_n476), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n477), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n474), .A2(new_n476), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n209), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT91), .A3(new_n490), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n483), .A2(new_n512), .A3(KEYINPUT17), .A4(G131), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n506), .B(new_n503), .C1(new_n513), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n508), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(G475), .A2(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT20), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n503), .B1(new_n513), .B2(new_n521), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n507), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n522), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n322), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n526), .A2(new_n528), .B1(new_n532), .B2(G475), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n463), .A2(new_n533), .A3(KEYINPUT98), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n527), .B1(new_n523), .B2(new_n524), .ZN(new_n536));
  INV_X1    g350(.A(new_n524), .ZN(new_n537));
  AOI211_X1 g351(.A(KEYINPUT20), .B(new_n537), .C1(new_n508), .C2(new_n522), .ZN(new_n538));
  INV_X1    g352(.A(G475), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n530), .B2(new_n522), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n536), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n449), .A2(new_n454), .A3(new_n462), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n400), .A2(new_n403), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT22), .B(G137), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n490), .A2(new_n499), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n326), .A2(new_n327), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n211), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n552), .A2(KEYINPUT77), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n326), .A2(G128), .A3(new_n327), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n552), .A2(KEYINPUT77), .B1(KEYINPUT23), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G110), .ZN(new_n557));
  INV_X1    g371(.A(G119), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G128), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT23), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n554), .B1(new_n558), .B2(G128), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT24), .B(G110), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n550), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n562), .A2(new_n563), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n518), .A2(new_n490), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n556), .A2(new_n560), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n568), .B1(new_n569), .B2(G110), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n549), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n553), .A2(new_n555), .B1(KEYINPUT23), .B2(new_n559), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n566), .B(new_n567), .C1(new_n572), .C2(new_n557), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n572), .A2(new_n557), .B1(new_n562), .B2(new_n563), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n573), .B(new_n548), .C1(new_n574), .C2(new_n550), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(new_n575), .A3(new_n322), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT25), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n405), .B1(G234), .B2(new_n322), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n575), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT78), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n338), .A2(new_n343), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n237), .A2(new_n280), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n245), .A2(new_n246), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n271), .B1(new_n590), .B2(new_n270), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n279), .B1(new_n591), .B2(new_n249), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n305), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n588), .B1(new_n593), .B2(KEYINPUT74), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(new_n589), .C1(new_n305), .C2(new_n592), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT28), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT71), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n305), .B2(new_n592), .ZN(new_n599));
  INV_X1    g413(.A(new_n592), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n259), .A2(KEYINPUT71), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n589), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n237), .A2(new_n280), .A3(KEYINPUT70), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n588), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n252), .A2(new_n359), .A3(new_n603), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT70), .B1(new_n237), .B2(new_n280), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(new_n599), .A3(new_n601), .A4(new_n587), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n597), .B1(new_n612), .B2(KEYINPUT28), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT26), .B(G101), .ZN(new_n614));
  INV_X1    g428(.A(G210), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n615), .A2(G237), .A3(G953), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT29), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(G902), .B1(new_n613), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n619), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n610), .A2(KEYINPUT30), .A3(new_n599), .A4(new_n601), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT30), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n587), .B1(new_n593), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT72), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n624), .A2(KEYINPUT72), .A3(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n623), .B1(new_n631), .B2(new_n611), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n593), .A2(new_n588), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n604), .A2(new_n605), .A3(new_n587), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n633), .B1(new_n602), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT28), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n593), .A2(KEYINPUT74), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n596), .A3(new_n587), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT28), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n636), .A2(new_n623), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n620), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n622), .B1(new_n632), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(G472), .ZN(new_n644));
  NOR2_X1   g458(.A1(G472), .A2(G902), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT75), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n639), .B1(new_n611), .B2(new_n633), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n646), .B(new_n619), .C1(new_n647), .C2(new_n597), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n611), .A2(new_n623), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n629), .B2(new_n630), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT31), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n649), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n624), .A2(KEYINPUT72), .A3(new_n626), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT72), .B1(new_n624), .B2(new_n626), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n651), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n623), .B1(new_n636), .B2(new_n640), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(new_n646), .ZN(new_n658));
  OAI211_X1 g472(.A(KEYINPUT32), .B(new_n645), .C1(new_n652), .C2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n645), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n661));
  AOI22_X1  g475(.A1(KEYINPUT31), .A2(new_n661), .B1(new_n657), .B2(new_n646), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n619), .B1(new_n647), .B2(new_n597), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n650), .A2(new_n651), .B1(new_n663), .B2(KEYINPUT75), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT76), .B(KEYINPUT32), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n644), .B(new_n659), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n324), .A2(new_n545), .A3(new_n586), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G101), .ZN(G3));
  AND3_X1   g483(.A1(new_n308), .A2(KEYINPUT83), .A3(new_n262), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT83), .B1(new_n308), .B2(new_n262), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n311), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(G469), .A3(new_n282), .ZN(new_n673));
  NAND2_X1  g487(.A1(G469), .A2(G902), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n323), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n189), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n661), .A2(KEYINPUT31), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n663), .A2(KEYINPUT75), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n648), .A3(new_n679), .A4(new_n656), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n645), .ZN(new_n681));
  AOI21_X1  g495(.A(G902), .B1(new_n662), .B2(new_n664), .ZN(new_n682));
  INV_X1    g496(.A(G472), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n586), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n398), .A2(new_n399), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n461), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n536), .A2(new_n538), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n540), .A2(new_n539), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n447), .A2(G902), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT33), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT99), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n692), .A2(KEYINPUT99), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n693), .B(new_n694), .C1(new_n441), .C2(new_n445), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT99), .A4(new_n692), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(G478), .B1(new_n452), .B2(new_n322), .ZN(new_n698));
  OAI22_X1  g512(.A1(new_n688), .A2(new_n689), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT100), .Z(new_n700));
  AND2_X1   g514(.A1(new_n687), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n685), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT34), .B(G104), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G6));
  NAND2_X1  g518(.A1(new_n689), .A2(KEYINPUT101), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n449), .A2(new_n454), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n540), .B2(new_n539), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n686), .A2(new_n688), .A3(new_n461), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n685), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT102), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT103), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT35), .B(G107), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G9));
  AOI21_X1  g529(.A(new_n683), .B1(new_n680), .B2(new_n322), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n565), .A2(new_n570), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n549), .A2(KEYINPUT36), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n717), .B(new_n718), .Z(new_n719));
  AOI22_X1  g533(.A1(new_n578), .A2(new_n579), .B1(new_n719), .B2(new_n583), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n716), .A2(new_n665), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n324), .A2(new_n545), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT37), .B(G110), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G12));
  INV_X1    g538(.A(new_n720), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n402), .B1(new_n391), .B2(new_n397), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n526), .A2(new_n528), .ZN(new_n727));
  INV_X1    g541(.A(new_n456), .ZN(new_n728));
  INV_X1    g542(.A(new_n460), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT104), .B(G900), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n709), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n725), .A2(new_n726), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n667), .A2(new_n676), .A3(new_n675), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G128), .ZN(G30));
  XNOR2_X1  g550(.A(new_n731), .B(KEYINPUT39), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n324), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n740));
  INV_X1    g554(.A(new_n666), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n681), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n612), .A2(new_n619), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n661), .A2(KEYINPUT106), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n322), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT106), .B1(new_n661), .B2(new_n743), .ZN(new_n746));
  OAI21_X1  g560(.A(G472), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n742), .A2(new_n659), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n398), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n541), .A2(new_n706), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n399), .A2(new_n750), .A3(new_n720), .A4(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n739), .A2(new_n740), .A3(new_n748), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n287), .ZN(G45));
  AOI22_X1  g569(.A1(new_n665), .A2(KEYINPUT32), .B1(G472), .B2(new_n643), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n720), .B1(new_n756), .B2(new_n742), .ZN(new_n757));
  INV_X1    g571(.A(new_n699), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n758), .A2(new_n731), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT107), .A3(new_n726), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n731), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n761), .B1(new_n686), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n757), .A2(new_n324), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G146), .ZN(G48));
  AOI21_X1  g580(.A(new_n585), .B1(new_n756), .B2(new_n742), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n318), .A2(new_n268), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n308), .A2(new_n316), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n314), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n771), .B2(G902), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT108), .A3(new_n323), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(G469), .C1(new_n771), .C2(G902), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n189), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n701), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT41), .B(G113), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT109), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n779), .B(new_n781), .ZN(G15));
  NAND2_X1  g596(.A1(new_n778), .A2(new_n710), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G116), .ZN(G18));
  INV_X1    g598(.A(new_n544), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n757), .A2(new_n726), .A3(new_n785), .A4(new_n776), .ZN(new_n786));
  XNOR2_X1  g600(.A(KEYINPUT110), .B(G119), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(G21));
  AOI21_X1  g602(.A(new_n639), .B1(new_n607), .B2(new_n611), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n619), .B1(new_n789), .B2(new_n597), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n678), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n790), .B(KEYINPUT112), .C1(new_n650), .C2(new_n651), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n656), .A3(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n645), .B(KEYINPUT111), .Z(new_n796));
  AOI21_X1  g610(.A(new_n716), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n726), .A2(new_n462), .A3(new_n752), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n776), .A2(new_n586), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G122), .ZN(G24));
  NAND2_X1  g614(.A1(new_n794), .A2(new_n656), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT112), .B1(new_n678), .B2(new_n790), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n680), .A2(new_n322), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(G472), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n803), .A2(new_n805), .A3(new_n725), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n776), .A3(new_n726), .A4(new_n759), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G125), .ZN(G27));
  NAND2_X1  g622(.A1(new_n644), .A2(new_n659), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT32), .B1(new_n680), .B2(new_n645), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n586), .B(new_n759), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n391), .A2(new_n399), .A3(new_n397), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n675), .A2(new_n676), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT42), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n675), .A2(new_n676), .A3(new_n813), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n762), .A2(KEYINPUT42), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n767), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(new_n249), .ZN(G33));
  NAND3_X1  g634(.A1(new_n767), .A2(new_n733), .A3(new_n816), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G134), .ZN(G36));
  OR2_X1    g636(.A1(new_n312), .A2(KEYINPUT45), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n312), .A2(KEYINPUT45), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(G469), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n674), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT46), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(KEYINPUT46), .A3(new_n674), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n828), .A2(KEYINPUT114), .B1(KEYINPUT113), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n831), .A3(new_n827), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n323), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n697), .A2(new_n698), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n533), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT43), .Z(new_n837));
  OAI211_X1 g651(.A(new_n837), .B(new_n725), .C1(new_n665), .C2(new_n716), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT44), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n812), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n834), .A2(new_n676), .A3(new_n737), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G137), .ZN(G39));
  NAND2_X1  g658(.A1(new_n834), .A2(new_n676), .ZN(new_n845));
  XNOR2_X1  g659(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n834), .A2(new_n676), .A3(new_n848), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n667), .A2(new_n586), .A3(new_n762), .A4(new_n812), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G140), .ZN(G42));
  NAND2_X1  g666(.A1(new_n773), .A2(new_n775), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT49), .Z(new_n854));
  OR2_X1    g668(.A1(new_n748), .A2(new_n585), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n835), .A2(new_n676), .A3(new_n399), .A4(new_n533), .ZN(new_n856));
  OR4_X1    g670(.A1(new_n750), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n777), .A2(new_n812), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n837), .A2(new_n456), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n806), .A3(new_n859), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n855), .A2(new_n777), .A3(new_n728), .A4(new_n812), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n835), .A2(new_n541), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n864));
  OR3_X1    g678(.A1(new_n777), .A2(new_n399), .A3(new_n750), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n797), .A2(new_n586), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n859), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n864), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n860), .B(new_n863), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n847), .A2(new_n849), .B1(new_n189), .B2(new_n853), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n866), .A2(new_n813), .A3(new_n859), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n586), .B1(new_n809), .B2(new_n810), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n858), .A2(new_n877), .A3(new_n859), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT48), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n776), .A2(new_n726), .ZN(new_n880));
  OAI211_X1 g694(.A(G952), .B(new_n264), .C1(new_n867), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n861), .B2(new_n700), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n874), .A2(new_n875), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n720), .A2(new_n676), .A3(new_n731), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n889), .A2(new_n686), .A3(new_n751), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n748), .A2(new_n675), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n667), .A2(new_n676), .A3(new_n675), .A4(new_n725), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n760), .A2(new_n763), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n891), .B(new_n735), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n803), .A2(new_n805), .A3(new_n725), .A4(new_n759), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n880), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n888), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(KEYINPUT117), .B(new_n888), .C1(new_n894), .C2(new_n896), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n807), .A2(new_n765), .A3(new_n735), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n891), .A2(KEYINPUT52), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n895), .A2(new_n814), .ZN(new_n905));
  INV_X1    g719(.A(new_n892), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n705), .A2(new_n708), .ZN(new_n907));
  NOR4_X1   g721(.A1(new_n812), .A2(new_n706), .A3(new_n907), .A4(new_n732), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n815), .A3(new_n818), .A4(new_n821), .ZN(new_n910));
  AND4_X1   g724(.A1(new_n586), .A2(new_n798), .A3(new_n803), .A4(new_n805), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n532), .A2(G475), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n706), .A2(new_n727), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n699), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT116), .B1(new_n835), .B2(new_n541), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n462), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n917), .A2(new_n400), .A3(new_n403), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n776), .A2(new_n911), .B1(new_n685), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n324), .B(new_n545), .C1(new_n767), .C2(new_n721), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n767), .B(new_n776), .C1(new_n701), .C2(new_n710), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n919), .A2(new_n786), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n910), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n904), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT53), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n891), .A2(new_n735), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n927), .A2(KEYINPUT52), .A3(new_n765), .A4(new_n807), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n897), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n923), .A2(KEYINPUT53), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n887), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n910), .A2(new_n922), .A3(new_n925), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n921), .A2(new_n786), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n716), .A2(new_n585), .A3(new_n665), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n918), .A2(new_n324), .A3(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n799), .A2(new_n668), .A3(new_n935), .A4(new_n722), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n806), .A2(new_n816), .A3(new_n759), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n324), .A2(new_n667), .A3(new_n725), .A4(new_n908), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n821), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n819), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n929), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  AOI22_X1  g756(.A1(new_n904), .A2(new_n932), .B1(new_n942), .B2(new_n925), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n931), .B1(new_n887), .B2(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n871), .B(KEYINPUT51), .C1(new_n872), .C2(new_n873), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n886), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(G952), .A2(G953), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n857), .B1(new_n946), .B2(new_n947), .ZN(G75));
  NOR2_X1   g762(.A1(new_n264), .A2(G952), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n943), .B2(new_n322), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n937), .A2(new_n941), .A3(KEYINPUT53), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n897), .A2(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n900), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT53), .B1(new_n923), .B2(new_n929), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT121), .B(G902), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n952), .A2(new_n957), .A3(new_n390), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n354), .A2(new_n367), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(new_n365), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT55), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n961), .A2(KEYINPUT56), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n950), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n943), .A2(new_n615), .A3(new_n322), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n964), .B2(KEYINPUT56), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT120), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(G51));
  INV_X1    g783(.A(new_n825), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n952), .A2(new_n957), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT54), .B1(new_n955), .B2(new_n956), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n904), .A2(new_n932), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n942), .A2(new_n925), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n974), .A3(new_n887), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n674), .B(KEYINPUT57), .Z(new_n977));
  AOI21_X1  g791(.A(new_n771), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n950), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT122), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT122), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n950), .C1(new_n971), .C2(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G54));
  NAND4_X1  g797(.A1(new_n952), .A2(new_n957), .A3(KEYINPUT58), .A4(G475), .ZN(new_n984));
  INV_X1    g798(.A(new_n523), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n986), .A2(new_n987), .A3(new_n949), .ZN(G60));
  NAND2_X1  g802(.A1(new_n695), .A2(new_n696), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(G478), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT59), .Z(new_n992));
  NOR2_X1   g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n949), .B1(new_n976), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(KEYINPUT123), .ZN(new_n995));
  INV_X1    g809(.A(new_n976), .ZN(new_n996));
  INV_X1    g810(.A(new_n993), .ZN(new_n997));
  OAI211_X1 g811(.A(KEYINPUT123), .B(new_n950), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n990), .B1(new_n944), .B2(new_n992), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(G63));
  NAND2_X1  g814(.A1(G217), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT124), .Z(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT60), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n943), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n719), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1005), .B(new_n950), .C1(new_n582), .C2(new_n1004), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G66));
  INV_X1    g822(.A(G224), .ZN(new_n1009));
  OAI21_X1  g823(.A(G953), .B1(new_n459), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n922), .B(KEYINPUT125), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(G953), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT126), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n959), .B1(G898), .B2(new_n264), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(G69));
  NAND2_X1  g829(.A1(new_n593), .A2(new_n625), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n624), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n469), .A2(new_n472), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n813), .B1(new_n915), .B2(new_n916), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n768), .A2(new_n738), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n754), .A2(new_n901), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT62), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n754), .A2(KEYINPUT62), .A3(new_n901), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n851), .A2(new_n843), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1020), .B1(new_n1028), .B2(new_n264), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n264), .B1(G227), .B2(G900), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n877), .A2(new_n726), .A3(new_n752), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n834), .A2(new_n676), .A3(new_n737), .A4(new_n1036), .ZN(new_n1037));
  AND4_X1   g851(.A1(new_n815), .A2(new_n901), .A3(new_n818), .A4(new_n821), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n843), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1039), .A2(new_n851), .A3(new_n264), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1019), .B1(G900), .B2(G953), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1042), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1044));
  AOI211_X1 g858(.A(KEYINPUT127), .B(new_n1020), .C1(new_n1028), .C2(new_n264), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1032), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1043), .A2(new_n1046), .ZN(G72));
  NAND2_X1  g861(.A1(new_n631), .A2(new_n611), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1039), .A2(new_n851), .A3(new_n1011), .ZN(new_n1049));
  NAND2_X1  g863(.A1(G472), .A2(G902), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1050), .B(KEYINPUT63), .Z(new_n1051));
  AOI211_X1 g865(.A(new_n623), .B(new_n1048), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1048), .A2(new_n623), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n851), .A2(new_n843), .A3(new_n1011), .A4(new_n1027), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1053), .B1(new_n1054), .B2(new_n1051), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1051), .B1(new_n632), .B2(new_n650), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1056), .B1(new_n926), .B2(new_n930), .ZN(new_n1057));
  NOR4_X1   g871(.A1(new_n1052), .A2(new_n1055), .A3(new_n949), .A4(new_n1057), .ZN(G57));
endmodule


