//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n209), .A2(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n205), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n214), .B(new_n215), .C1(new_n211), .C2(new_n213), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n205), .A2(KEYINPUT88), .A3(new_n211), .A4(new_n213), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G1gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  INV_X1    g021(.A(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT16), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n221), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n221), .B2(new_n225), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT90), .B1(new_n218), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT89), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n205), .A2(new_n211), .A3(new_n213), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n215), .B1(new_n211), .B2(new_n213), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n230), .B(new_n217), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n216), .A2(new_n230), .A3(KEYINPUT17), .A4(new_n217), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n229), .B1(new_n237), .B2(new_n228), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n226), .A2(new_n227), .ZN(new_n239));
  AOI211_X1 g038(.A(KEYINPUT90), .B(new_n239), .C1(new_n235), .C2(new_n236), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n202), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n218), .B(new_n228), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n202), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT18), .B(new_n202), .C1(new_n238), .C2(new_n240), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G169gat), .B(G197gat), .Z(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n243), .A2(new_n246), .A3(new_n247), .A4(new_n254), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT34), .ZN(new_n260));
  NAND2_X1  g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n261), .B(KEYINPUT64), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G113gat), .ZN(new_n266));
  INV_X1    g065(.A(G113gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G120gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT1), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n264), .B1(new_n269), .B2(KEYINPUT67), .ZN(new_n270));
  INV_X1    g069(.A(G134gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G127gat), .ZN(new_n272));
  INV_X1    g071(.A(G127gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G134gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  XNOR2_X1  g075(.A(G113gat), .B(G120gat), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n275), .B(new_n276), .C1(new_n277), .C2(KEYINPUT1), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n270), .A2(KEYINPUT68), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n266), .A2(new_n268), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n270), .A2(new_n278), .B1(KEYINPUT68), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n280), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n278), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT69), .B1(new_n289), .B2(new_n279), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT23), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(KEYINPUT66), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT23), .B1(new_n291), .B2(new_n292), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n295), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT66), .B1(new_n293), .B2(new_n294), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT25), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n292), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT26), .ZN(new_n308));
  OR3_X1    g107(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n294), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT27), .B(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT28), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n315));
  OAI211_X1 g114(.A(KEYINPUT28), .B(new_n312), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n310), .B(new_n296), .C1(new_n313), .C2(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n302), .B1(new_n321), .B2(new_n299), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT23), .B(new_n292), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n322), .A2(new_n323), .A3(new_n294), .A4(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n318), .A3(new_n327), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n286), .A2(new_n290), .A3(new_n328), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n306), .A2(new_n318), .A3(new_n327), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n285), .B1(new_n280), .B2(new_n284), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n289), .A2(KEYINPUT69), .A3(new_n279), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n260), .B(new_n263), .C1(new_n329), .C2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n263), .B1(new_n329), .B2(new_n333), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT34), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n328), .B1(new_n286), .B2(new_n290), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n331), .A2(new_n330), .A3(new_n332), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n262), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(KEYINPUT71), .A3(new_n260), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n336), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n262), .A3(new_n340), .ZN(new_n344));
  XNOR2_X1  g143(.A(G15gat), .B(G43gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G71gat), .B(G99gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT33), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(KEYINPUT32), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT32), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT33), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n350), .B1(new_n353), .B2(new_n347), .ZN(new_n354));
  INV_X1    g153(.A(new_n347), .ZN(new_n355));
  AOI211_X1 g154(.A(KEYINPUT70), .B(new_n355), .C1(new_n344), .C2(new_n352), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n343), .B(new_n349), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(G211gat), .A2(G218gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G197gat), .A2(G204gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G197gat), .A2(G204gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G197gat), .B(G204gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n364), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G141gat), .B(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT2), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G155gat), .ZN(new_n375));
  INV_X1    g174(.A(G162gat), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT2), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n378));
  INV_X1    g177(.A(G141gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(G148gat), .ZN(new_n380));
  INV_X1    g179(.A(G148gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(G141gat), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n377), .B(new_n378), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G155gat), .B(G162gat), .Z(new_n384));
  OAI21_X1  g183(.A(KEYINPUT75), .B1(new_n380), .B2(new_n382), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n374), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n384), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n377), .B1(new_n380), .B2(new_n382), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(new_n378), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT3), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n371), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n371), .B2(KEYINPUT29), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n381), .A2(G141gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n379), .A2(G148gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n373), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n385), .A2(new_n394), .A3(new_n384), .A4(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n383), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n389), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n391), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT82), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n365), .B2(KEYINPUT82), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n392), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n401), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n404), .B1(new_n391), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(G22gat), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n405), .A2(new_n411), .A3(G22gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G50gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT84), .B(G22gat), .C1(new_n405), .C2(new_n411), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n415), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G22gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n391), .A2(new_n410), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n403), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n391), .A2(new_n402), .A3(new_n404), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n419), .B1(new_n413), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT83), .B(new_n419), .C1(new_n413), .C2(new_n427), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n422), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n349), .B1(new_n354), .B2(new_n356), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n336), .A2(new_n338), .A3(new_n342), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n357), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437));
  INV_X1    g236(.A(G85gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT0), .B(G57gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n289), .A2(new_n400), .A3(new_n279), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n400), .B1(new_n289), .B2(new_n279), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT5), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n289), .A2(new_n400), .A3(new_n279), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n448), .A2(KEYINPUT4), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n401), .B1(new_n331), .B2(new_n332), .ZN(new_n450));
  XOR2_X1   g249(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n449), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n289), .A2(new_n279), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n400), .A2(new_n392), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n386), .A2(KEYINPUT3), .A3(new_n389), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n442), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n447), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n461), .A3(new_n442), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n400), .B(new_n452), .C1(new_n286), .C2(new_n290), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT4), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n441), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(new_n401), .B(new_n451), .C1(new_n331), .C2(new_n332), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n448), .A2(KEYINPUT4), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n459), .B(new_n461), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n441), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n400), .B1(new_n286), .B2(new_n290), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n451), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n458), .B1(new_n472), .B2(new_n449), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n469), .B(new_n470), .C1(new_n473), .C2(new_n447), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n466), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n466), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n475), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT80), .B1(new_n466), .B2(new_n476), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n466), .A2(new_n474), .A3(KEYINPUT79), .A4(new_n476), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n479), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G8gat), .B(G36gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G64gat), .B(G92gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G226gat), .A2(G233gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n330), .B2(KEYINPUT29), .ZN(new_n491));
  INV_X1    g290(.A(new_n490), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n328), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n370), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n328), .A2(new_n492), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n328), .B2(new_n407), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n371), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n489), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n494), .A2(new_n497), .A3(new_n489), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT73), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT30), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT74), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT73), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n498), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT30), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n436), .A2(new_n485), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n482), .A2(new_n483), .A3(new_n477), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n436), .A2(new_n511), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n485), .A2(new_n508), .ZN(new_n515));
  INV_X1    g314(.A(new_n432), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT39), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT85), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n457), .B1(new_n467), .B2(new_n468), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(new_n443), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n463), .B2(new_n464), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n523), .A2(KEYINPUT85), .A3(new_n442), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n518), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n519), .A3(new_n443), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT85), .B1(new_n523), .B2(new_n442), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n444), .A2(new_n445), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n518), .B1(new_n528), .B2(new_n442), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n470), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT40), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n480), .B1(new_n506), .B2(new_n507), .ZN(new_n535));
  INV_X1    g334(.A(new_n533), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n525), .A2(new_n470), .A3(new_n536), .A4(new_n530), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n494), .A2(new_n497), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT37), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n494), .A2(new_n497), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n488), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT38), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT38), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n540), .A2(new_n545), .A3(new_n488), .A4(new_n542), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n544), .A2(new_n499), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n547), .A2(new_n482), .A3(new_n483), .A4(new_n477), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n538), .A2(new_n432), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n435), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n433), .A2(new_n434), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552));
  OAI22_X1  g351(.A1(new_n550), .A2(new_n551), .B1(KEYINPUT72), .B2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n554));
  NAND3_X1  g353(.A1(new_n357), .A2(new_n435), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n517), .A2(new_n549), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n259), .B1(new_n514), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT91), .ZN(new_n566));
  XOR2_X1   g365(.A(G71gat), .B(G78gat), .Z(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(KEYINPUT91), .B2(new_n565), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n569), .A2(new_n562), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n568), .A2(new_n570), .B1(new_n571), .B2(new_n567), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n239), .B1(KEYINPUT21), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n568), .A2(new_n570), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n567), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n575), .A2(new_n580), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n561), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n575), .A2(new_n580), .ZN(new_n584));
  INV_X1    g383(.A(new_n561), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n575), .A2(new_n580), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n583), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n583), .B2(new_n587), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(KEYINPUT7), .C1(G85gat), .C2(G92gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n595), .B1(new_n438), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G99gat), .ZN(new_n598));
  INV_X1    g397(.A(G106gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT95), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT95), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(G99gat), .A3(G106gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(KEYINPUT8), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n594), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n597), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G99gat), .B(G106gat), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n608), .A2(new_n603), .A3(new_n597), .A4(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n237), .A2(new_n610), .B1(KEYINPUT41), .B2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n218), .A2(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT96), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n617), .A3(new_n613), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n616), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n612), .A2(new_n617), .A3(new_n620), .A4(new_n613), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n611), .A2(KEYINPUT41), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT93), .ZN(new_n623));
  XOR2_X1   g422(.A(G134gat), .B(G162gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n619), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n619), .A2(new_n621), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n626), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n628), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n610), .A2(new_n578), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT10), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n610), .A2(new_n578), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n572), .A2(new_n609), .A3(new_n607), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n635), .B(new_n636), .C1(new_n639), .C2(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(KEYINPUT98), .A3(KEYINPUT10), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n593), .A2(new_n633), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n558), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n485), .B(KEYINPUT99), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  INV_X1    g459(.A(new_n508), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT16), .B(G8gat), .ZN(new_n664));
  OR3_X1    g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(G8gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n663), .B1(new_n662), .B2(new_n664), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT100), .Z(G1325gat));
  NOR2_X1   g468(.A1(new_n550), .A2(new_n551), .ZN(new_n670));
  AOI21_X1  g469(.A(G15gat), .B1(new_n656), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n556), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n672), .A2(G15gat), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n656), .B2(new_n673), .ZN(G1326gat));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n516), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n514), .A2(new_n557), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n632), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT44), .B(new_n633), .C1(new_n514), .C2(new_n557), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n258), .A2(KEYINPUT101), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n256), .A2(new_n684), .A3(new_n257), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(new_n593), .A3(new_n652), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n688), .A2(KEYINPUT102), .A3(new_n657), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT102), .B1(new_n688), .B2(new_n657), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(G29gat), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n593), .ZN(new_n692));
  AND4_X1   g491(.A1(new_n558), .A2(new_n692), .A3(new_n632), .A4(new_n653), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n207), .A3(new_n658), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n208), .A3(new_n661), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT46), .Z(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n688), .B2(new_n508), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1329gat));
  OAI21_X1  g499(.A(G43gat), .B1(new_n688), .B2(new_n556), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT47), .B1(new_n701), .B2(KEYINPUT103), .ZN(new_n702));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n693), .A2(new_n703), .A3(new_n670), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n702), .B(new_n705), .ZN(G1330gat));
  OAI21_X1  g505(.A(G50gat), .B1(new_n688), .B2(new_n432), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n432), .A2(G50gat), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT104), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g511(.A1(new_n593), .A2(new_n633), .ZN(new_n713));
  AOI211_X1 g512(.A(new_n713), .B(new_n653), .C1(new_n514), .C2(new_n557), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n686), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n658), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g517(.A(new_n508), .B(KEYINPUT105), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n719), .B(new_n715), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n720), .B(KEYINPUT106), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(G1333gat));
  NOR3_X1   g526(.A1(new_n715), .A2(new_n563), .A3(new_n556), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n716), .A2(new_n670), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n563), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1334gat));
  NOR2_X1   g531(.A1(new_n715), .A2(new_n432), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT108), .B(G78gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1335gat));
  INV_X1    g534(.A(new_n686), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n593), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n652), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n682), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740), .B2(new_n657), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n679), .A2(new_n632), .A3(new_n737), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT109), .Z(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(new_n438), .A3(new_n658), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n741), .B1(new_n746), .B2(new_n653), .ZN(G1336gat));
  OAI21_X1  g546(.A(G92gat), .B1(new_n740), .B2(new_n508), .ZN(new_n748));
  INV_X1    g547(.A(new_n719), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n744), .A2(new_n596), .A3(new_n652), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT52), .ZN(new_n752));
  OAI21_X1  g551(.A(G92gat), .B1(new_n740), .B2(new_n719), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n750), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(G1337gat));
  NAND4_X1  g555(.A1(new_n745), .A2(new_n598), .A3(new_n670), .A4(new_n652), .ZN(new_n757));
  OAI21_X1  g556(.A(G99gat), .B1(new_n740), .B2(new_n556), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1338gat));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n516), .B(new_n739), .C1(new_n680), .C2(new_n681), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n761), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT111), .B1(new_n761), .B2(G106gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n744), .A2(new_n599), .A3(new_n516), .A4(new_n652), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n761), .A2(G106gat), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT113), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n761), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(new_n765), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT53), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n769), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n771), .A2(new_n778), .ZN(G1339gat));
  NOR2_X1   g578(.A1(new_n654), .A2(new_n736), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n256), .A2(new_n684), .A3(new_n257), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n684), .B1(new_n256), .B2(new_n257), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n640), .A2(new_n642), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n644), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(KEYINPUT54), .A3(new_n643), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n640), .A2(new_n786), .A3(new_n641), .A4(new_n642), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n649), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n785), .A2(new_n788), .A3(KEYINPUT55), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n650), .A3(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n781), .A2(new_n782), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n238), .A2(new_n240), .A3(new_n202), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n244), .A2(new_n245), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n253), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n257), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n652), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n633), .B1(new_n794), .B2(new_n800), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n619), .A2(new_n621), .A3(new_n627), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n631), .B1(new_n619), .B2(new_n621), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n257), .B(new_n797), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT114), .B1(new_n804), .B2(new_n793), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n791), .A2(new_n650), .A3(new_n792), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n806), .A2(new_n807), .A3(new_n632), .A4(new_n798), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n801), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n780), .B1(new_n810), .B2(new_n692), .ZN(new_n811));
  INV_X1    g610(.A(new_n436), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n811), .A2(new_n812), .A3(new_n657), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n813), .A2(new_n267), .A3(new_n736), .A4(new_n719), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n805), .A2(new_n808), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n683), .A2(new_n806), .A3(new_n685), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n632), .B1(new_n818), .B2(new_n799), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n692), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n780), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n816), .B1(new_n822), .B2(new_n432), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT115), .B(new_n516), .C1(new_n820), .C2(new_n821), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n749), .A2(new_n657), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n825), .A2(new_n258), .A3(new_n670), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n815), .B1(new_n827), .B2(G113gat), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n811), .B2(new_n516), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n593), .B1(new_n801), .B2(new_n809), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n816), .B(new_n432), .C1(new_n830), .C2(new_n780), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n829), .A2(new_n670), .A3(new_n826), .A4(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n815), .B(G113gat), .C1(new_n832), .C2(new_n259), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n814), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT117), .B(new_n814), .C1(new_n828), .C2(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1340gat));
  OAI21_X1  g638(.A(G120gat), .B1(new_n832), .B2(new_n653), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n813), .A2(new_n265), .A3(new_n719), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n653), .B2(new_n841), .ZN(G1341gat));
  AND3_X1   g641(.A1(new_n813), .A2(new_n593), .A3(new_n719), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n593), .A2(G127gat), .ZN(new_n844));
  OAI22_X1  g643(.A1(new_n843), .A2(G127gat), .B1(new_n832), .B2(new_n844), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT118), .Z(G1342gat));
  NOR2_X1   g645(.A1(new_n633), .A2(new_n661), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n813), .A2(new_n271), .A3(new_n847), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT56), .Z(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n832), .B2(new_n633), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n799), .B1(new_n259), .B2(new_n793), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n633), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n809), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n780), .B1(new_n855), .B2(new_n692), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n432), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n749), .A2(new_n657), .A3(new_n672), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n822), .A2(new_n860), .A3(new_n516), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n258), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G141gat), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n672), .A2(new_n432), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT119), .Z(new_n865));
  AND3_X1   g664(.A1(new_n865), .A2(new_n658), .A3(new_n822), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n866), .A2(new_n379), .A3(new_n258), .A4(new_n719), .ZN(new_n867));
  XNOR2_X1  g666(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n859), .A2(new_n736), .A3(new_n861), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G141gat), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n867), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n852), .B(new_n869), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n873), .B1(new_n871), .B2(new_n867), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(G1344gat));
  AND2_X1   g677(.A1(new_n859), .A2(new_n861), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n381), .C1(new_n879), .C2(new_n652), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n654), .A2(new_n258), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n854), .B1(new_n793), .B2(new_n804), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n692), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(KEYINPUT57), .A3(new_n432), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n811), .B2(new_n432), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n652), .A4(new_n858), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n881), .B1(new_n888), .B2(G148gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n866), .A2(new_n719), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n652), .A2(new_n381), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n880), .A2(new_n889), .B1(new_n890), .B2(new_n891), .ZN(G1345gat));
  OAI21_X1  g691(.A(new_n375), .B1(new_n890), .B2(new_n692), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n879), .A2(G155gat), .A3(new_n593), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT122), .ZN(G1346gat));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n632), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n879), .A2(KEYINPUT123), .A3(new_n632), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(G162gat), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n866), .A2(new_n376), .A3(new_n847), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n811), .A2(new_n658), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT124), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(new_n436), .A3(new_n749), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n906), .B(new_n736), .C1(new_n325), .C2(new_n324), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n658), .A2(new_n508), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n825), .A2(new_n670), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n259), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(G1348gat));
  NOR3_X1   g710(.A1(new_n909), .A2(new_n292), .A3(new_n653), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n906), .A2(new_n652), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n292), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n909), .B2(new_n692), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n593), .A2(new_n311), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n905), .A2(new_n436), .A3(new_n749), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n906), .A2(new_n312), .A3(new_n632), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n909), .A2(new_n633), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(G190gat), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n921), .B(G190gat), .C1(new_n909), .C2(new_n633), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n920), .B1(new_n923), .B2(new_n925), .ZN(G1351gat));
  AND3_X1   g725(.A1(new_n905), .A2(new_n749), .A3(new_n864), .ZN(new_n927));
  INV_X1    g726(.A(G197gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(new_n736), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n886), .A2(new_n930), .A3(new_n887), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n860), .B1(new_n822), .B2(new_n516), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT125), .B1(new_n932), .B2(new_n885), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n658), .A2(new_n508), .A3(new_n672), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n934), .A2(new_n258), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n929), .B1(new_n936), .B2(new_n928), .ZN(G1352gat));
  INV_X1    g736(.A(G204gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n938), .A3(new_n652), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n652), .A3(new_n935), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G204gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n927), .A2(new_n943), .A3(new_n938), .A4(new_n652), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n940), .A2(new_n942), .A3(new_n944), .ZN(G1353gat));
  NOR2_X1   g744(.A1(new_n692), .A2(G211gat), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n905), .A2(new_n749), .A3(new_n864), .A4(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n886), .A2(new_n887), .A3(new_n593), .A4(new_n935), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g753(.A(KEYINPUT126), .B(new_n947), .C1(new_n950), .C2(new_n951), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1354gat));
  NAND4_X1  g755(.A1(new_n931), .A2(new_n933), .A3(new_n632), .A4(new_n935), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G218gat), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n633), .A2(G218gat), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n905), .A2(new_n749), .A3(new_n864), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(G1355gat));
endmodule


