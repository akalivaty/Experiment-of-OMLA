//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT65), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT66), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT67), .Z(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n209), .B1(new_n213), .B2(new_n216), .C1(new_n223), .C2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n237), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G222), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n253), .B1(new_n202), .B2(new_n251), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT69), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n257), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n266), .A2(new_n260), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n265), .B1(G226), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT70), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n270), .A2(G179), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n210), .B1(new_n206), .B2(new_n246), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n211), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n277), .A2(new_n279), .B1(new_n201), .B2(new_n211), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n272), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT72), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT72), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n284), .A2(new_n259), .A3(G13), .A4(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n272), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n211), .A2(G1), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G50), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n281), .B1(G50), .B2(new_n286), .C1(new_n288), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n271), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n270), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n292), .B(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n270), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n270), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n286), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n240), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT12), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n279), .A2(new_n238), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n275), .A2(new_n202), .B1(new_n211), .B2(G68), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n272), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT11), .ZN(new_n309));
  INV_X1    g0109(.A(new_n288), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(G68), .A3(new_n290), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(new_n312), .B(KEYINPUT76), .Z(new_n313));
  AOI21_X1  g0113(.A(new_n265), .B1(G238), .B2(new_n267), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n251), .A2(G226), .A3(new_n252), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n314), .B1(new_n266), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT13), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G169), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n321), .A2(new_n322), .B1(new_n323), .B2(new_n320), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n321), .A2(new_n322), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n313), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n320), .A2(new_n298), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(new_n312), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT74), .B1(new_n320), .B2(G200), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n320), .A2(KEYINPUT74), .A3(G200), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n286), .A2(G77), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n288), .A2(new_n202), .A3(new_n289), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G20), .A2(G77), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT15), .B(G87), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n335), .B1(new_n273), .B2(new_n279), .C1(new_n275), .C2(new_n336), .ZN(new_n337));
  AOI211_X1 g0137(.A(new_n333), .B(new_n334), .C1(new_n272), .C2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n251), .A2(G232), .A3(new_n252), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT73), .B(G107), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G238), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n339), .B1(new_n251), .B2(new_n341), .C1(new_n254), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n257), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n265), .B1(G244), .B2(new_n267), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n338), .B1(new_n294), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n345), .A3(new_n323), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(G200), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n338), .C1(new_n298), .C2(new_n346), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n302), .A2(new_n326), .A3(new_n332), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G58), .A2(G68), .ZN(new_n354));
  XOR2_X1   g0154(.A(new_n354), .B(KEYINPUT81), .Z(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G58), .B2(G68), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT77), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n248), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(G33), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT78), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n359), .A2(KEYINPUT78), .A3(G33), .A4(new_n360), .ZN(new_n364));
  NOR2_X1   g0164(.A1(KEYINPUT79), .A2(KEYINPUT7), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n363), .A2(new_n211), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n366), .A2(G68), .ZN(new_n367));
  AND2_X1   g0167(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n368), .A2(new_n369), .A3(new_n246), .ZN(new_n370));
  INV_X1    g0170(.A(new_n362), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n211), .B(new_n364), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  XOR2_X1   g0172(.A(KEYINPUT79), .B(KEYINPUT7), .Z(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT80), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  AND4_X1   g0175(.A1(KEYINPUT80), .A2(new_n374), .A3(G68), .A4(new_n366), .ZN(new_n376));
  OAI211_X1 g0176(.A(KEYINPUT16), .B(new_n357), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  INV_X1    g0178(.A(new_n357), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n246), .B1(new_n368), .B2(new_n369), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n249), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n250), .B2(new_n211), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n240), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n378), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n377), .A2(new_n386), .A3(new_n272), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n274), .A2(new_n289), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n310), .B1(new_n303), .B2(new_n274), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n363), .A2(new_n364), .ZN(new_n390));
  MUX2_X1   g0190(.A(G223), .B(G226), .S(G1698), .Z(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  XOR2_X1   g0193(.A(new_n393), .B(KEYINPUT82), .Z(new_n394));
  AOI21_X1  g0194(.A(new_n266), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n267), .A2(G232), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n262), .A2(new_n264), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(G169), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n395), .A2(new_n398), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G179), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n387), .A2(new_n389), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT18), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n298), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(G200), .B2(new_n400), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n387), .A2(new_n389), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n404), .B1(new_n407), .B2(KEYINPUT83), .ZN(new_n408));
  INV_X1    g0208(.A(new_n389), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n374), .A2(G68), .A3(new_n366), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT80), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n374), .A2(KEYINPUT80), .A3(G68), .A4(new_n366), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n379), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n287), .B1(new_n414), .B2(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n409), .B1(new_n415), .B2(new_n386), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT83), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT84), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(new_n406), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n408), .A2(new_n419), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n407), .A2(KEYINPUT84), .A3(KEYINPUT17), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n403), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n353), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n251), .A2(new_n211), .A3(G87), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT90), .B(KEYINPUT22), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n390), .A2(new_n211), .A3(G87), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(KEYINPUT22), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n211), .A2(KEYINPUT23), .A3(G107), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT91), .ZN(new_n431));
  INV_X1    g0231(.A(G116), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n246), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n211), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT23), .B1(new_n340), .B2(new_n211), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT24), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G87), .ZN(new_n438));
  AOI211_X1 g0238(.A(G20), .B(new_n438), .C1(new_n363), .C2(new_n364), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT22), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n439), .A2(new_n440), .B1(new_n426), .B2(new_n425), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT24), .ZN(new_n442));
  INV_X1    g0242(.A(new_n436), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n437), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n272), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT92), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(KEYINPUT92), .A3(new_n272), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n246), .A2(G1), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n288), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n303), .A2(KEYINPUT25), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT25), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n286), .B2(G107), .ZN(new_n456));
  AOI22_X1  g0256(.A1(G107), .A2(new_n452), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G257), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n252), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n390), .A2(new_n459), .B1(G33), .B2(G294), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT93), .ZN(new_n461));
  INV_X1    g0261(.A(G250), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1698), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n390), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n390), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n257), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT5), .B(G41), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n264), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n257), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G264), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n467), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT94), .ZN(new_n475));
  INV_X1    g0275(.A(new_n473), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n466), .B2(new_n257), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT94), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n471), .ZN(new_n479));
  AOI21_X1  g0279(.A(G190), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n474), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G200), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n450), .B(new_n457), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n470), .A2(new_n469), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(new_n266), .A3(KEYINPUT88), .A4(G270), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n471), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT88), .B1(new_n472), .B2(G270), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G264), .A2(G1698), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n390), .A2(new_n490), .B1(G303), .B2(new_n250), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(G1698), .B1(new_n363), .B2(new_n364), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT89), .B1(new_n493), .B2(G257), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(KEYINPUT89), .A3(G257), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G190), .B(new_n488), .C1(new_n497), .C2(new_n266), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n286), .A2(G116), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n452), .B2(G116), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  INV_X1    g0301(.A(G97), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n211), .C1(G33), .C2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n272), .C1(new_n211), .C2(G116), .ZN(new_n504));
  XOR2_X1   g0304(.A(new_n504), .B(KEYINPUT20), .Z(new_n505));
  NAND2_X1  g0305(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n488), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n493), .A2(KEYINPUT89), .A3(G257), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n491), .B1(new_n509), .B2(new_n494), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n510), .B2(new_n257), .ZN(new_n511));
  INV_X1    g0311(.A(G200), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n498), .B(new_n507), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n257), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n508), .A2(new_n323), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n506), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n506), .A2(G169), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT21), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n511), .A2(new_n517), .A3(KEYINPUT21), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n513), .B(new_n516), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G238), .A2(G1698), .ZN(new_n523));
  INV_X1    g0323(.A(G244), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(G1698), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n363), .B2(new_n364), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n257), .B1(new_n527), .B2(new_n433), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n264), .A2(new_n469), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n469), .A2(new_n462), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n266), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n512), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n532), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n535), .B2(G190), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n288), .A2(new_n438), .A3(new_n451), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n390), .A2(new_n211), .A3(G68), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n211), .B1(new_n317), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n438), .A2(new_n502), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n340), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n540), .B1(new_n275), .B2(new_n502), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT87), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT87), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n546), .B(new_n540), .C1(new_n275), .C2(new_n502), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n287), .B1(new_n539), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n336), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n286), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n536), .A2(new_n538), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n452), .A2(new_n550), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n535), .A2(new_n323), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n534), .A2(new_n294), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT85), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n452), .A2(new_n502), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n303), .A2(G97), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n562), .ZN(new_n564));
  OAI211_X1 g0364(.A(KEYINPUT85), .B(new_n564), .C1(new_n452), .C2(new_n502), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n453), .A2(KEYINPUT6), .A3(G97), .ZN(new_n566));
  XOR2_X1   g0366(.A(G97), .B(G107), .Z(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(KEYINPUT6), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(G20), .B1(G77), .B2(new_n278), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n384), .B2(new_n341), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n563), .A2(new_n565), .B1(new_n272), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n471), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(G257), .B2(new_n472), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n252), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n501), .A3(new_n576), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n524), .B(G1698), .C1(new_n363), .C2(new_n364), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT86), .B1(new_n578), .B2(KEYINPUT4), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n390), .A2(G244), .A3(new_n252), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT86), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT4), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n577), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n323), .B(new_n574), .C1(new_n584), .C2(new_n266), .ZN(new_n585));
  INV_X1    g0385(.A(new_n574), .ZN(new_n586));
  INV_X1    g0386(.A(new_n577), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n578), .A2(KEYINPUT86), .A3(KEYINPUT4), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n581), .B1(new_n580), .B2(new_n582), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n590), .B2(new_n257), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n572), .B(new_n585), .C1(new_n591), .C2(G169), .ZN(new_n592));
  OAI211_X1 g0392(.A(G190), .B(new_n574), .C1(new_n584), .C2(new_n266), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n571), .C1(new_n591), .C2(new_n512), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n559), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n475), .A2(G169), .A3(new_n479), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n481), .A2(G179), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT92), .B1(new_n445), .B2(new_n272), .ZN(new_n599));
  AOI211_X1 g0399(.A(new_n447), .B(new_n287), .C1(new_n437), .C2(new_n444), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n457), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n483), .A2(new_n522), .A3(new_n595), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n424), .A2(new_n603), .ZN(G372));
  INV_X1    g0404(.A(KEYINPUT26), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT95), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n552), .B2(new_n538), .ZN(new_n607));
  NOR4_X1   g0407(.A1(new_n549), .A2(KEYINPUT95), .A3(new_n537), .A4(new_n551), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n536), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n558), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n605), .B1(new_n610), .B2(new_n592), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT96), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n574), .B1(new_n584), .B2(new_n266), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n571), .B1(new_n614), .B2(new_n294), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n559), .A2(new_n615), .A3(KEYINPUT26), .A4(new_n585), .ZN(new_n616));
  OAI211_X1 g0416(.A(KEYINPUT96), .B(new_n605), .C1(new_n610), .C2(new_n592), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n592), .A2(new_n594), .A3(new_n609), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n450), .A2(new_n457), .B1(new_n596), .B2(new_n597), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n514), .A2(new_n488), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(G169), .A4(new_n506), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n518), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n516), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n483), .B(new_n620), .C1(new_n621), .C2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n618), .A2(new_n627), .A3(new_n558), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n423), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n332), .A2(new_n348), .A3(new_n347), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n630), .A2(new_n326), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n407), .A2(KEYINPUT84), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n408), .A2(new_n419), .B1(new_n632), .B2(new_n404), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n403), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n300), .A2(new_n301), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n295), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n629), .A2(new_n636), .ZN(G369));
  INV_X1    g0437(.A(G13), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n638), .A2(G1), .A3(G20), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(KEYINPUT97), .A3(KEYINPUT27), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT97), .B1(new_n640), .B2(KEYINPUT27), .ZN(new_n643));
  OAI221_X1 g0443(.A(G213), .B1(KEYINPUT27), .B2(new_n640), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n507), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n626), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n649), .B(KEYINPUT98), .C1(new_n521), .C2(new_n648), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(G330), .ZN(new_n653));
  INV_X1    g0453(.A(new_n601), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n483), .B(new_n602), .C1(new_n654), .C2(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n621), .A2(new_n646), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n621), .A2(new_n647), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n625), .A2(new_n516), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n646), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n602), .A3(new_n483), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n207), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n340), .A2(G116), .A3(new_n542), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n214), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n628), .A2(new_n647), .ZN(new_n671));
  INV_X1    g0471(.A(new_n558), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n475), .A2(new_n479), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n298), .ZN(new_n674));
  INV_X1    g0474(.A(new_n482), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n619), .B1(new_n676), .B2(new_n654), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n660), .A2(new_n602), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n672), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n559), .A2(new_n615), .A3(new_n605), .A4(new_n585), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT26), .B1(new_n610), .B2(new_n592), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n646), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  MUX2_X1   g0483(.A(new_n671), .B(new_n683), .S(KEYINPUT29), .Z(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n514), .A2(new_n477), .A3(new_n515), .A4(new_n535), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(new_n614), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n390), .A2(new_n463), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT93), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n390), .A2(new_n461), .A3(new_n463), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n266), .B1(new_n691), .B2(new_n460), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n488), .A2(G179), .A3(new_n528), .A4(new_n532), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n692), .A2(new_n693), .A3(new_n476), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n591), .A3(KEYINPUT30), .A4(new_n514), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n535), .A2(G179), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n614), .A2(new_n622), .A3(new_n474), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n687), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n646), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n699), .B(new_n702), .C1(new_n603), .C2(new_n646), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n684), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n670), .B1(new_n706), .B2(G1), .ZN(G364));
  NAND3_X1  g0507(.A1(new_n251), .A2(G355), .A3(new_n207), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n215), .A2(new_n468), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n244), .B2(new_n468), .ZN(new_n710));
  INV_X1    g0510(.A(new_n390), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n207), .ZN(new_n712));
  OAI221_X1 g0512(.A(new_n708), .B1(G116), .B2(new_n207), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n210), .B1(G20), .B2(new_n294), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n638), .A2(G20), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n259), .B1(new_n720), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n665), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n716), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n652), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n211), .A2(new_n323), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n298), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G326), .ZN(new_n731));
  INV_X1    g0531(.A(G294), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n298), .A2(G179), .A3(G200), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n211), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n730), .A2(new_n731), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n728), .A2(G190), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT33), .B(G317), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n211), .A2(G179), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(G190), .A3(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n251), .B1(new_n741), .B2(G303), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT100), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n298), .A3(G200), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT99), .Z(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G283), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n727), .A2(G190), .A3(new_n512), .ZN(new_n747));
  INV_X1    g0547(.A(G322), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G190), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n727), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G311), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n747), .A2(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n739), .A2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n752), .B1(G329), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n738), .A2(new_n743), .A3(new_n746), .A4(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n736), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n757), .A2(new_n240), .B1(new_n740), .B2(new_n438), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(G159), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n730), .A2(new_n238), .B1(new_n759), .B2(KEYINPUT32), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n745), .A2(G107), .ZN(new_n762));
  INV_X1    g0562(.A(G58), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n251), .B1(new_n747), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n750), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n764), .B1(G77), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n734), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n759), .A2(KEYINPUT32), .B1(new_n767), .B2(G97), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n761), .A2(new_n762), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n756), .A2(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n724), .B(new_n726), .C1(new_n717), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n653), .A2(new_n723), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n652), .A2(G330), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(G396));
  NOR2_X1   g0576(.A1(new_n349), .A2(new_n646), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n351), .B1(new_n338), .B2(new_n647), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n777), .B1(new_n349), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n628), .A2(new_n647), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT103), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n646), .B1(new_n679), .B2(new_n618), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(KEYINPUT103), .A3(new_n779), .ZN(new_n784));
  INV_X1    g0584(.A(new_n779), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n782), .A2(new_n784), .B1(new_n671), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n723), .B1(new_n787), .B2(new_n704), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n704), .B2(new_n787), .ZN(new_n789));
  INV_X1    g0589(.A(new_n717), .ZN(new_n790));
  INV_X1    g0590(.A(new_n745), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n438), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n250), .B1(new_n750), .B2(new_n432), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n729), .A2(G303), .B1(new_n741), .B2(G107), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n502), .B2(new_n734), .C1(new_n795), .C2(new_n757), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n747), .A2(new_n732), .B1(new_n753), .B2(new_n751), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n792), .A2(new_n793), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G137), .A2(new_n729), .B1(new_n736), .B2(G150), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT101), .Z(new_n801));
  INV_X1    g0601(.A(G143), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n802), .B2(new_n747), .C1(new_n803), .C2(new_n750), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT34), .Z(new_n805));
  NAND2_X1  g0605(.A1(new_n745), .A2(G68), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n741), .A2(G50), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n767), .A2(G58), .B1(G132), .B2(new_n754), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n806), .A2(new_n390), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n799), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT102), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n790), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  INV_X1    g0613(.A(new_n723), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n717), .A2(new_n714), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n202), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n813), .B(new_n816), .C1(new_n715), .C2(new_n779), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n789), .A2(new_n817), .ZN(G384));
  NOR2_X1   g0618(.A1(new_n720), .A2(new_n259), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n407), .A2(KEYINPUT83), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n377), .A2(new_n272), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n414), .A2(KEYINPUT16), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n389), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n401), .A2(new_n399), .A3(new_n644), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n387), .A2(new_n406), .A3(new_n417), .A4(new_n389), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n820), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT104), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT104), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n827), .A2(new_n830), .A3(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n820), .A2(new_n826), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n387), .A2(new_n389), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n401), .A2(new_n399), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n644), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n829), .A2(new_n831), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n823), .A2(new_n837), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n422), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n842), .A2(new_n844), .A3(KEYINPUT38), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT38), .B1(new_n842), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n699), .ZN(new_n848));
  AND4_X1   g0648(.A1(new_n602), .A2(new_n522), .A3(new_n483), .A4(new_n595), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n647), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n700), .A2(KEYINPUT107), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT107), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n698), .A2(new_n852), .A3(new_n646), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n701), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(KEYINPUT108), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT108), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT31), .B1(new_n700), .B2(KEYINPUT107), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n853), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n850), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT40), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n313), .A2(new_n646), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n326), .B2(new_n332), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n326), .A2(new_n332), .A3(new_n861), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n785), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n859), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n847), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n326), .A2(new_n332), .A3(new_n861), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n779), .B1(new_n868), .B2(new_n862), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n854), .A2(KEYINPUT108), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n857), .A2(new_n856), .A3(new_n853), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n869), .B1(new_n872), .B2(new_n850), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n842), .A2(new_n844), .A3(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n838), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT18), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n402), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n633), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n402), .B1(new_n416), .B2(new_n406), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n839), .B1(new_n879), .B2(new_n838), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n832), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n874), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n860), .B1(new_n873), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n867), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n423), .A2(new_n859), .ZN(new_n891));
  OAI21_X1  g0691(.A(G330), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n403), .A2(new_n837), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n868), .A2(new_n862), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n782), .A2(new_n784), .ZN(new_n897));
  INV_X1    g0697(.A(new_n777), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n847), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n895), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n326), .A2(new_n646), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n885), .B1(new_n878), .B2(new_n880), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n828), .A2(KEYINPUT104), .B1(new_n833), .B2(new_n840), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n905), .A2(new_n831), .B1(new_n422), .B2(new_n843), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n904), .B1(new_n906), .B2(KEYINPUT38), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(KEYINPUT106), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT106), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n888), .B2(KEYINPUT39), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n842), .A2(new_n844), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n908), .B1(new_n914), .B2(new_n874), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n903), .B(new_n909), .C1(new_n911), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n901), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n636), .B1(new_n684), .B2(new_n424), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n917), .B(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n819), .B1(new_n894), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n894), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n568), .A2(KEYINPUT35), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n568), .A2(KEYINPUT35), .ZN(new_n923));
  NOR4_X1   g0723(.A1(new_n922), .A2(new_n923), .A3(new_n432), .A4(new_n213), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT36), .Z(new_n925));
  INV_X1    g0725(.A(new_n214), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n355), .A2(G77), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n239), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(G1), .A3(new_n638), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n925), .A3(new_n929), .ZN(G367));
  OAI211_X1 g0730(.A(new_n592), .B(new_n594), .C1(new_n571), .C2(new_n647), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n615), .A2(new_n585), .A3(new_n646), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n662), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n592), .B1(new_n602), .B2(new_n931), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n935), .A2(KEYINPUT42), .B1(new_n647), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n607), .A2(new_n608), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n646), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(new_n558), .A3(new_n609), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n558), .B2(new_n940), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n936), .A2(new_n938), .B1(KEYINPUT43), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n658), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n933), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n945), .B(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n665), .B(KEYINPUT41), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n662), .A2(new_n659), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT44), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n933), .B1(KEYINPUT109), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT110), .Z(new_n954));
  INV_X1    g0754(.A(KEYINPUT109), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n950), .A2(new_n934), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT45), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n953), .B(KEYINPUT110), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n955), .A3(KEYINPUT44), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n957), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n946), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT111), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n662), .B1(new_n657), .B2(new_n661), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n653), .B(new_n965), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n964), .B1(new_n966), .B2(new_n705), .ZN(new_n967));
  INV_X1    g0767(.A(new_n966), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(KEYINPUT111), .A3(new_n706), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n957), .A2(new_n658), .A3(new_n961), .A4(new_n959), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n963), .A2(new_n967), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n949), .B1(new_n971), .B2(new_n706), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n948), .B1(new_n972), .B2(new_n722), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n718), .B1(new_n207), .B2(new_n336), .C1(new_n712), .C2(new_n233), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n974), .A2(new_n723), .ZN(new_n975));
  INV_X1    g0775(.A(new_n744), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n767), .A2(new_n340), .B1(new_n976), .B2(G97), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n732), .B2(new_n757), .C1(new_n751), .C2(new_n730), .ZN(new_n978));
  INV_X1    g0778(.A(new_n747), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n979), .A2(G303), .B1(new_n765), .B2(G283), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n754), .A2(G317), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n711), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n740), .A2(new_n432), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT46), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n978), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G50), .A2(new_n765), .B1(new_n754), .B2(G137), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n251), .C1(new_n277), .C2(new_n747), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n730), .A2(new_n802), .B1(new_n740), .B2(new_n763), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n757), .A2(new_n803), .B1(new_n240), .B2(new_n734), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n744), .A2(new_n202), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n975), .B1(new_n790), .B2(new_n993), .C1(new_n942), .C2(new_n725), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT112), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n973), .A2(new_n995), .ZN(G387));
  OR3_X1    g0796(.A1(new_n966), .A2(KEYINPUT113), .A3(new_n721), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT113), .B1(new_n966), .B2(new_n721), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n655), .A2(new_n656), .A3(new_n716), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n979), .A2(G317), .B1(new_n765), .B2(G303), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n751), .A2(new_n757), .B1(new_n730), .B2(new_n748), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT114), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n1002), .B2(new_n1001), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT48), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(KEYINPUT48), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n767), .A2(G283), .B1(new_n741), .B2(G294), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n744), .A2(new_n432), .B1(new_n753), .B2(new_n731), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1010), .A2(new_n390), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n747), .A2(new_n238), .B1(new_n750), .B2(new_n240), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1015), .B(new_n711), .C1(G150), .C2(new_n754), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n274), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n736), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n745), .A2(G97), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n740), .A2(new_n202), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n734), .A2(new_n336), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(G159), .C2(new_n729), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n790), .B1(new_n1014), .B2(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n230), .A2(G45), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n251), .A2(new_n207), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1025), .A2(new_n712), .B1(new_n667), .B2(new_n1026), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n273), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT50), .B1(new_n273), .B2(G50), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1028), .A2(new_n667), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(G107), .B2(new_n207), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n814), .B(new_n1024), .C1(new_n718), .C2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n997), .A2(new_n998), .B1(new_n999), .B2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n969), .A2(new_n967), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n665), .B1(new_n968), .B2(new_n706), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(G393));
  AND2_X1   g0838(.A1(new_n963), .A2(new_n970), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n722), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n718), .B1(new_n502), .B2(new_n207), .C1(new_n712), .C2(new_n237), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n723), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n792), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n750), .A2(new_n273), .B1(new_n753), .B2(new_n802), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G68), .B2(new_n741), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G77), .A2(new_n767), .B1(new_n736), .B2(G50), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1043), .A2(new_n1045), .A3(new_n390), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G150), .A2(new_n729), .B1(new_n979), .B2(G159), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G317), .A2(new_n729), .B1(new_n979), .B2(G311), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1051));
  XNOR2_X1  g0851(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n250), .B1(new_n750), .B2(new_n732), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G322), .B2(new_n754), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n736), .A2(G303), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n767), .A2(G116), .B1(new_n741), .B2(G283), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n762), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1047), .A2(new_n1049), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1042), .B1(new_n1058), .B2(new_n717), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n933), .B2(new_n725), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1039), .A2(new_n1036), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n971), .A2(new_n665), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1040), .B(new_n1060), .C1(new_n1061), .C2(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(G330), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n872), .B2(new_n850), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n423), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n636), .C1(new_n424), .C2(new_n684), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n859), .A2(G330), .A3(new_n865), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n896), .B1(new_n704), .B2(new_n785), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT103), .B1(new_n783), .B2(new_n779), .ZN(new_n1071));
  AND4_X1   g0871(.A1(KEYINPUT103), .A2(new_n628), .A3(new_n647), .A4(new_n779), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n898), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n704), .A2(new_n896), .A3(new_n785), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n627), .A2(new_n558), .A3(new_n682), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n778), .A2(new_n349), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n647), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n898), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1064), .B(new_n785), .C1(new_n872), .C2(new_n850), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n896), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1067), .B1(new_n1074), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(new_n902), .A3(new_n888), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n909), .B1(new_n911), .B2(new_n915), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n777), .B1(new_n782), .B2(new_n784), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n902), .B1(new_n1090), .B2(new_n896), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1088), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1092), .A2(new_n1068), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1075), .ZN(new_n1094));
  AND4_X1   g0894(.A1(KEYINPUT106), .A2(new_n874), .A3(new_n908), .A4(new_n887), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT106), .B1(new_n907), .B2(new_n908), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT39), .B1(new_n845), .B2(new_n846), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n903), .B1(new_n1073), .B2(new_n1082), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1087), .B(new_n1094), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1085), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1100), .B(new_n1084), .C1(new_n1092), .C2(new_n1068), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n665), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n806), .B1(new_n732), .B2(new_n753), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT116), .Z(new_n1106));
  OAI221_X1 g0906(.A(new_n250), .B1(new_n750), .B2(new_n502), .C1(new_n432), .C2(new_n747), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n734), .A2(new_n202), .B1(new_n740), .B2(new_n438), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n341), .A2(new_n757), .B1(new_n730), .B2(new_n795), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n767), .A2(G159), .B1(new_n976), .B2(G50), .ZN(new_n1111));
  INV_X1    g0911(.A(G128), .ZN(new_n1112));
  INV_X1    g0912(.A(G137), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n730), .C1(new_n1113), .C2(new_n757), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n741), .A2(G150), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  INV_X1    g0916(.A(G132), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n251), .B1(new_n747), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  INV_X1    g0919(.A(G125), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n750), .A2(new_n1119), .B1(new_n753), .B2(new_n1120), .ZN(new_n1121));
  NOR4_X1   g0921(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .A4(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n717), .B1(new_n1110), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n815), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n723), .C1(new_n1017), .C2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1089), .B2(new_n714), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1093), .A2(new_n1101), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n722), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1104), .A2(new_n1128), .ZN(G378));
  NAND2_X1  g0929(.A1(new_n292), .A2(new_n837), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n302), .B(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT118), .ZN(new_n1134));
  OAI21_X1  g0934(.A(G330), .B1(new_n867), .B2(new_n889), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n901), .A2(new_n1135), .A3(new_n916), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n916), .B2(new_n901), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1135), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n917), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1134), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n901), .A2(new_n1135), .A3(new_n916), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1133), .A2(new_n714), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n723), .B1(new_n1124), .B2(G50), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n976), .A2(G58), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n202), .B2(new_n740), .C1(new_n795), .C2(new_n753), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n390), .A2(G41), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT117), .Z(new_n1151));
  OAI22_X1  g0951(.A1(new_n747), .A2(new_n453), .B1(new_n750), .B2(new_n336), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G68), .B2(new_n767), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G97), .A2(new_n736), .B1(new_n729), .B2(G116), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT58), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n747), .A2(new_n1112), .B1(new_n750), .B2(new_n1113), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G150), .B2(new_n767), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1119), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n736), .A2(G132), .B1(new_n741), .B2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(new_n1120), .C2(new_n730), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(G33), .A2(G41), .ZN(new_n1165));
  INV_X1    g0965(.A(G124), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1165), .B1(new_n753), .B2(new_n1166), .C1(new_n803), .C2(new_n744), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1163), .B2(KEYINPUT59), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1165), .A2(G50), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1164), .A2(new_n1168), .B1(new_n1149), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1157), .A2(new_n1158), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1146), .B1(new_n1171), .B2(new_n717), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1144), .A2(new_n722), .B1(new_n1145), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1067), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1103), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT119), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1103), .A2(new_n1178), .A3(new_n1175), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n666), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1103), .A2(new_n1178), .A3(new_n1175), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1178), .B1(new_n1103), .B2(new_n1175), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1144), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n1181), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1174), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(G375));
  AOI21_X1  g0989(.A(new_n721), .B1(new_n1083), .B2(new_n1074), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT120), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT120), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n723), .B1(new_n1124), .B2(G68), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n730), .A2(new_n732), .B1(new_n740), .B2(new_n502), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1021), .B(new_n1194), .C1(G116), .C2(new_n736), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n341), .A2(new_n750), .B1(new_n747), .B2(new_n795), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n251), .B(new_n1196), .C1(G303), .C2(new_n754), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(new_n202), .C2(new_n791), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n734), .A2(new_n238), .B1(new_n750), .B2(new_n277), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT121), .Z(new_n1200));
  OAI22_X1  g1000(.A1(new_n730), .A2(new_n1117), .B1(new_n740), .B2(new_n803), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n736), .B2(new_n1161), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n979), .A2(G137), .B1(new_n754), .B2(G128), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n390), .A3(new_n1147), .A4(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1198), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1193), .B1(new_n1205), .B2(new_n717), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1082), .B2(new_n715), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1191), .A2(new_n1192), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n949), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1083), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1085), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1208), .A2(new_n1211), .ZN(G381));
  OR4_X1    g1012(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1104), .A2(new_n1128), .A3(KEYINPUT122), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT122), .B1(new_n1104), .B2(new_n1128), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1213), .A2(new_n1217), .A3(G387), .A4(G381), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1188), .ZN(G407));
  INV_X1    g1019(.A(G213), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(G343), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1188), .A2(new_n1216), .A3(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT123), .Z(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1024(.A(G390), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G387), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(G390), .A2(new_n973), .A3(new_n995), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(G393), .B(new_n775), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT125), .B1(G387), .B2(new_n1225), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1229), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1226), .A2(new_n1232), .A3(KEYINPUT125), .A4(new_n1227), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1210), .B1(new_n1084), .B2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1083), .A2(new_n1067), .A3(new_n1074), .A4(KEYINPUT60), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n665), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT124), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1208), .A2(new_n1239), .B1(new_n1240), .B2(G384), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1240), .B2(G384), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1208), .A2(KEYINPUT124), .A3(new_n1243), .A4(new_n1239), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1221), .A2(G2897), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1242), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1173), .B1(new_n1186), .B2(new_n949), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1188), .A2(G378), .B1(new_n1216), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1250), .B2(new_n1221), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT57), .B1(new_n1180), .B2(new_n1144), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1182), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n665), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G378), .B(new_n1173), .C1(new_n1253), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1216), .A2(new_n1249), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1221), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1251), .A2(new_n1252), .A3(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1221), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1265), .B2(new_n1261), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1235), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1261), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT61), .B1(new_n1269), .B2(new_n1248), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1261), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1234), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1274), .ZN(G405));
  NAND2_X1  g1075(.A1(new_n1234), .A2(new_n1270), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1231), .A2(new_n1261), .A3(new_n1233), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1256), .B1(new_n1188), .B2(new_n1217), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1278), .B(new_n1279), .ZN(G402));
endmodule


