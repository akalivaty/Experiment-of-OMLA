

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578;

  XNOR2_X1 U319 ( .A(n428), .B(KEYINPUT118), .ZN(n429) );
  XOR2_X1 U320 ( .A(KEYINPUT28), .B(n450), .Z(n511) );
  XOR2_X1 U321 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n287) );
  XNOR2_X1 U322 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U323 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U324 ( .A(n430), .B(n429), .ZN(n442) );
  XOR2_X1 U325 ( .A(n568), .B(KEYINPUT41), .Z(n547) );
  XOR2_X1 U326 ( .A(n441), .B(n440), .Z(n520) );
  XNOR2_X1 U327 ( .A(n408), .B(n407), .ZN(n558) );
  XNOR2_X1 U328 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n443) );
  XNOR2_X1 U329 ( .A(n444), .B(n443), .ZN(G1348GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n289) );
  XNOR2_X1 U331 ( .A(G22GAT), .B(G197GAT), .ZN(n288) );
  XOR2_X1 U332 ( .A(n289), .B(n288), .Z(n306) );
  XOR2_X1 U333 ( .A(G141GAT), .B(G15GAT), .Z(n291) );
  XNOR2_X1 U334 ( .A(G169GAT), .B(G113GAT), .ZN(n290) );
  XNOR2_X1 U335 ( .A(n291), .B(n290), .ZN(n293) );
  XOR2_X1 U336 ( .A(G43GAT), .B(G50GAT), .Z(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n302) );
  XNOR2_X1 U338 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n294), .B(KEYINPUT67), .ZN(n295) );
  XOR2_X1 U340 ( .A(n295), .B(KEYINPUT65), .Z(n300) );
  XOR2_X1 U341 ( .A(G29GAT), .B(G36GAT), .Z(n297) );
  XNOR2_X1 U342 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n337) );
  XNOR2_X1 U344 ( .A(G8GAT), .B(G1GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n298), .B(KEYINPUT68), .ZN(n362) );
  XNOR2_X1 U346 ( .A(n337), .B(n362), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n304) );
  NAND2_X1 U349 ( .A1(G229GAT), .A2(G233GAT), .ZN(n303) );
  XOR2_X1 U350 ( .A(n304), .B(n303), .Z(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n562) );
  INV_X1 U352 ( .A(KEYINPUT54), .ZN(n385) );
  XOR2_X1 U353 ( .A(G176GAT), .B(G183GAT), .Z(n308) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U356 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n310) );
  XNOR2_X1 U357 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U359 ( .A(n312), .B(n311), .Z(n440) );
  XNOR2_X1 U360 ( .A(G211GAT), .B(G218GAT), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n313), .B(KEYINPUT86), .ZN(n314) );
  XOR2_X1 U362 ( .A(n314), .B(KEYINPUT21), .Z(n316) );
  XNOR2_X1 U363 ( .A(G197GAT), .B(G204GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n421) );
  XNOR2_X1 U365 ( .A(n440), .B(n421), .ZN(n323) );
  XOR2_X1 U366 ( .A(KEYINPUT94), .B(G92GAT), .Z(n318) );
  XNOR2_X1 U367 ( .A(G36GAT), .B(G8GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U369 ( .A(G64GAT), .B(n319), .Z(n321) );
  NAND2_X1 U370 ( .A1(G226GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U372 ( .A(n323), .B(n322), .Z(n507) );
  INV_X1 U373 ( .A(n507), .ZN(n383) );
  XOR2_X1 U374 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n325) );
  XNOR2_X1 U375 ( .A(G190GAT), .B(G99GAT), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U377 ( .A(G85GAT), .B(G92GAT), .Z(n343) );
  XOR2_X1 U378 ( .A(KEYINPUT9), .B(n343), .Z(n327) );
  XOR2_X1 U379 ( .A(G43GAT), .B(G134GAT), .Z(n436) );
  XNOR2_X1 U380 ( .A(n436), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U382 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U383 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U385 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n333) );
  XNOR2_X1 U386 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U388 ( .A(n335), .B(n334), .Z(n339) );
  XNOR2_X1 U389 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n336), .B(G162GAT), .ZN(n409) );
  XNOR2_X1 U391 ( .A(n337), .B(n409), .ZN(n338) );
  XOR2_X1 U392 ( .A(n339), .B(n338), .Z(n551) );
  INV_X1 U393 ( .A(n551), .ZN(n542) );
  XOR2_X1 U394 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n341) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G204GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n356) );
  XNOR2_X1 U397 ( .A(G57GAT), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n287), .B(n342), .ZN(n358) );
  XNOR2_X1 U399 ( .A(n358), .B(n343), .ZN(n345) );
  AND2_X1 U400 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n354) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G71GAT), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n346), .B(G120GAT), .ZN(n431) );
  XOR2_X1 U404 ( .A(G78GAT), .B(G148GAT), .Z(n348) );
  XNOR2_X1 U405 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n418) );
  XNOR2_X1 U407 ( .A(n431), .B(n418), .ZN(n352) );
  XOR2_X1 U408 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n350) );
  XNOR2_X1 U409 ( .A(KEYINPUT71), .B(KEYINPUT73), .ZN(n349) );
  XOR2_X1 U410 ( .A(n350), .B(n349), .Z(n351) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n568) );
  NOR2_X1 U412 ( .A1(n562), .A2(n547), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n357), .B(KEYINPUT46), .ZN(n373) );
  XOR2_X1 U414 ( .A(n358), .B(KEYINPUT79), .Z(n360) );
  NAND2_X1 U415 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U417 ( .A(G22GAT), .B(G155GAT), .Z(n415) );
  XOR2_X1 U418 ( .A(n361), .B(n415), .Z(n364) );
  XOR2_X1 U419 ( .A(G15GAT), .B(G127GAT), .Z(n434) );
  XNOR2_X1 U420 ( .A(n362), .B(n434), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n372) );
  XOR2_X1 U422 ( .A(G78GAT), .B(G211GAT), .Z(n366) );
  XNOR2_X1 U423 ( .A(G183GAT), .B(G71GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U425 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n368) );
  XNOR2_X1 U426 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U428 ( .A(n370), .B(n369), .Z(n371) );
  XOR2_X1 U429 ( .A(n372), .B(n371), .Z(n572) );
  INV_X1 U430 ( .A(n572), .ZN(n540) );
  NOR2_X1 U431 ( .A1(n373), .A2(n540), .ZN(n374) );
  XOR2_X1 U432 ( .A(KEYINPUT114), .B(n374), .Z(n375) );
  NOR2_X1 U433 ( .A1(n542), .A2(n375), .ZN(n376) );
  XNOR2_X1 U434 ( .A(KEYINPUT47), .B(n376), .ZN(n381) );
  INV_X1 U435 ( .A(n562), .ZN(n534) );
  XNOR2_X1 U436 ( .A(KEYINPUT36), .B(n551), .ZN(n575) );
  NOR2_X1 U437 ( .A1(n575), .A2(n572), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n377), .B(KEYINPUT45), .ZN(n378) );
  NAND2_X1 U439 ( .A1(n378), .A2(n568), .ZN(n379) );
  OR2_X1 U440 ( .A1(n534), .A2(n379), .ZN(n380) );
  AND2_X1 U441 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U442 ( .A(KEYINPUT48), .B(n382), .ZN(n517) );
  NOR2_X1 U443 ( .A1(n383), .A2(n517), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n557) );
  XOR2_X1 U445 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n387) );
  XNOR2_X1 U446 ( .A(KEYINPUT5), .B(KEYINPUT93), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n400) );
  XOR2_X1 U448 ( .A(G57GAT), .B(G155GAT), .Z(n389) );
  XNOR2_X1 U449 ( .A(G1GAT), .B(G148GAT), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U451 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n391) );
  XNOR2_X1 U452 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U454 ( .A(n393), .B(n392), .Z(n398) );
  XOR2_X1 U455 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n395) );
  XNOR2_X1 U456 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n437) );
  XNOR2_X1 U458 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n396), .B(KEYINPUT2), .ZN(n420) );
  XNOR2_X1 U460 ( .A(n437), .B(n420), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n408) );
  NAND2_X1 U463 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XOR2_X1 U464 ( .A(G162GAT), .B(G120GAT), .Z(n402) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(G127GAT), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U467 ( .A(G134GAT), .B(G85GAT), .Z(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  INV_X1 U470 ( .A(n558), .ZN(n426) );
  XOR2_X1 U471 ( .A(KEYINPUT24), .B(n409), .Z(n411) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n425) );
  XOR2_X1 U474 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n413) );
  XNOR2_X1 U475 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U477 ( .A(n414), .B(KEYINPUT89), .Z(n417) );
  XNOR2_X1 U478 ( .A(n415), .B(KEYINPUT85), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U480 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n450) );
  NAND2_X1 U484 ( .A1(n426), .A2(n450), .ZN(n427) );
  NOR2_X1 U485 ( .A1(n557), .A2(n427), .ZN(n430) );
  INV_X1 U486 ( .A(KEYINPUT55), .ZN(n428) );
  XOR2_X1 U487 ( .A(KEYINPUT20), .B(n431), .Z(n433) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n441) );
  NAND2_X1 U493 ( .A1(n442), .A2(n520), .ZN(n552) );
  NOR2_X1 U494 ( .A1(n562), .A2(n552), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n462) );
  AND2_X1 U496 ( .A1(n568), .A2(n534), .ZN(n479) );
  INV_X1 U497 ( .A(n511), .ZN(n519) );
  XOR2_X1 U498 ( .A(n507), .B(KEYINPUT27), .Z(n516) );
  XNOR2_X1 U499 ( .A(KEYINPUT84), .B(n520), .ZN(n445) );
  NOR2_X1 U500 ( .A1(n516), .A2(n445), .ZN(n446) );
  NAND2_X1 U501 ( .A1(n519), .A2(n446), .ZN(n447) );
  NAND2_X1 U502 ( .A1(n447), .A2(n558), .ZN(n457) );
  NAND2_X1 U503 ( .A1(n520), .A2(n507), .ZN(n448) );
  NAND2_X1 U504 ( .A1(n450), .A2(n448), .ZN(n449) );
  XOR2_X1 U505 ( .A(KEYINPUT25), .B(n449), .Z(n455) );
  NOR2_X1 U506 ( .A1(n520), .A2(n450), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT95), .B(n451), .Z(n452) );
  XOR2_X1 U508 ( .A(KEYINPUT26), .B(n452), .Z(n556) );
  NOR2_X1 U509 ( .A1(n556), .A2(n516), .ZN(n453) );
  NOR2_X1 U510 ( .A1(n558), .A2(n453), .ZN(n454) );
  NAND2_X1 U511 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U512 ( .A1(n457), .A2(n456), .ZN(n475) );
  NAND2_X1 U513 ( .A1(n540), .A2(n551), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n458), .B(KEYINPUT80), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT16), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n475), .A2(n460), .ZN(n492) );
  AND2_X1 U517 ( .A1(n479), .A2(n492), .ZN(n470) );
  NAND2_X1 U518 ( .A1(n470), .A2(n558), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U520 ( .A(G1GAT), .B(n463), .Z(G1324GAT) );
  XOR2_X1 U521 ( .A(G8GAT), .B(KEYINPUT97), .Z(n465) );
  NAND2_X1 U522 ( .A1(n470), .A2(n507), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n465), .B(n464), .ZN(G1325GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n467) );
  NAND2_X1 U525 ( .A1(n470), .A2(n520), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(n469) );
  XOR2_X1 U527 ( .A(G15GAT), .B(KEYINPUT98), .Z(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(G1326GAT) );
  NAND2_X1 U529 ( .A1(n511), .A2(n470), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n473) );
  XNOR2_X1 U532 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT100), .B(n474), .Z(n483) );
  XOR2_X1 U535 ( .A(KEYINPUT38), .B(KEYINPUT102), .Z(n481) );
  NOR2_X1 U536 ( .A1(n575), .A2(n475), .ZN(n476) );
  NAND2_X1 U537 ( .A1(n572), .A2(n476), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT37), .B(KEYINPUT101), .Z(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n504) );
  NAND2_X1 U540 ( .A1(n479), .A2(n504), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n489) );
  NAND2_X1 U542 ( .A1(n489), .A2(n558), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(G1328GAT) );
  XOR2_X1 U544 ( .A(G36GAT), .B(KEYINPUT105), .Z(n485) );
  NAND2_X1 U545 ( .A1(n489), .A2(n507), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(G1329GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n487) );
  NAND2_X1 U548 ( .A1(n489), .A2(n520), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U550 ( .A(G43GAT), .B(n488), .Z(G1330GAT) );
  XOR2_X1 U551 ( .A(G50GAT), .B(KEYINPUT107), .Z(n491) );
  NAND2_X1 U552 ( .A1(n489), .A2(n511), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1331GAT) );
  NOR2_X1 U554 ( .A1(n534), .A2(n547), .ZN(n503) );
  AND2_X1 U555 ( .A1(n503), .A2(n492), .ZN(n499) );
  NAND2_X1 U556 ( .A1(n558), .A2(n499), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n494) );
  XNOR2_X1 U558 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(G1332GAT) );
  NAND2_X1 U561 ( .A1(n507), .A2(n499), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n497), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U563 ( .A1(n499), .A2(n520), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n498), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n501) );
  NAND2_X1 U566 ( .A1(n499), .A2(n511), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(n502), .ZN(G1335GAT) );
  XOR2_X1 U569 ( .A(G85GAT), .B(KEYINPUT111), .Z(n506) );
  AND2_X1 U570 ( .A1(n504), .A2(n503), .ZN(n512) );
  NAND2_X1 U571 ( .A1(n512), .A2(n558), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1336GAT) );
  NAND2_X1 U573 ( .A1(n507), .A2(n512), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n520), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(KEYINPUT112), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G99GAT), .B(n510), .ZN(G1338GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G106GAT), .B(n515), .ZN(G1339GAT) );
  NOR2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n518) );
  NAND2_X1 U583 ( .A1(n518), .A2(n558), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U585 ( .A1(n533), .A2(n521), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n530), .A2(n534), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n524) );
  INV_X1 U589 ( .A(n547), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n530), .A2(n536), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U592 ( .A(G120GAT), .B(n525), .Z(G1341GAT) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n527) );
  NAND2_X1 U595 ( .A1(n530), .A2(n540), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .Z(n532) );
  NAND2_X1 U599 ( .A1(n530), .A2(n542), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(G1343GAT) );
  NOR2_X1 U601 ( .A1(n556), .A2(n533), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n534), .A2(n543), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(n535), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n538) );
  NAND2_X1 U605 ( .A1(n543), .A2(n536), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(n539), .ZN(G1345GAT) );
  NAND2_X1 U608 ( .A1(n540), .A2(n543), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n541), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n544), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n546) );
  XNOR2_X1 U613 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n549) );
  NOR2_X1 U615 ( .A1(n547), .A2(n552), .ZN(n548) );
  XOR2_X1 U616 ( .A(n549), .B(n548), .Z(G1349GAT) );
  NOR2_X1 U617 ( .A1(n572), .A2(n552), .ZN(n550) );
  XOR2_X1 U618 ( .A(G183GAT), .B(n550), .Z(G1350GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT121), .B(KEYINPUT58), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G190GAT), .B(n555), .ZN(G1351GAT) );
  INV_X1 U623 ( .A(n556), .ZN(n560) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT122), .ZN(n574) );
  NOR2_X1 U627 ( .A1(n574), .A2(n562), .ZN(n564) );
  XNOR2_X1 U628 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(n565), .ZN(G1352GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n567) );
  XNOR2_X1 U632 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n574), .A2(n568), .ZN(n569) );
  XOR2_X1 U635 ( .A(n570), .B(n569), .Z(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT123), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n574), .ZN(n573) );
  XOR2_X1 U638 ( .A(G211GAT), .B(n573), .Z(G1354GAT) );
  XNOR2_X1 U639 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n577) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(G218GAT), .B(n578), .Z(G1355GAT) );
endmodule

