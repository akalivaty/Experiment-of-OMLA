//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(new_n461), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n470), .A2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT71), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(KEYINPUT70), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(KEYINPUT70), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n482), .A2(new_n483), .B1(new_n472), .B2(new_n471), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n482), .A2(new_n483), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(G136), .B2(new_n488), .ZN(G162));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n468), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n473), .A2(new_n481), .A3(new_n496), .A4(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OR2_X1    g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n500), .A2(new_n501), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT72), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n503), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(G62), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(new_n522), .B1(G75), .B2(G543), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n514), .A2(KEYINPUT73), .A3(G62), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT7), .Z(new_n528));
  AND3_X1   g103(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n529));
  AOI211_X1 g104(.A(new_n528), .B(new_n529), .C1(G51), .C2(new_n502), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n511), .A2(new_n516), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n507), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G651), .B1(G52), .B2(new_n502), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n517), .B2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n507), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G651), .B1(G43), .B2(new_n502), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n517), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT75), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n502), .A2(new_n557), .A3(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n531), .A2(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n514), .B(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n520), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND3_X1  g143(.A1(new_n511), .A2(G87), .A3(new_n516), .ZN(new_n569));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n512), .A2(new_n570), .A3(new_n513), .ZN(new_n571));
  AOI22_X1  g146(.A1(G49), .A2(new_n502), .B1(new_n571), .B2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n507), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G48), .B2(new_n502), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n517), .B2(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(new_n502), .A2(G47), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  OAI221_X1 g157(.A(new_n580), .B1(new_n520), .B2(new_n581), .C1(new_n517), .C2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n531), .A2(G92), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G79), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT79), .B1(new_n588), .B2(new_n499), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n588), .A2(new_n499), .A3(KEYINPUT79), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n507), .B(KEYINPUT77), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n502), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(KEYINPUT78), .ZN(new_n595));
  INV_X1    g170(.A(G54), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n594), .B2(KEYINPUT78), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n593), .A2(G651), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n584), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n584), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n566), .B2(G868), .ZN(G297));
  XNOR2_X1  g179(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n600), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n600), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n488), .A2(G135), .ZN(new_n612));
  INV_X1    g187(.A(new_n484), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G123), .ZN(new_n614));
  OAI221_X1 g189(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G2096), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(G2096), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT83), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2427), .B(G2430), .Z(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n630), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT82), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n634), .A2(new_n638), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(G401));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT84), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n642), .B1(new_n644), .B2(KEYINPUT85), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(KEYINPUT85), .B2(new_n644), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2084), .B(G2090), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n644), .B(KEYINPUT17), .Z(new_n648));
  INV_X1    g223(.A(new_n642), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n642), .A2(new_n647), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n660), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n660), .B2(new_n666), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1981), .B(G1986), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G32), .ZN(new_n678));
  NAND3_X1  g253(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT95), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT26), .Z(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n488), .B2(G141), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT94), .Z(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n613), .B2(G129), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n678), .B1(new_n687), .B2(new_n677), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT96), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT27), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n677), .A2(G35), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G162), .B2(new_n677), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT29), .B(G2090), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT30), .B(G28), .ZN(new_n696));
  OR2_X1    g271(.A1(KEYINPUT31), .A2(G11), .ZN(new_n697));
  NAND2_X1  g272(.A1(KEYINPUT31), .A2(G11), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n696), .A2(new_n677), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n616), .B2(new_n677), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT98), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NOR2_X1   g278(.A1(G168), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n703), .B2(G21), .ZN(new_n705));
  INV_X1    g280(.A(G1966), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT97), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n677), .A2(G26), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n488), .A2(G140), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n613), .A2(G128), .ZN(new_n712));
  OAI221_X1 g287(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n710), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT93), .B(G2067), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n691), .A2(new_n702), .A3(new_n708), .A4(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT24), .ZN(new_n719));
  INV_X1    g294(.A(G34), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G160), .B2(new_n677), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2084), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n488), .A2(G139), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT25), .Z(new_n727));
  AOI22_X1  g302(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n725), .B(new_n727), .C1(new_n473), .C2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G33), .B(new_n729), .S(G29), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2072), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n724), .B(new_n731), .C1(new_n706), .C2(new_n705), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n703), .A2(G20), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT23), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n566), .B2(new_n703), .ZN(new_n735));
  INV_X1    g310(.A(G1956), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G171), .A2(new_n703), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G5), .B2(new_n703), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT99), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n677), .A2(G27), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT100), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n677), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n743), .B1(G2078), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G2078), .B2(new_n746), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n732), .A2(new_n737), .A3(new_n742), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G4), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n600), .B2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT91), .B(G1348), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n703), .A2(G19), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT92), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n550), .B2(new_n703), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n718), .A2(new_n749), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(G25), .A2(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n488), .A2(G131), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n473), .A2(G107), .ZN(new_n761));
  OAI21_X1  g336(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n613), .A2(G119), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(KEYINPUT87), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(KEYINPUT87), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n760), .B1(new_n761), .B2(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n677), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT35), .B(G1991), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n770));
  MUX2_X1   g345(.A(G24), .B(G290), .S(G16), .Z(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G1986), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n769), .B(new_n772), .C1(G1986), .C2(new_n771), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n767), .A2(new_n768), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G23), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n569), .A2(KEYINPUT88), .A3(new_n572), .ZN(new_n777));
  AOI21_X1  g352(.A(KEYINPUT88), .B1(new_n569), .B2(new_n572), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n776), .B1(new_n779), .B2(G16), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT33), .B(G1976), .Z(new_n781));
  XOR2_X1   g356(.A(new_n780), .B(new_n781), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n703), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n703), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G6), .B(G305), .S(G16), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n782), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(KEYINPUT89), .B1(new_n790), .B2(KEYINPUT34), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n790), .A2(KEYINPUT89), .A3(KEYINPUT34), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n775), .B1(KEYINPUT34), .B2(new_n790), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n758), .A2(new_n796), .A3(new_n797), .ZN(G150));
  INV_X1    g373(.A(G150), .ZN(G311));
  NAND2_X1  g374(.A1(new_n502), .A2(G55), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  INV_X1    g376(.A(G93), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n800), .B1(new_n520), .B2(new_n801), .C1(new_n517), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G860), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT102), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT37), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n549), .A2(new_n803), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n547), .B2(new_n803), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n600), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT101), .ZN(new_n814));
  INV_X1    g389(.A(G860), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n812), .B2(KEYINPUT39), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n806), .B1(new_n814), .B2(new_n816), .ZN(G145));
  OAI221_X1 g392(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n473), .C2(G118), .ZN(new_n818));
  INV_X1    g393(.A(G130), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n484), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G142), .B2(new_n488), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT103), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n620), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n686), .B(new_n729), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n714), .B(G164), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n766), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n616), .B(G160), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G162), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(G37), .B1(new_n828), .B2(new_n830), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n832), .A2(KEYINPUT40), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT40), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(G395));
  XNOR2_X1  g411(.A(new_n599), .B(G299), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n599), .B(new_n566), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT41), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n608), .B(new_n808), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G166), .B(KEYINPUT105), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G305), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n779), .B(G290), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT106), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n849), .A2(new_n850), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n848), .A2(new_n853), .A3(new_n851), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT42), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n844), .A2(new_n837), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n852), .A2(new_n854), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT42), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND4_X1   g435(.A1(new_n846), .A2(new_n856), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n856), .A2(new_n860), .B1(new_n846), .B2(new_n857), .ZN(new_n862));
  OAI21_X1  g437(.A(G868), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n864));
  INV_X1    g439(.A(G868), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n803), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n863), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(G295));
  NAND2_X1  g444(.A1(new_n863), .A2(new_n866), .ZN(G331));
  XNOR2_X1  g445(.A(G286), .B(G171), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n808), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n840), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n843), .B2(new_n872), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n855), .B1(new_n874), .B2(KEYINPUT108), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(KEYINPUT108), .B2(new_n874), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n874), .B2(new_n858), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT43), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n873), .B(KEYINPUT110), .ZN(new_n881));
  INV_X1    g456(.A(new_n872), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n837), .A2(KEYINPUT41), .ZN(new_n883));
  OAI22_X1  g458(.A1(new_n883), .A2(KEYINPUT109), .B1(new_n837), .B2(new_n838), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n883), .A2(KEYINPUT109), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n855), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n887), .A2(new_n878), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT44), .B1(new_n880), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n876), .B2(new_n879), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n887), .A2(new_n878), .A3(KEYINPUT43), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n890), .B1(new_n893), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g469(.A1(new_n495), .A2(new_n497), .ZN(new_n895));
  INV_X1    g470(.A(new_n493), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G1384), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT45), .ZN(new_n900));
  INV_X1    g475(.A(G40), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n470), .A2(new_n476), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n686), .B(G1996), .Z(new_n904));
  XOR2_X1   g479(.A(new_n714), .B(G2067), .Z(new_n905));
  AND2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n768), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n766), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n766), .A2(new_n907), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(G290), .B(G1986), .Z(new_n911));
  AOI21_X1  g486(.A(new_n903), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n902), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(new_n899), .B2(KEYINPUT50), .ZN(new_n914));
  INV_X1    g489(.A(G2090), .ZN(new_n915));
  AOI21_X1  g490(.A(G1384), .B1(new_n895), .B2(new_n896), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT50), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT111), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n919));
  NOR4_X1   g494(.A1(G164), .A2(new_n919), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n914), .B(new_n915), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(KEYINPUT45), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n900), .B1(G164), .B2(G1384), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n902), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n785), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(G8), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n928));
  OAI211_X1 g503(.A(G8), .B(new_n928), .C1(new_n519), .C2(new_n525), .ZN(new_n929));
  INV_X1    g504(.A(G8), .ZN(new_n930));
  NOR2_X1   g505(.A1(G166), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G2084), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n914), .B(new_n936), .C1(new_n918), .C2(new_n920), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n924), .A2(new_n706), .ZN(new_n938));
  AOI211_X1 g513(.A(new_n930), .B(G286), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(KEYINPUT63), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1976), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n777), .A2(new_n778), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(G8), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT52), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n778), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n569), .A2(KEYINPUT88), .A3(new_n572), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(G1976), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n930), .B1(new_n916), .B2(new_n902), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT52), .B1(G288), .B2(new_n941), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n511), .A2(G86), .A3(new_n516), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n502), .A2(G48), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(new_n520), .ZN(new_n956));
  OAI21_X1  g531(.A(G1981), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1981), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n577), .B(new_n958), .C1(new_n578), .C2(new_n517), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(G305), .A2(KEYINPUT113), .A3(G1981), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT49), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n966), .A2(new_n949), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n952), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n926), .A2(G8), .A3(new_n933), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT115), .B1(new_n940), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n970), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n939), .A2(KEYINPUT63), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n935), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n897), .A2(new_n917), .A3(new_n898), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n976), .A2(new_n902), .A3(new_n977), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n978), .A2(new_n915), .B1(new_n924), .B2(new_n785), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n934), .B1(new_n979), .B2(new_n930), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n968), .A2(new_n939), .A3(new_n969), .A4(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT63), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n981), .A2(KEYINPUT114), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT114), .B1(new_n981), .B2(new_n982), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n971), .B(new_n975), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(G286), .A2(G8), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n986), .B2(KEYINPUT122), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n977), .A2(new_n902), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n976), .A2(new_n919), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n916), .A2(KEYINPUT111), .A3(new_n917), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n991), .A2(new_n936), .B1(new_n706), .B2(new_n924), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n986), .B(new_n987), .C1(new_n992), .C2(new_n930), .ZN(new_n993));
  INV_X1    g568(.A(new_n987), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n937), .A2(new_n938), .ZN(new_n995));
  OAI211_X1 g570(.A(G8), .B(new_n994), .C1(new_n995), .C2(G286), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT121), .B1(new_n992), .B2(new_n986), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT121), .ZN(new_n999));
  INV_X1    g574(.A(new_n986), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n997), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n918), .A2(new_n920), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT118), .B1(new_n1007), .B2(new_n988), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n914), .B(new_n1009), .C1(new_n918), .C2(new_n920), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n740), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n924), .B2(G2078), .ZN(new_n1013));
  OR3_X1    g588(.A1(new_n924), .A2(new_n1012), .A3(G2078), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G171), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n968), .A2(new_n980), .A3(new_n969), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1004), .A2(new_n1006), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n967), .A2(new_n964), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1020), .A2(new_n941), .A3(new_n569), .A4(new_n572), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n944), .B1(new_n1021), .B2(new_n959), .ZN(new_n1022));
  INV_X1    g597(.A(new_n969), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(new_n968), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n985), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1348), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1008), .A2(new_n1026), .A3(new_n1010), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n943), .A2(G2067), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT117), .Z(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n922), .A2(new_n923), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT56), .B(G2072), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n902), .A4(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT57), .B1(new_n561), .B2(new_n565), .ZN(new_n1035));
  INV_X1    g610(.A(G65), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n591), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n564), .ZN(new_n1038));
  OAI21_X1  g613(.A(G651), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n559), .A4(new_n560), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1035), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n922), .A2(new_n902), .A3(new_n923), .A4(new_n1033), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1044));
  INV_X1    g619(.A(new_n976), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n736), .B1(new_n1045), .B2(new_n988), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1034), .A2(new_n1042), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1030), .A2(new_n600), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1034), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1034), .A2(KEYINPUT119), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1042), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT60), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n600), .B2(KEYINPUT120), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n600), .A2(KEYINPUT120), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1030), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1060), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(KEYINPUT60), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1058), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT58), .B(G1341), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n943), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n924), .B2(G1996), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n550), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1069), .B2(new_n550), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1047), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT61), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1047), .A2(KEYINPUT61), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1054), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1056), .B1(new_n1066), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1017), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1003), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT123), .B1(new_n474), .B2(new_n475), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(new_n473), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n474), .A2(KEYINPUT123), .A3(new_n475), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR4_X1   g663(.A1(new_n470), .A2(new_n1012), .A3(new_n901), .A4(G2078), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1031), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1011), .A2(G301), .A3(new_n1013), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT54), .B1(new_n1016), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1011), .A2(new_n1013), .A3(new_n1090), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1011), .A2(KEYINPUT124), .A3(new_n1013), .A4(new_n1090), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(G171), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1011), .A2(G301), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1099), .A2(KEYINPUT54), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1098), .A2(KEYINPUT125), .A3(new_n1100), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1082), .A2(new_n1093), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n912), .B1(new_n1025), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n903), .B1(new_n905), .B2(new_n687), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT46), .B1(new_n903), .B2(G1996), .ZN(new_n1108));
  OR3_X1    g683(.A1(new_n903), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT47), .Z(new_n1111));
  NOR3_X1   g686(.A1(new_n903), .A2(G1986), .A3(G290), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n1112), .B(KEYINPUT48), .Z(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n910), .B2(new_n903), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n908), .A2(KEYINPUT126), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n906), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n908), .A2(KEYINPUT126), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1116), .A2(new_n1117), .B1(G2067), .B2(new_n714), .ZN(new_n1118));
  INV_X1    g693(.A(new_n903), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1111), .A2(new_n1114), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT127), .B1(new_n1106), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT127), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1121), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n983), .A2(new_n984), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n975), .A2(new_n971), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1019), .B(new_n1024), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1042), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1078), .B1(new_n1128), .B2(new_n1052), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT61), .B1(new_n1074), .B2(new_n1047), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1129), .A2(new_n1130), .A3(new_n1073), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1063), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1060), .B1(new_n1030), .B2(new_n1057), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1030), .A2(new_n1059), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1055), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1127), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1123), .B(new_n1124), .C1(new_n1140), .C2(new_n912), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1122), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g717(.A(G319), .ZN(new_n1144));
  NOR4_X1   g718(.A1(G229), .A2(new_n1144), .A3(G401), .A4(G227), .ZN(new_n1145));
  NAND2_X1  g719(.A1(new_n828), .A2(new_n830), .ZN(new_n1146));
  NAND2_X1  g720(.A1(new_n1146), .A2(new_n877), .ZN(new_n1147));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1147), .B2(new_n831), .ZN(new_n1148));
  NOR2_X1   g722(.A1(new_n1148), .A2(new_n893), .ZN(G308));
  OAI221_X1 g723(.A(new_n1145), .B1(new_n1147), .B2(new_n831), .C1(new_n891), .C2(new_n892), .ZN(G225));
endmodule


