//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  AND2_X1   g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(KEYINPUT22), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G211gat), .A2(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n204), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208));
  XNOR2_X1  g007(.A(G141gat), .B(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n210), .B1(G155gat), .B2(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n209), .A2(new_n211), .B1(KEYINPUT80), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G155gat), .B(G162gat), .Z(new_n216));
  AND2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n208), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT29), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n207), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n207), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n208), .B1(new_n222), .B2(KEYINPUT29), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n217), .A2(new_n218), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G78gat), .B(G106gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G228gat), .A2(G233gat), .ZN(new_n228));
  INV_X1    g027(.A(G22gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT31), .B(G50gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n227), .A2(new_n232), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G1gat), .B(G29gat), .Z(new_n237));
  XNOR2_X1  g036(.A(G57gat), .B(G85gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT86), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n243));
  INV_X1    g042(.A(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G113gat), .ZN(new_n245));
  INV_X1    g044(.A(G113gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G120gat), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT1), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G127gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G134gat), .ZN(new_n250));
  INV_X1    g049(.A(G134gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G127gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n252), .B2(KEYINPUT72), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n248), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n253), .B2(new_n254), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT74), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n246), .B2(G120gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(KEYINPUT74), .A3(G113gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n247), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n250), .A4(new_n252), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT75), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n256), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n243), .A2(new_n266), .A3(new_n219), .ZN(new_n267));
  OAI221_X1 g066(.A(new_n256), .B1(new_n217), .B2(new_n218), .C1(new_n264), .C2(new_n265), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(KEYINPUT4), .A3(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n268), .A2(KEYINPUT4), .ZN(new_n270));
  NAND2_X1  g069(.A1(G225gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT87), .B(KEYINPUT39), .Z(new_n275));
  AOI21_X1  g074(.A(new_n242), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n266), .A2(new_n224), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(new_n268), .A3(KEYINPUT81), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n266), .A2(new_n279), .A3(new_n224), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n272), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n273), .A2(KEYINPUT39), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT40), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(KEYINPUT5), .A3(new_n271), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n278), .A2(new_n272), .A3(new_n280), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n271), .A2(new_n286), .B1(new_n289), .B2(KEYINPUT5), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n242), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n283), .A2(new_n284), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT78), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  INV_X1    g098(.A(G226gat), .ZN(new_n300));
  INV_X1    g099(.A(G233gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT29), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  AND2_X1   g104(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n306));
  NOR2_X1   g105(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n307));
  OAI22_X1  g106(.A1(new_n306), .A2(new_n307), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT24), .ZN(new_n313));
  XOR2_X1   g112(.A(G183gat), .B(G190gat), .Z(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(KEYINPUT24), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(KEYINPUT23), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n305), .B1(new_n310), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n308), .B(KEYINPUT66), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n319), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT23), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n318), .A2(new_n305), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n323), .A2(new_n315), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n322), .A2(new_n328), .A3(KEYINPUT68), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n318), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT26), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n319), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n335), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(KEYINPUT71), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n325), .A2(new_n339), .A3(new_n335), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n338), .A2(new_n340), .B1(G183gat), .B2(G190gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT27), .B(G183gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n311), .B2(KEYINPUT27), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n312), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n342), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(KEYINPUT28), .A3(new_n312), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n348), .A2(KEYINPUT70), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT70), .B1(new_n348), .B2(new_n349), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n341), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n304), .B1(new_n333), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n302), .A3(new_n329), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n353), .A2(new_n355), .A3(new_n207), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n333), .A2(new_n302), .A3(new_n352), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n329), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n303), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n222), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n299), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n359), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n207), .ZN(new_n363));
  INV_X1    g162(.A(new_n332), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT68), .B1(new_n322), .B2(new_n328), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n352), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n303), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n222), .A3(new_n354), .ZN(new_n368));
  INV_X1    g167(.A(new_n299), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n363), .A2(KEYINPUT30), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(new_n368), .A3(new_n369), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(KEYINPUT79), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT79), .B1(new_n371), .B2(new_n372), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n361), .B(new_n370), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n236), .B1(new_n295), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n356), .A2(new_n360), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT37), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(KEYINPUT88), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n379), .A3(new_n368), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n353), .A2(new_n355), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n379), .B1(new_n385), .B2(new_n207), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n222), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT38), .B(new_n369), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n299), .B1(new_n378), .B2(new_n379), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n383), .B2(new_n380), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT38), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n371), .B(new_n389), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT89), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n291), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n241), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n286), .A2(new_n271), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n289), .A2(KEYINPUT5), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n398), .A2(KEYINPUT6), .A3(new_n241), .A4(new_n287), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n401), .A3(new_n394), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405));
  INV_X1    g204(.A(new_n241), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n288), .B2(new_n290), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n292), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n403), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n377), .B1(new_n393), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n366), .B2(new_n266), .ZN(new_n413));
  INV_X1    g212(.A(new_n266), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n333), .A2(KEYINPUT76), .A3(new_n414), .A4(new_n352), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n366), .A2(new_n266), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G227gat), .A2(G233gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n418), .B(KEYINPUT64), .Z(new_n419));
  OR2_X1    g218(.A1(new_n419), .A2(KEYINPUT34), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n418), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT34), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT32), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n417), .B2(new_n419), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT33), .B1(new_n417), .B2(new_n419), .ZN(new_n427));
  XOR2_X1   g226(.A(G15gat), .B(G43gat), .Z(new_n428));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n426), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  AOI221_X4 g231(.A(new_n425), .B1(KEYINPUT33), .B2(new_n430), .C1(new_n417), .C2(new_n419), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n424), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n427), .A2(new_n431), .ZN(new_n435));
  INV_X1    g234(.A(new_n426), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(new_n424), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT77), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n434), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n437), .A2(new_n439), .A3(KEYINPUT77), .A4(new_n438), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n291), .A2(new_n241), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n291), .A2(KEYINPUT83), .A3(new_n241), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n405), .A3(new_n450), .A4(new_n407), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n395), .A2(new_n401), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n370), .A2(new_n361), .ZN(new_n455));
  INV_X1    g254(.A(new_n375), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n373), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n235), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n445), .B1(new_n434), .B2(new_n440), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n411), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT36), .B1(new_n442), .B2(new_n443), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(KEYINPUT85), .A3(new_n459), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n454), .A2(new_n457), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n434), .A2(new_n440), .A3(new_n235), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT35), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n457), .A2(new_n471), .A3(new_n235), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n404), .A2(new_n408), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n402), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n444), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n464), .A2(new_n467), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n478));
  INV_X1    g277(.A(G29gat), .ZN(new_n479));
  INV_X1    g278(.A(G36gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G29gat), .A2(G36gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n483), .B(new_n488), .C1(KEYINPUT91), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n483), .B2(new_n488), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT15), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n483), .A2(new_n488), .ZN(new_n498));
  INV_X1    g297(.A(new_n489), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n495), .B1(new_n500), .B2(new_n490), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n490), .A2(new_n495), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT17), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G15gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n229), .ZN(new_n505));
  NAND2_X1  g304(.A1(G15gat), .A2(G22gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT16), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(G1gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G8gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT92), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(G1gat), .A3(new_n506), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n511), .A2(KEYINPUT92), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n515), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n510), .A2(new_n517), .A3(new_n512), .A4(new_n513), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n497), .A2(new_n503), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n501), .A2(new_n502), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523));
  AOI211_X1 g322(.A(KEYINPUT92), .B(new_n511), .C1(new_n510), .C2(new_n513), .ZN(new_n524));
  INV_X1    g323(.A(new_n518), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n516), .A2(KEYINPUT93), .A3(new_n518), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n520), .A2(new_n521), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n520), .A2(KEYINPUT18), .A3(new_n528), .A4(new_n521), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n516), .A2(KEYINPUT93), .A3(new_n518), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT93), .B1(new_n516), .B2(new_n518), .ZN(new_n534));
  OAI22_X1  g333(.A1(new_n533), .A2(new_n534), .B1(new_n501), .B2(new_n502), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n528), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n521), .B(KEYINPUT13), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G197gat), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT11), .B(G169gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT12), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n531), .A2(new_n544), .A3(new_n538), .A4(new_n532), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n477), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT9), .ZN(new_n551));
  INV_X1    g350(.A(G71gat), .ZN(new_n552));
  INV_X1    g351(.A(G78gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT94), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT94), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n556), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  INV_X1    g356(.A(G57gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G64gat), .ZN(new_n559));
  INV_X1    g358(.A(G64gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G57gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n560), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n559), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n570), .A2(new_n555), .A3(new_n564), .A4(new_n557), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n249), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n566), .A2(new_n571), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n526), .A2(new_n527), .B1(new_n578), .B2(KEYINPUT21), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n577), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n212), .ZN(new_n582));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n580), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT100), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT8), .ZN(new_n590));
  OR2_X1    g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n593));
  OR2_X1    g392(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  AND2_X1   g396(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n598));
  NOR2_X1   g397(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n592), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT98), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G99gat), .ZN(new_n605));
  INV_X1    g404(.A(G106gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n589), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT99), .B1(new_n601), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n600), .ZN(new_n612));
  INV_X1    g411(.A(new_n592), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n612), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n613), .ZN(new_n616));
  INV_X1    g415(.A(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n610), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(KEYINPUT99), .A3(new_n619), .ZN(new_n620));
  AND4_X1   g419(.A1(new_n497), .A2(new_n503), .A3(new_n615), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n611), .A2(new_n614), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT99), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n522), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n588), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G134gat), .B(G162gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n587), .A2(KEYINPUT100), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n629), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n588), .B(new_n634), .C1(new_n621), .C2(new_n627), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n630), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n633), .B1(new_n630), .B2(new_n635), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n585), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n615), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n572), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n601), .A2(new_n610), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n619), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n601), .A2(KEYINPUT101), .A3(new_n610), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n578), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT103), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n642), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT104), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n642), .A2(new_n647), .A3(new_n652), .A4(new_n649), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  NAND3_X1  g455(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n649), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n566), .A2(KEYINPUT10), .A3(new_n571), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT102), .B1(new_n641), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n663), .B(new_n660), .C1(new_n620), .C2(new_n615), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT10), .B1(new_n642), .B2(new_n647), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n659), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n658), .A2(KEYINPUT105), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n661), .B1(new_n622), .B2(new_n623), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n663), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n641), .A2(KEYINPUT102), .A3(new_n661), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT10), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n618), .B1(new_n614), .B2(KEYINPUT101), .ZN(new_n675));
  INV_X1    g474(.A(new_n646), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n572), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n578), .B1(new_n620), .B2(new_n615), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n649), .B1(new_n673), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n669), .B1(new_n657), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n656), .ZN(new_n683));
  INV_X1    g482(.A(new_n650), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n640), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n550), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n454), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g490(.A(KEYINPUT16), .B(G8gat), .Z(new_n692));
  NAND4_X1  g491(.A1(new_n550), .A2(new_n376), .A3(new_n687), .A4(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n550), .A2(new_n376), .A3(new_n687), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G8gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n693), .ZN(new_n696));
  MUX2_X1   g495(.A(new_n693), .B(new_n696), .S(KEYINPUT42), .Z(G1325gat));
  NAND3_X1  g496(.A1(new_n688), .A2(new_n504), .A3(new_n444), .ZN(new_n698));
  INV_X1    g497(.A(new_n466), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n688), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n700), .B2(new_n504), .ZN(G1326gat));
  NOR3_X1   g500(.A1(new_n477), .A2(new_n549), .A3(new_n235), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n687), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT43), .B(G22gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  INV_X1    g504(.A(new_n686), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n585), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n638), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n550), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n479), .A3(new_n689), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n446), .A2(new_n459), .A3(new_n410), .A4(new_n461), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n476), .A2(new_n470), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n638), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n707), .A2(new_n549), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n708), .A2(new_n718), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n719), .B(new_n720), .C1(new_n477), .C2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n454), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n710), .A2(KEYINPUT45), .A3(new_n479), .A4(new_n689), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n713), .A2(new_n724), .A3(new_n725), .ZN(G1328gat));
  NAND4_X1  g525(.A1(new_n550), .A2(new_n480), .A3(new_n376), .A4(new_n709), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT46), .Z(new_n728));
  OR3_X1    g527(.A1(new_n723), .A2(KEYINPUT106), .A3(new_n457), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT106), .B1(new_n723), .B2(new_n457), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(G36gat), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(G1329gat));
  NAND2_X1  g531(.A1(new_n699), .A2(G43gat), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n723), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n464), .A2(new_n467), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n715), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n736), .A2(new_n548), .A3(new_n444), .A4(new_n709), .ZN(new_n737));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(KEYINPUT47), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(KEYINPUT47), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n734), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n734), .B2(new_n740), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(G1330gat));
  OAI21_X1  g543(.A(G50gat), .B1(new_n723), .B2(new_n235), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n707), .A2(G50gat), .A3(new_n708), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n702), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1331gat));
  NOR3_X1   g550(.A1(new_n640), .A2(new_n548), .A3(new_n706), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n716), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n454), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n558), .ZN(G1332gat));
  XNOR2_X1  g554(.A(new_n457), .B(KEYINPUT109), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n753), .B2(new_n466), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n444), .A2(new_n552), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n753), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g564(.A1(new_n753), .A2(new_n235), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(new_n553), .ZN(G1335gat));
  INV_X1    g566(.A(new_n585), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n768), .A2(new_n548), .A3(new_n706), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n719), .B(new_n769), .C1(new_n477), .C2(new_n722), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n454), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n708), .B1(new_n714), .B2(new_n715), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n768), .A2(new_n548), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT51), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n454), .A2(G85gat), .A3(new_n706), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT110), .Z(new_n778));
  OAI21_X1  g577(.A(new_n771), .B1(new_n776), .B2(new_n778), .ZN(G1336gat));
  OAI21_X1  g578(.A(G92gat), .B1(new_n770), .B2(new_n457), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n756), .A2(G92gat), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n686), .B(new_n781), .C1(new_n774), .C2(new_n775), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n716), .A2(new_n638), .A3(new_n773), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n773), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n706), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(KEYINPUT111), .A3(new_n781), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n780), .A2(new_n784), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT52), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(new_n789), .B2(new_n781), .ZN(new_n793));
  OAI21_X1  g592(.A(G92gat), .B1(new_n770), .B2(new_n756), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT112), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n792), .A2(new_n797), .A3(new_n798), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n770), .B2(new_n466), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n789), .A2(new_n605), .A3(new_n444), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1338gat));
  OAI21_X1  g601(.A(G106gat), .B1(new_n770), .B2(new_n235), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n789), .A2(new_n606), .A3(new_n236), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n807), .A3(KEYINPUT53), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n803), .B(new_n804), .C1(new_n806), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(G1339gat));
  NAND3_X1  g610(.A1(new_n639), .A2(new_n549), .A3(new_n706), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n536), .A2(new_n537), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n521), .B1(new_n520), .B2(new_n528), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n543), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n547), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n686), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n673), .A2(new_n649), .A3(new_n679), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n667), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n822), .B(new_n659), .C1(new_n665), .C2(new_n666), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n823), .A2(KEYINPUT114), .A3(new_n683), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT114), .B1(new_n823), .B2(new_n683), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT55), .B(new_n821), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n548), .A3(new_n682), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n667), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829));
  AOI211_X1 g628(.A(KEYINPUT54), .B(new_n649), .C1(new_n673), .C2(new_n679), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n656), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n823), .A2(KEYINPUT114), .A3(new_n683), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(KEYINPUT55), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n819), .B1(new_n827), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n708), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n636), .A2(new_n637), .A3(new_n817), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n833), .B2(KEYINPUT55), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n826), .A2(new_n682), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n813), .B1(new_n842), .B2(new_n585), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n454), .ZN(new_n844));
  INV_X1    g643(.A(new_n469), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n756), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n548), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n840), .B1(new_n835), .B2(new_n708), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n812), .B1(new_n849), .B2(new_n768), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n235), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT115), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(new_n689), .A3(new_n444), .A4(new_n756), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n549), .A2(new_n246), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n848), .B1(new_n854), .B2(new_n855), .ZN(G1340gat));
  NAND3_X1  g655(.A1(new_n847), .A2(new_n244), .A3(new_n686), .ZN(new_n857));
  OAI21_X1  g656(.A(G120gat), .B1(new_n853), .B2(new_n706), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(KEYINPUT116), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(KEYINPUT116), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(G1341gat));
  NAND3_X1  g660(.A1(new_n847), .A2(new_n249), .A3(new_n768), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n854), .A2(new_n768), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(new_n249), .ZN(G1342gat));
  NAND2_X1  g664(.A1(new_n844), .A2(new_n845), .ZN(new_n866));
  NOR4_X1   g665(.A1(new_n866), .A2(G134gat), .A3(new_n376), .A4(new_n708), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n854), .A2(new_n638), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n870), .B2(new_n251), .ZN(G1343gat));
  NAND4_X1  g670(.A1(new_n844), .A2(new_n236), .A3(new_n466), .A4(new_n756), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(G141gat), .A3(new_n549), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n236), .A2(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n833), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n877), .B(new_n821), .C1(new_n824), .C2(new_n825), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT119), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n827), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT55), .B1(new_n883), .B2(KEYINPUT118), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n879), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n638), .B1(new_n887), .B2(new_n819), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n585), .B1(new_n888), .B2(new_n840), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n875), .B1(new_n889), .B2(new_n812), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n850), .A2(new_n236), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT117), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n894), .B(KEYINPUT57), .C1(new_n850), .C2(new_n236), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n890), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n466), .A2(new_n689), .A3(new_n756), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n896), .A2(new_n549), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(G141gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n874), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT120), .B1(new_n896), .B2(new_n897), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n891), .A2(KEYINPUT117), .A3(new_n892), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n876), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n903), .A2(new_n548), .A3(new_n682), .A4(new_n826), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n638), .B1(new_n904), .B2(new_n819), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n585), .B1(new_n905), .B2(new_n840), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n235), .B1(new_n906), .B2(new_n812), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n894), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n887), .A2(new_n819), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n708), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n841), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n813), .B1(new_n911), .B2(new_n585), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n902), .B(new_n908), .C1(new_n912), .C2(new_n875), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  INV_X1    g713(.A(new_n897), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n548), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n873), .B1(new_n917), .B2(G141gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n900), .B1(new_n918), .B2(new_n919), .ZN(G1344gat));
  NOR2_X1   g719(.A1(new_n872), .A2(new_n706), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n921), .A2(new_n922), .A3(G148gat), .ZN(new_n923));
  INV_X1    g722(.A(G148gat), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n843), .A2(new_n875), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT121), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n889), .A2(new_n812), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(new_n927), .B2(new_n236), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n686), .A3(new_n915), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n924), .B1(new_n930), .B2(KEYINPUT59), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n901), .A2(new_n916), .A3(new_n922), .A4(new_n686), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n923), .B1(new_n931), .B2(new_n932), .ZN(G1345gat));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n901), .A2(new_n768), .A3(new_n916), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G155gat), .ZN(new_n936));
  NOR4_X1   g735(.A1(new_n699), .A2(new_n843), .A3(new_n454), .A4(new_n235), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n937), .A2(new_n938), .A3(new_n768), .A4(new_n756), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT122), .B1(new_n872), .B2(new_n585), .ZN(new_n940));
  AOI21_X1  g739(.A(G155gat), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n934), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  AOI211_X1 g742(.A(KEYINPUT123), .B(new_n941), .C1(new_n935), .C2(G155gat), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(G1346gat));
  NAND4_X1  g744(.A1(new_n937), .A2(new_n213), .A3(new_n457), .A4(new_n638), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n901), .A2(new_n638), .A3(new_n916), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(new_n213), .ZN(G1347gat));
  NOR3_X1   g747(.A1(new_n843), .A2(new_n689), .A3(new_n756), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n845), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(G169gat), .B1(new_n951), .B2(new_n548), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n454), .A2(new_n376), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n953), .B1(new_n443), .B2(new_n442), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n852), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n549), .A2(new_n316), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(G1348gat));
  OAI21_X1  g757(.A(G176gat), .B1(new_n955), .B2(new_n706), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n951), .A2(new_n317), .A3(new_n686), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT124), .Z(G1349gat));
  OAI21_X1  g761(.A(G183gat), .B1(new_n955), .B2(new_n585), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n951), .A2(new_n343), .A3(new_n768), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n312), .A3(new_n638), .ZN(new_n967));
  OAI21_X1  g766(.A(G190gat), .B1(new_n955), .B2(new_n708), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  INV_X1    g770(.A(G197gat), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n699), .A2(new_n953), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n929), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n972), .B1(new_n974), .B2(new_n548), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n949), .A2(new_n236), .A3(new_n466), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(new_n972), .A3(new_n548), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT125), .Z(new_n978));
  OR2_X1    g777(.A1(new_n975), .A2(new_n978), .ZN(G1352gat));
  INV_X1    g778(.A(G204gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n976), .A2(new_n980), .A3(new_n686), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n981), .B(new_n982), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n686), .B(new_n973), .C1(new_n926), .C2(new_n928), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT126), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n983), .A2(new_n988), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(G1353gat));
  INV_X1    g789(.A(G211gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n991), .A3(new_n768), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n929), .A2(new_n768), .A3(new_n973), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n993), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n994));
  AOI21_X1  g793(.A(KEYINPUT63), .B1(new_n993), .B2(G211gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n976), .B2(new_n638), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT127), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n638), .A2(G218gat), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n998), .B1(new_n974), .B2(new_n999), .ZN(G1355gat));
endmodule


