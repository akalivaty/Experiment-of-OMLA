//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  AND2_X1   g0023(.A1(G87), .A2(G250), .ZN(new_n224));
  NOR4_X1   g0024(.A1(new_n219), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G107), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n202), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G238), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n203), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(new_n209), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n204), .A2(new_n205), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n236), .A2(new_n220), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n214), .B(new_n233), .C1(new_n235), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  INV_X1    g0047(.A(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT66), .B(G107), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT65), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G50), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  NAND3_X1  g0056(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n234), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(KEYINPUT69), .A3(new_n257), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n208), .A2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT69), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(new_n258), .B2(new_n261), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n259), .B1(new_n267), .B2(G50), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT70), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT8), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G58), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n273));
  MUX2_X1   g0073(.A(new_n272), .B(KEYINPUT68), .S(new_n273), .Z(new_n274));
  NAND2_X1  g0074(.A1(new_n209), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n209), .B1(new_n236), .B2(new_n220), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n261), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n269), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT67), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n283), .A2(KEYINPUT67), .A3(G1), .A4(G13), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G223), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G222), .B2(G1698), .ZN(new_n291));
  OR2_X1    g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n288), .B(new_n295), .C1(G77), .C2(new_n294), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n284), .A2(new_n297), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n296), .B(new_n300), .C1(new_n221), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n282), .B(new_n304), .C1(G179), .C2(new_n302), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n282), .B(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n302), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT72), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n311), .A2(new_n314), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n305), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n277), .A2(G50), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT75), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n275), .A2(new_n215), .B1(new_n209), .B2(G68), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n261), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g0121(.A(new_n321), .B(KEYINPUT11), .Z(new_n322));
  INV_X1    g0122(.A(new_n264), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n323), .A2(new_n261), .A3(new_n203), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n257), .A2(G68), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n292), .A2(new_n293), .B1(new_n226), .B2(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(G1698), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n221), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G33), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n217), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n330), .B(new_n288), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n288), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n337), .B1(new_n331), .B2(new_n333), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT73), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n301), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n299), .B1(new_n342), .B2(G238), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT13), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n338), .A2(new_n341), .A3(new_n346), .A4(new_n343), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n329), .B1(new_n348), .B2(G169), .ZN(new_n349));
  AOI211_X1 g0149(.A(KEYINPUT14), .B(new_n303), .C1(new_n345), .C2(new_n347), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n345), .A2(new_n353), .A3(new_n347), .ZN(new_n354));
  OR3_X1    g0154(.A1(new_n344), .A2(new_n353), .A3(KEYINPUT13), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n328), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(G200), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n354), .A2(new_n355), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n327), .B(new_n358), .C1(new_n359), .C2(new_n308), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n230), .A2(G1698), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G232), .B2(G1698), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n294), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n288), .B(new_n364), .C1(G107), .C2(new_n294), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n300), .C1(new_n216), .C2(new_n301), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n303), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n323), .A2(new_n261), .A3(new_n215), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G20), .A2(G77), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n271), .A2(new_n273), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n369), .B1(new_n370), .B2(new_n275), .C1(new_n371), .C2(new_n278), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n368), .B1(new_n372), .B2(new_n261), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G77), .B2(new_n257), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT71), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n366), .A2(G179), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT71), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n367), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n366), .A2(G200), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n308), .B2(new_n366), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(new_n374), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n204), .A2(new_n205), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n277), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT76), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n292), .A2(new_n209), .A3(new_n293), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  NOR2_X1   g0194(.A1(KEYINPUT3), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT7), .B1(new_n396), .B2(new_n209), .ZN(new_n397));
  OAI21_X1  g0197(.A(G68), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n387), .A2(new_n399), .A3(new_n388), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n391), .A2(new_n392), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n396), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n203), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n402), .B1(new_n405), .B2(new_n389), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(new_n261), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n267), .A2(new_n274), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n258), .B2(new_n274), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n289), .A2(new_n332), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n221), .A2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n394), .C2(new_n395), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G87), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT77), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT77), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n413), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n288), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n284), .A2(G232), .A3(new_n297), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT78), .B1(new_n300), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n300), .A2(new_n421), .A3(KEYINPUT78), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(G169), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n424), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n422), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(new_n419), .A3(G179), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n410), .A2(new_n430), .A3(KEYINPUT18), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT18), .B1(new_n410), .B2(new_n430), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G200), .B1(new_n420), .B2(new_n425), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n428), .A2(new_n419), .A3(G190), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n407), .A2(new_n434), .A3(new_n435), .A4(new_n409), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n317), .A2(new_n361), .A3(new_n384), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n216), .A2(G1698), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n440), .B1(G238), .B2(G1698), .C1(new_n394), .C2(new_n395), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n288), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT82), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n208), .A2(KEYINPUT82), .A3(G45), .A4(G274), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n208), .A2(G45), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n284), .A2(G250), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT83), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n444), .B(G179), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n441), .A2(new_n442), .B1(new_n286), .B2(new_n287), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n451), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT83), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n449), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n454), .B1(new_n460), .B2(new_n303), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n454), .B(KEYINPUT84), .C1(new_n460), .C2(new_n303), .ZN(new_n464));
  INV_X1    g0264(.A(new_n370), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n257), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G97), .A2(G107), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT85), .A2(G87), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT85), .A2(G87), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(KEYINPUT19), .C1(G20), .C2(new_n337), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n294), .A2(new_n209), .A3(G68), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT19), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n275), .B2(new_n217), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n466), .B1(new_n475), .B2(new_n261), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n208), .A2(G33), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n257), .A2(new_n477), .A3(new_n234), .A4(new_n260), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n370), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n463), .A2(new_n464), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n460), .A2(G190), .ZN(new_n481));
  INV_X1    g0281(.A(G87), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  AOI211_X1 g0283(.A(new_n483), .B(new_n466), .C1(new_n475), .C2(new_n261), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n444), .B1(new_n452), .B2(new_n453), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G200), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n478), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n258), .A2(new_n248), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n260), .A2(new_n234), .B1(G20), .B2(new_n248), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(new_n209), .C1(G33), .C2(new_n217), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n492), .A2(KEYINPUT20), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT20), .B1(new_n492), .B2(new_n494), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n490), .B(new_n491), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n294), .A2(G303), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G257), .A2(G1698), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n228), .A2(G1698), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n500), .A2(new_n501), .B1(new_n292), .B2(new_n293), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT87), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n332), .A2(G264), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n504), .A2(new_n499), .B1(new_n394), .B2(new_n395), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT87), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n506), .C1(G303), .C2(new_n294), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n288), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G41), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n208), .B(G45), .C1(new_n509), .C2(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT79), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G41), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT79), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n208), .A4(G45), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n298), .B1(KEYINPUT5), .B2(new_n509), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n511), .A2(new_n515), .A3(new_n284), .A4(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n512), .A2(G41), .ZN(new_n518));
  OAI211_X1 g0318(.A(G270), .B(new_n284), .C1(new_n510), .C2(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n517), .A2(KEYINPUT86), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT86), .B1(new_n517), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n508), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n497), .B1(new_n522), .B2(G200), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT88), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n508), .B(G190), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n522), .A2(G169), .A3(new_n497), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT21), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT21), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n522), .A2(new_n531), .A3(G169), .A4(new_n497), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n497), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n522), .A2(new_n534), .A3(new_n352), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G244), .B(new_n332), .C1(new_n394), .C2(new_n395), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n294), .A2(KEYINPUT4), .A3(G244), .A4(new_n332), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n294), .A2(G250), .A3(G1698), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n493), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n288), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(new_n284), .C1(new_n510), .C2(new_n518), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n517), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT80), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n517), .A2(new_n549), .A3(new_n546), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n545), .A2(new_n548), .A3(new_n352), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT81), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n517), .A2(new_n549), .A3(new_n546), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n549), .B1(new_n517), .B2(new_n546), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(KEYINPUT81), .A3(new_n352), .A4(new_n545), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n545), .A2(new_n548), .A3(new_n550), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n303), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n257), .A2(G97), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n478), .A2(new_n217), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n227), .B1(new_n403), .B2(new_n404), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n278), .A2(new_n215), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT6), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n217), .A2(new_n227), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n467), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n227), .A2(KEYINPUT6), .A3(G97), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n209), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n564), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n561), .B(new_n563), .C1(new_n571), .C2(new_n262), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n553), .A2(new_n557), .A3(new_n559), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n403), .A2(new_n404), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G107), .ZN(new_n575));
  INV_X1    g0375(.A(new_n565), .ZN(new_n576));
  INV_X1    g0376(.A(new_n570), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI211_X1 g0378(.A(new_n560), .B(new_n562), .C1(new_n578), .C2(new_n261), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n558), .A2(G200), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n556), .A2(G190), .A3(new_n545), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n573), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n528), .A2(new_n537), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G264), .B(new_n284), .C1(new_n510), .C2(new_n518), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G250), .A2(G1698), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n396), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n218), .A2(G1698), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n588), .B1(G33), .B2(G294), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n517), .B(new_n585), .C1(new_n589), .C2(new_n339), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n303), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(G179), .B2(new_n590), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT90), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT90), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT23), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n594), .A2(new_n596), .B1(G20), .B2(new_n227), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n593), .A2(KEYINPUT90), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n227), .A2(G20), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n209), .B(G87), .C1(new_n394), .C2(new_n395), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT22), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n275), .A2(new_n248), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n294), .A2(KEYINPUT22), .A3(new_n209), .A4(G87), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n601), .A2(new_n604), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT91), .ZN(new_n609));
  XNOR2_X1  g0409(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n611), .A2(new_n261), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n609), .ZN(new_n613));
  INV_X1    g0413(.A(new_n602), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n605), .B1(new_n614), .B2(KEYINPUT22), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n615), .A2(KEYINPUT91), .A3(new_n604), .A4(new_n601), .ZN(new_n616));
  INV_X1    g0416(.A(new_n610), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n612), .A2(new_n618), .B1(G107), .B2(new_n489), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n257), .A2(G107), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT25), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n592), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n489), .A2(G107), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n618), .A2(new_n261), .A3(new_n611), .ZN(new_n624));
  INV_X1    g0424(.A(G200), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n590), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n585), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n294), .B(new_n588), .C1(G250), .C2(G1698), .ZN(new_n628));
  NAND2_X1  g0428(.A1(G33), .A2(G294), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n630), .B2(new_n288), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n308), .A3(new_n517), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n623), .A2(new_n624), .A3(new_n621), .A4(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT92), .B1(new_n622), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n624), .A2(new_n623), .A3(new_n621), .ZN(new_n636));
  INV_X1    g0436(.A(new_n592), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n624), .A2(new_n623), .A3(new_n621), .A4(new_n633), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n439), .A2(new_n488), .A3(new_n584), .A4(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n380), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n360), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n356), .A2(new_n349), .A3(new_n350), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n327), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n437), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n433), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n316), .B2(new_n315), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n305), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n461), .A2(new_n479), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n487), .A2(new_n640), .A3(new_n573), .A4(new_n582), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n535), .B1(new_n530), .B2(new_n532), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n638), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n487), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n573), .A2(new_n658), .A3(KEYINPUT26), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n553), .A2(new_n557), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n559), .A2(new_n572), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n480), .A2(new_n660), .A3(new_n487), .A4(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n659), .B1(KEYINPUT26), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n439), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n651), .A2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G13), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G20), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .A3(G1), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT27), .B1(new_n669), .B2(G1), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n636), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n642), .A2(new_n675), .B1(new_n622), .B2(new_n674), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n497), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n655), .B(new_n677), .C1(new_n527), .C2(new_n526), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n655), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n674), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n642), .A2(new_n537), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n622), .A2(new_n683), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n212), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n468), .A2(new_n469), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n248), .A3(new_n467), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n689), .A2(new_n691), .A3(new_n208), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n237), .B2(new_n689), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT28), .Z(new_n694));
  AND2_X1   g0494(.A1(new_n638), .A2(new_n655), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n640), .A2(new_n573), .A3(new_n582), .A4(new_n487), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n652), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT26), .B1(new_n573), .B2(new_n658), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n683), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n642), .A2(new_n584), .A3(new_n488), .A4(new_n683), .ZN(new_n703));
  INV_X1    g0503(.A(new_n558), .ZN(new_n704));
  INV_X1    g0504(.A(new_n522), .ZN(new_n705));
  INV_X1    g0505(.A(new_n454), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .A4(new_n631), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n556), .A2(new_n545), .A3(new_n631), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n706), .A4(new_n705), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n522), .A2(new_n590), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n352), .A3(new_n485), .A4(new_n558), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT31), .B1(new_n714), .B2(new_n674), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n702), .B1(new_n703), .B2(new_n717), .ZN(new_n718));
  AOI211_X1 g0518(.A(KEYINPUT29), .B(new_n674), .C1(new_n657), .C2(new_n663), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n701), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n694), .B1(new_n720), .B2(G1), .ZN(G364));
  AOI21_X1  g0521(.A(new_n208), .B1(new_n668), .B2(G45), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n689), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(KEYINPUT93), .B(G169), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n234), .B1(new_n726), .B2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(G20), .A3(G179), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n729), .B1(G20), .B2(G179), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G190), .A2(G200), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n308), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n738), .A2(new_n215), .B1(new_n202), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT95), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n209), .A2(G179), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n625), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(G107), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n308), .A2(new_n625), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n743), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(new_n690), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n733), .A2(KEYINPUT96), .A3(new_n744), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT96), .B1(new_n733), .B2(new_n744), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT32), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n750), .A2(new_n736), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G159), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n756), .A2(new_n203), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n396), .B(new_n762), .C1(new_n757), .C2(new_n761), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n209), .B1(new_n739), .B2(new_n352), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n217), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n734), .A2(new_n749), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(G50), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n747), .A2(new_n753), .A3(new_n763), .A4(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT33), .B(G317), .Z(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n756), .A2(new_n769), .B1(new_n770), .B2(new_n745), .ZN(new_n771));
  INV_X1    g0571(.A(new_n764), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(G294), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n751), .A2(G303), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n737), .A2(G311), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n766), .A2(G326), .B1(G329), .B2(new_n758), .ZN(new_n776));
  INV_X1    g0576(.A(new_n740), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n294), .B1(new_n777), .B2(G322), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n728), .B1(new_n768), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n727), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n255), .A2(G45), .ZN(new_n786));
  INV_X1    g0586(.A(G45), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n237), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n688), .A2(new_n294), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n212), .A2(G355), .A3(new_n294), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n791), .C1(G116), .C2(new_n212), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n725), .B(new_n781), .C1(new_n785), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n784), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n679), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n724), .B1(new_n679), .B2(G330), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G330), .B2(new_n679), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  NAND2_X1  g0599(.A1(new_n374), .A2(new_n674), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n380), .A2(new_n383), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n380), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n662), .A2(KEYINPUT26), .ZN(new_n803));
  INV_X1    g0603(.A(new_n659), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n683), .B(new_n802), .C1(new_n697), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT98), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n674), .B1(new_n657), .B2(new_n663), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n809), .A2(KEYINPUT98), .A3(new_n802), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n809), .B2(new_n802), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(new_n718), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n725), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G159), .A2(new_n737), .B1(new_n777), .B2(G143), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  INV_X1    g0616(.A(new_n766), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n817), .C1(new_n276), .C2(new_n756), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT34), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n751), .A2(G50), .B1(new_n746), .B2(G68), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n202), .B2(new_n764), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n396), .B(new_n821), .C1(G132), .C2(new_n758), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n738), .A2(new_n248), .B1(new_n824), .B2(new_n740), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G303), .B2(new_n766), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n294), .B1(new_n746), .B2(G87), .ZN(new_n827));
  INV_X1    g0627(.A(new_n756), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G283), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n759), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n765), .B(new_n831), .C1(G107), .C2(new_n751), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n826), .A2(new_n827), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n728), .B1(new_n823), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n727), .A2(new_n782), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n725), .B(new_n834), .C1(new_n215), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT97), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n783), .B2(new_n802), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n814), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  OAI21_X1  g0640(.A(new_n439), .B1(new_n701), .B2(new_n719), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n651), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n703), .A2(new_n717), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n439), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT107), .Z(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  INV_X1    g0647(.A(new_n672), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n410), .B1(new_n430), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n850), .A3(new_n436), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n401), .A2(new_n261), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n277), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n574), .A2(G68), .B1(new_n854), .B2(new_n399), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT16), .B1(new_n855), .B2(new_n390), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n409), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n848), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT101), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(KEYINPUT101), .A3(new_n848), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n857), .A2(new_n430), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n860), .A2(new_n436), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n852), .B1(new_n863), .B2(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n398), .A2(new_n400), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n854), .A2(new_n399), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n402), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(new_n261), .A3(new_n401), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n859), .B(new_n672), .C1(new_n868), .C2(new_n409), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT101), .B1(new_n857), .B2(new_n848), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n433), .B2(new_n437), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n847), .B1(new_n864), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n860), .A2(new_n861), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT17), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n436), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n431), .A2(new_n432), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n862), .A2(new_n436), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n850), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n878), .B(KEYINPUT38), .C1(new_n880), .C2(new_n852), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT100), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n328), .A2(new_n884), .A3(new_n674), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n360), .B(new_n885), .C1(new_n646), .C2(new_n327), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n328), .B2(new_n674), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n886), .A2(new_n887), .B1(new_n357), .B2(new_n683), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n844), .A2(new_n888), .A3(new_n802), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(KEYINPUT40), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n410), .B(new_n848), .C1(new_n876), .C2(new_n877), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n850), .B1(new_n849), .B2(new_n436), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT102), .B1(new_n852), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n849), .A2(new_n436), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(new_n851), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n894), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n847), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n851), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(KEYINPUT103), .A3(KEYINPUT38), .A4(new_n878), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n893), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT105), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT105), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n893), .A2(new_n902), .A3(new_n905), .A4(new_n908), .ZN(new_n909));
  AND4_X1   g0709(.A1(KEYINPUT40), .A2(new_n844), .A3(new_n888), .A4(new_n802), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT106), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT106), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n907), .A2(new_n913), .A3(new_n909), .A4(new_n910), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n891), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n846), .B(new_n915), .Z(new_n916));
  OAI21_X1  g0716(.A(new_n843), .B1(new_n916), .B2(new_n702), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n433), .A2(new_n848), .ZN(new_n919));
  INV_X1    g0719(.A(new_n888), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n380), .A2(new_n674), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n920), .B1(new_n811), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n919), .B1(new_n923), .B2(new_n882), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n906), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n357), .A2(new_n674), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT104), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(KEYINPUT104), .A3(new_n929), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n916), .A2(new_n702), .A3(new_n843), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n918), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n933), .B1(new_n918), .B2(new_n934), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n208), .C2(new_n668), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n568), .A2(new_n569), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n248), .B1(new_n938), .B2(KEYINPUT35), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n939), .B(new_n235), .C1(KEYINPUT35), .C2(new_n938), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT36), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n237), .A2(G77), .A3(new_n385), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(G50), .B2(new_n203), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n667), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT99), .Z(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(new_n941), .A3(new_n945), .ZN(G367));
  NOR2_X1   g0746(.A1(new_n579), .A2(new_n683), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n583), .A2(new_n947), .B1(new_n573), .B2(new_n683), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT108), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n684), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT42), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n573), .B1(new_n949), .B2(new_n638), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n683), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n484), .A2(new_n683), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(new_n652), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n652), .A3(new_n487), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n951), .A2(new_n953), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n949), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n681), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n960), .B(new_n962), .Z(new_n963));
  XNOR2_X1  g0763(.A(new_n689), .B(KEYINPUT41), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n686), .A2(new_n961), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT45), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n686), .A2(new_n961), .ZN(new_n969));
  XNOR2_X1  g0769(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n966), .B1(new_n972), .B2(new_n681), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n968), .A2(KEYINPUT110), .A3(new_n971), .A4(new_n682), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n676), .B1(new_n655), .B2(new_n674), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n684), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n681), .B1(new_n977), .B2(new_n680), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n978), .A2(new_n720), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n965), .B1(new_n980), .B2(new_n720), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n963), .B1(new_n981), .B2(new_n723), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n957), .A2(new_n794), .ZN(new_n983));
  INV_X1    g0783(.A(new_n245), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n784), .B(new_n727), .C1(new_n984), .C2(new_n789), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n688), .A2(new_n465), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n724), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n752), .A2(new_n248), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n828), .A2(G294), .B1(KEYINPUT46), .B2(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(KEYINPUT46), .B2(new_n989), .C1(new_n830), .C2(new_n817), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n777), .A2(G303), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n764), .A2(new_n227), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n738), .A2(new_n770), .ZN(new_n994));
  NOR4_X1   g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n746), .A2(G97), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n758), .A2(G317), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n995), .A2(new_n396), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n756), .A2(new_n760), .B1(new_n738), .B2(new_n220), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT111), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n999), .A2(new_n1000), .B1(G150), .B2(new_n777), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n294), .B1(new_n745), .B2(new_n215), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1001), .B1(KEYINPUT112), .B2(new_n1002), .C1(new_n203), .C2(new_n764), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G143), .B2(new_n766), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1002), .A2(KEYINPUT112), .B1(new_n751), .B2(G58), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n816), .C2(new_n759), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n999), .A2(new_n1000), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n998), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n983), .B(new_n988), .C1(new_n1009), .C2(new_n727), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n982), .A2(new_n1011), .ZN(G387));
  NAND2_X1  g0812(.A1(new_n676), .A2(new_n784), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n371), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n220), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT50), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n203), .A2(new_n215), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1016), .A2(G45), .A3(new_n1017), .A4(new_n691), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n691), .A2(new_n212), .A3(new_n294), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n789), .B1(new_n242), .B2(new_n787), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n212), .A2(G107), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n785), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1013), .A2(new_n724), .A3(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G303), .A2(new_n737), .B1(new_n777), .B2(G317), .ZN(new_n1025));
  INV_X1    g0825(.A(G322), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1025), .B1(new_n1026), .B2(new_n817), .C1(new_n830), .C2(new_n756), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n770), .B2(new_n764), .C1(new_n824), .C2(new_n752), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n294), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n758), .A2(G326), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n746), .A2(G116), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n756), .A2(new_n274), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n996), .B1(new_n752), .B2(new_n215), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1036), .A2(new_n396), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n276), .B2(new_n759), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G68), .B2(new_n737), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n772), .A2(new_n465), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n220), .C2(new_n740), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n766), .A2(G159), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT113), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1035), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1024), .B1(new_n1045), .B2(new_n727), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n723), .B2(new_n978), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n689), .B1(new_n978), .B2(new_n720), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n979), .ZN(G393));
  AOI22_X1  g0849(.A1(new_n973), .A2(new_n974), .B1(new_n681), .B2(new_n972), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n980), .B(new_n689), .C1(new_n979), .C2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n396), .B1(new_n745), .B2(new_n227), .C1(new_n764), .C2(new_n248), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G317), .A2(new_n766), .B1(new_n777), .B2(G311), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT52), .Z(new_n1054));
  AOI22_X1  g0854(.A1(new_n737), .A2(G294), .B1(G283), .B2(new_n751), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n1026), .C2(new_n759), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1052), .B(new_n1056), .C1(G303), .C2(new_n828), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G150), .A2(new_n766), .B1(new_n777), .B2(G159), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n294), .B1(new_n215), .B2(new_n764), .C1(new_n1058), .C2(KEYINPUT51), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n828), .A2(G50), .B1(G68), .B2(new_n751), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G143), .A2(new_n758), .B1(new_n746), .B2(G87), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1059), .B(new_n1063), .C1(new_n1014), .C2(new_n737), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(new_n728), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n724), .B1(new_n961), .B2(new_n794), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n251), .A2(new_n789), .B1(G97), .B2(new_n688), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1066), .B(new_n1067), .C1(new_n785), .C2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1050), .B2(new_n723), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1051), .A2(new_n1070), .ZN(G390));
  NAND2_X1  g0871(.A1(new_n926), .A2(new_n927), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n928), .B2(new_n923), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n802), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n922), .B1(new_n700), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n928), .B1(new_n1075), .B2(new_n888), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n907), .A2(new_n909), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n718), .A2(new_n802), .A3(new_n888), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT114), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1073), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(KEYINPUT115), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n718), .A2(new_n802), .A3(new_n888), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT115), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1073), .A2(new_n1085), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1081), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n722), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1072), .A2(new_n782), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G128), .A2(new_n766), .B1(new_n777), .B2(G132), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT53), .B1(new_n752), .B2(new_n276), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G125), .A2(new_n758), .B1(new_n746), .B2(G50), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1090), .A2(new_n294), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  OR3_X1    g0893(.A1(new_n752), .A2(KEYINPUT53), .A3(new_n276), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n760), .B2(new_n764), .C1(new_n756), .C2(new_n816), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT54), .B(G143), .Z(new_n1096));
  AOI211_X1 g0896(.A(new_n1093), .B(new_n1095), .C1(new_n737), .C2(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n396), .B1(new_n203), .B2(new_n745), .C1(new_n752), .C2(new_n482), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n828), .A2(G107), .B1(G294), .B2(new_n758), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n215), .B2(new_n764), .C1(new_n248), .C2(new_n740), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(G283), .C2(new_n766), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n737), .A2(G97), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1097), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT118), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n727), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1089), .A2(new_n724), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n274), .B2(new_n835), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1088), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n841), .B(new_n651), .C1(new_n702), .C2(new_n845), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n806), .A2(new_n807), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT98), .B1(new_n809), .B2(new_n802), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n922), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n888), .B1(new_n718), .B2(new_n802), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n1083), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT116), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1112), .B(new_n1116), .C1(new_n1083), .C2(new_n1113), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1075), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1113), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1079), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1109), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1087), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1122), .A2(new_n1081), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n689), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1108), .B1(new_n1128), .B2(new_n1129), .ZN(G378));
  XNOR2_X1  g0930(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT121), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT55), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n317), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n282), .A2(new_n848), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1133), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n782), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n740), .A2(new_n227), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n828), .A2(G97), .B1(G58), .B2(new_n746), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n203), .B2(new_n764), .C1(new_n370), .C2(new_n738), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1145), .B(new_n1147), .C1(G116), .C2(new_n766), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n509), .B(new_n396), .C1(new_n752), .C2(new_n215), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT119), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(new_n770), .C2(new_n759), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT58), .Z(new_n1152));
  OAI21_X1  g0952(.A(new_n220), .B1(new_n394), .B2(G41), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n828), .A2(G132), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n777), .A2(G128), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G125), .A2(new_n766), .B1(new_n737), .B2(G137), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n772), .A2(G150), .B1(new_n751), .B2(new_n1096), .ZN(new_n1157));
  AND4_X1   g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT59), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G33), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G41), .B1(new_n758), .B2(G124), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n760), .C2(new_n745), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1153), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n727), .B1(new_n1152), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n835), .A2(new_n220), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1144), .A2(new_n724), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n912), .A2(new_n914), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n891), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(G330), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n931), .A3(new_n932), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n924), .A2(KEYINPUT104), .A3(new_n929), .ZN(new_n1172));
  OAI211_X1 g0972(.A(G330), .B(new_n915), .C1(new_n1172), .C2(new_n930), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1142), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n1173), .A3(new_n1143), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1167), .B1(new_n1177), .B2(new_n722), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n689), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1109), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1125), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(new_n1176), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1175), .A2(KEYINPUT57), .A3(new_n1176), .A4(new_n1181), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1178), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  NAND3_X1  g0987(.A1(new_n1118), .A2(new_n1109), .A3(new_n1121), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1123), .A2(new_n964), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n722), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n920), .A2(new_n782), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n828), .A2(G116), .B1(G303), .B2(new_n758), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1041), .C1(new_n770), .C2(new_n740), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n294), .B(new_n1193), .C1(G107), .C2(new_n737), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n751), .A2(G97), .B1(new_n746), .B2(G77), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n824), .C2(new_n817), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT122), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n738), .A2(new_n276), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n828), .A2(new_n1096), .B1(G50), .B2(new_n772), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n758), .A2(G128), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n816), .C2(new_n740), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(G159), .C2(new_n751), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n766), .A2(G132), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n294), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G58), .B2(new_n746), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n727), .B1(new_n1197), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n835), .A2(new_n203), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n724), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT123), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1190), .B1(new_n1191), .B2(new_n1209), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1189), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(G381));
  NAND2_X1  g1012(.A1(new_n1108), .A2(new_n1126), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G375), .A2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n982), .A2(new_n1011), .A3(new_n1070), .A4(new_n1051), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1215), .A2(G396), .A3(G393), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n839), .A3(new_n1211), .A4(new_n1216), .ZN(G407));
  INV_X1    g1017(.A(G213), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1214), .B2(new_n673), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(G407), .ZN(G409));
  XNOR2_X1  g1020(.A(G393), .B(new_n798), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(G387), .A2(G390), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(KEYINPUT127), .A3(new_n1215), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT127), .B1(new_n1223), .B2(new_n1215), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1222), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1222), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1188), .B1(new_n1122), .B2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1118), .A2(new_n1121), .A3(KEYINPUT60), .A4(new_n1109), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n689), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT124), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1232), .A2(new_n1236), .A3(new_n689), .A4(new_n1233), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1210), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n839), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(G384), .A3(new_n1210), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1218), .A2(G343), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT126), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(G2897), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1240), .A2(new_n1241), .A3(new_n1246), .A4(new_n1244), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1167), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1171), .A2(new_n1143), .A3(new_n1173), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1143), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1250), .B1(new_n1253), .B2(new_n723), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n964), .A3(new_n1181), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1213), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1186), .B2(G378), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1248), .B(new_n1249), .C1(new_n1257), .C2(new_n1242), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n689), .A3(new_n1185), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(G378), .A3(new_n1254), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1182), .A2(new_n965), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1108), .B(new_n1126), .C1(new_n1178), .C2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1243), .A4(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1258), .A2(new_n1259), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1242), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1266), .B1(new_n1271), .B2(new_n1268), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1230), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1257), .A2(new_n1242), .A3(new_n1267), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(KEYINPUT63), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1271), .A2(new_n1268), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(KEYINPUT125), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1227), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1271), .A2(KEYINPUT63), .A3(new_n1268), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1259), .A3(new_n1258), .A4(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1273), .B1(new_n1280), .B2(new_n1283), .ZN(G405));
  OAI21_X1  g1084(.A(new_n1262), .B1(new_n1186), .B2(new_n1213), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1267), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1281), .ZN(G402));
endmodule


