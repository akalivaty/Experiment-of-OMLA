//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT77), .Z(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT69), .B(KEYINPUT26), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n205), .B1(new_n209), .B2(KEYINPUT70), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT26), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n210), .B(new_n212), .C1(KEYINPUT70), .C2(new_n209), .ZN(new_n213));
  XOR2_X1   g012(.A(KEYINPUT27), .B(G183gat), .Z(new_n214));
  OAI21_X1  g013(.A(KEYINPUT28), .B1(new_n214), .B2(G190gat), .ZN(new_n215));
  AOI21_X1  g014(.A(G190gat), .B1(new_n214), .B2(KEYINPUT68), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT68), .B1(new_n217), .B2(KEYINPUT27), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT28), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n216), .A2(new_n219), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n213), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT23), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n225), .A3(new_n204), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(KEYINPUT24), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n223), .A2(new_n225), .A3(new_n235), .A4(new_n204), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n227), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n211), .B2(new_n224), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n223), .A2(new_n241), .A3(new_n204), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n223), .B2(new_n204), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n234), .B(new_n240), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n230), .A2(G183gat), .A3(G190gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n228), .A2(KEYINPUT24), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n232), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n224), .A2(G169gat), .A3(G176gat), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT65), .B1(new_n250), .B2(new_n205), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n223), .A2(new_n241), .A3(new_n204), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT66), .B1(new_n253), .B2(new_n240), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n239), .B1(new_n246), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n244), .A2(new_n245), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(KEYINPUT66), .A3(new_n240), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(new_n239), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n222), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n203), .B1(new_n262), .B2(KEYINPUT29), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT78), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G211gat), .B(G218gat), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G197gat), .B(G204gat), .Z(new_n268));
  AOI21_X1  g067(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n270), .A2(KEYINPUT76), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n268), .A2(new_n269), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n266), .B1(new_n272), .B2(KEYINPUT76), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n255), .A2(new_n221), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n275), .A2(new_n203), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT78), .B(new_n203), .C1(new_n262), .C2(KEYINPUT29), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n265), .A2(new_n274), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n203), .B1(new_n275), .B2(KEYINPUT29), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n262), .B2(new_n203), .ZN(new_n280));
  INV_X1    g079(.A(new_n274), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G8gat), .B(G36gat), .ZN(new_n284));
  INV_X1    g083(.A(G92gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT79), .B(G64gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(KEYINPUT30), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n278), .A2(new_n282), .A3(new_n288), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(KEYINPUT80), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT30), .B1(new_n283), .B2(new_n289), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G134gat), .ZN(new_n299));
  INV_X1    g098(.A(G120gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G113gat), .ZN(new_n301));
  INV_X1    g100(.A(G113gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G120gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT71), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT1), .ZN(new_n305));
  INV_X1    g104(.A(G127gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n304), .B2(new_n305), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n299), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n302), .A2(G120gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n300), .A2(G113gat), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n311), .B(new_n305), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G127gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(new_n307), .A3(G134gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G141gat), .B(G148gat), .Z(new_n318));
  XOR2_X1   g117(.A(KEYINPUT81), .B(KEYINPUT2), .Z(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(new_n319), .B1(G155gat), .B2(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G141gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT82), .B(G141gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(new_n324), .ZN(new_n327));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(new_n323), .B2(KEYINPUT2), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n320), .A2(new_n323), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n318), .A2(new_n319), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(new_n328), .A3(new_n323), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n327), .A2(new_n329), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n317), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n310), .A2(new_n330), .A3(new_n316), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n315), .A2(G134gat), .A3(new_n307), .ZN(new_n341));
  AOI21_X1  g140(.A(G134gat), .B1(new_n315), .B2(new_n307), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n341), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n298), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n296), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n330), .B1(new_n310), .B2(new_n316), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT84), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT5), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n336), .B1(new_n341), .B2(new_n342), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n296), .B1(new_n352), .B2(new_n339), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT84), .B1(new_n353), .B2(new_n297), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n344), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n310), .A2(new_n330), .A3(KEYINPUT4), .A4(new_n316), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n338), .A2(new_n356), .A3(new_n296), .A4(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n346), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT87), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n367));
  INV_X1    g166(.A(new_n358), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n351), .B2(new_n354), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n364), .C1(new_n369), .C2(new_n346), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n350), .B1(new_n349), .B2(KEYINPUT5), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n353), .A2(KEYINPUT84), .A3(new_n297), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n358), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n346), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n365), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(KEYINPUT86), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT86), .B1(new_n376), .B2(new_n377), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n371), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT6), .B(new_n364), .C1(new_n369), .C2(new_n346), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n371), .B(KEYINPUT88), .C1(new_n378), .C2(new_n379), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n290), .A2(new_n291), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n295), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G78gat), .B(G106gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G22gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n332), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n274), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n272), .A2(new_n266), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n397), .A2(new_n270), .A3(new_n394), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n336), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT3), .B1(new_n281), .B2(new_n394), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n393), .B(new_n396), .C1(new_n405), .C2(new_n330), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n402), .B2(new_n406), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n392), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n409), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(new_n391), .A3(new_n407), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI221_X4 g212(.A(KEYINPUT67), .B1(new_n237), .B2(new_n238), .C1(new_n257), .C2(new_n258), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n260), .B1(new_n259), .B2(new_n239), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n221), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n317), .ZN(new_n417));
  NAND2_X1  g216(.A1(G227gat), .A2(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n317), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n419), .B(new_n221), .C1(new_n414), .C2(new_n415), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT73), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT34), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n421), .B2(KEYINPUT34), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT34), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n417), .A2(new_n427), .A3(new_n418), .A4(new_n420), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT74), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(G71gat), .B(G99gat), .Z(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT72), .ZN(new_n432));
  XNOR2_X1  g231(.A(G15gat), .B(G43gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n418), .B1(new_n417), .B2(new_n420), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n434), .B1(new_n435), .B2(KEYINPUT33), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n420), .ZN(new_n440));
  INV_X1    g239(.A(new_n418), .ZN(new_n441));
  AOI221_X4 g240(.A(new_n437), .B1(KEYINPUT33), .B2(new_n434), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  OAI22_X1  g241(.A1(new_n426), .A2(new_n430), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n441), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT32), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n447), .A3(new_n434), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n421), .A2(KEYINPUT34), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT73), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n423), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n438), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n428), .B(KEYINPUT74), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n448), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n413), .A2(new_n443), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT35), .B1(new_n389), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT6), .B1(new_n359), .B2(new_n365), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n359), .A2(new_n365), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NOR4_X1   g259(.A1(new_n386), .A2(new_n460), .A3(new_n293), .A4(KEYINPUT35), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n454), .A3(KEYINPUT75), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT75), .ZN(new_n463));
  OAI221_X1 g262(.A(new_n463), .B1(new_n439), .B2(new_n442), .C1(new_n426), .C2(new_n430), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n413), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n413), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n389), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n340), .A2(new_n347), .A3(new_n345), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n470), .A2(KEYINPUT90), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(KEYINPUT90), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n352), .A2(new_n339), .A3(new_n296), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT39), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT91), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n474), .A2(KEYINPUT91), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n471), .A2(new_n472), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n471), .A2(new_n472), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n365), .B(new_n477), .C1(new_n478), .C2(KEYINPUT39), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n459), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n481), .B(new_n482), .C1(new_n386), .C2(new_n293), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n280), .A2(new_n281), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n265), .A2(new_n276), .A3(new_n277), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT37), .B(new_n484), .C1(new_n485), .C2(new_n274), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n283), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT38), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n486), .A2(new_n488), .A3(new_n489), .A4(new_n288), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n283), .A2(new_n289), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n460), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n289), .B1(new_n283), .B2(new_n487), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n278), .A2(KEYINPUT37), .A3(new_n282), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n483), .B(new_n413), .C1(new_n492), .C2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n443), .B2(new_n454), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n465), .B2(new_n497), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n469), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n467), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G8gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(G1gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n504), .B2(KEYINPUT94), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT16), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n503), .B1(new_n506), .B2(G1gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(G1gat), .B2(new_n503), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n505), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G71gat), .B(G78gat), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(KEYINPUT97), .ZN(new_n512));
  XOR2_X1   g311(.A(G57gat), .B(G64gat), .Z(new_n513));
  INV_X1    g312(.A(KEYINPUT9), .ZN(new_n514));
  INV_X1    g313(.A(G71gat), .ZN(new_n515));
  INV_X1    g314(.A(G78gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n511), .A2(KEYINPUT97), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n512), .A2(new_n513), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(KEYINPUT9), .ZN(new_n520));
  INV_X1    g319(.A(new_n511), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT21), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G127gat), .B(G155gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT20), .Z(new_n530));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n526), .A3(new_n523), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n528), .B2(new_n531), .ZN(new_n533));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(G211gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  OR3_X1    g335(.A1(new_n532), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT99), .B(G183gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n536), .B1(new_n532), .B2(new_n533), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n540), .B1(new_n537), .B2(new_n541), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT102), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  AOI22_X1  g351(.A1(KEYINPUT8), .A2(new_n551), .B1(new_n552), .B2(new_n285), .ZN(new_n553));
  NAND2_X1  g352(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n552), .B2(new_n285), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n551), .ZN(new_n558));
  OR2_X1    g357(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n559));
  NAND3_X1  g358(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n560), .A2(new_n554), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n556), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n561), .A2(new_n553), .A3(new_n559), .A4(new_n555), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n551), .A3(new_n557), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n566));
  INV_X1    g365(.A(G29gat), .ZN(new_n567));
  INV_X1    g366(.A(G36gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(KEYINPUT92), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n571), .A2(KEYINPUT93), .A3(new_n572), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(G29gat), .A2(G36gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G50gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G43gat), .ZN(new_n581));
  INV_X1    g380(.A(G43gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(G50gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n583), .A3(KEYINPUT15), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n572), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n584), .A3(new_n578), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT15), .B1(new_n581), .B2(new_n583), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n565), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT17), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n586), .A2(new_n594), .A3(new_n591), .ZN(new_n595));
  INV_X1    g394(.A(new_n578), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n574), .B2(new_n575), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n584), .B1(new_n597), .B2(new_n577), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT17), .B1(new_n598), .B2(new_n590), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  AOI211_X1 g399(.A(new_n592), .B(new_n593), .C1(new_n600), .C2(new_n565), .ZN(new_n601));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n550), .B(new_n603), .C1(new_n605), .C2(new_n549), .ZN(new_n606));
  INV_X1    g405(.A(new_n603), .ZN(new_n607));
  OAI211_X1 g406(.A(KEYINPUT102), .B(new_n549), .C1(new_n607), .C2(new_n604), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n545), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n501), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n586), .A2(new_n591), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n509), .ZN(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n600), .B2(new_n510), .ZN(new_n618));
  AOI211_X1 g417(.A(KEYINPUT95), .B(new_n509), .C1(new_n595), .C2(new_n599), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT18), .B(new_n616), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n594), .B1(new_n586), .B2(new_n591), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n598), .A2(KEYINPUT17), .A3(new_n590), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n510), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT95), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n600), .A2(new_n617), .A3(new_n510), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n628), .A2(KEYINPUT96), .A3(KEYINPUT18), .A4(new_n616), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G113gat), .B(G141gat), .ZN(new_n631));
  INV_X1    g430(.A(G197gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT11), .B(G169gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  OAI21_X1  g435(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n612), .B(new_n509), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n614), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n630), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n636), .B1(new_n630), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n565), .A2(new_n523), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n519), .A2(new_n562), .A3(new_n564), .A4(new_n522), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n565), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n524), .A3(KEYINPUT10), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n646), .A2(new_n648), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n654), .B1(new_n655), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n656), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n611), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n385), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(G1gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1324gat));
  NOR2_X1   g464(.A1(new_n386), .A2(new_n293), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n502), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT104), .Z(new_n669));
  NAND2_X1  g468(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n506), .A2(new_n502), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT42), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(new_n662), .ZN(new_n675));
  INV_X1    g474(.A(new_n499), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n675), .A2(G15gat), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(G15gat), .B1(new_n675), .B2(new_n465), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(G1326gat));
  NOR2_X1   g478(.A1(new_n662), .A2(new_n413), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  AND2_X1   g481(.A1(new_n499), .A2(new_n496), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n683), .A2(new_n469), .B1(new_n457), .B2(new_n466), .ZN(new_n684));
  INV_X1    g483(.A(new_n609), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n684), .A2(new_n544), .A3(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(new_n661), .ZN(new_n687));
  INV_X1    g486(.A(new_n385), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n567), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT44), .B1(new_n501), .B2(new_n609), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n692), .B(new_n685), .C1(new_n467), .C2(new_n500), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n661), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n544), .B(KEYINPUT105), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n385), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n690), .A2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(new_n666), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n687), .A2(new_n568), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT46), .Z(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n701), .B2(new_n666), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n687), .A2(new_n582), .A3(new_n465), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n692), .B1(new_n684), .B2(new_n685), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n501), .A2(KEYINPUT44), .A3(new_n609), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n711), .A2(new_n676), .A3(new_n712), .A4(new_n698), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G43gat), .B1(new_n713), .B2(new_n714), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n710), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(G43gat), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n710), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n709), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n694), .A2(KEYINPUT106), .A3(new_n676), .A4(new_n698), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n715), .A3(G43gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n720), .B1(new_n726), .B2(new_n710), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(KEYINPUT107), .A3(new_n722), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n724), .A2(new_n728), .ZN(G1330gat));
  NAND2_X1  g528(.A1(new_n700), .A2(new_n468), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n413), .A2(G50gat), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(G50gat), .B1(new_n687), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g532(.A(new_n645), .ZN(new_n734));
  INV_X1    g533(.A(new_n660), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n611), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n688), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(G57gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n704), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT49), .B(G64gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1333gat));
  NAND3_X1  g543(.A1(new_n737), .A2(new_n515), .A3(new_n465), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n737), .A2(new_n676), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n515), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g547(.A1(new_n737), .A2(new_n468), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g549(.A1(new_n694), .A2(new_n545), .A3(new_n736), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(new_n552), .A3(new_n385), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n686), .A2(new_n645), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n753), .A2(KEYINPUT51), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(KEYINPUT51), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(new_n660), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n688), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n752), .B1(new_n757), .B2(new_n552), .ZN(G1336gat));
  OAI21_X1  g557(.A(G92gat), .B1(new_n751), .B2(new_n666), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n754), .A2(new_n660), .A3(new_n755), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n704), .A2(new_n285), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT52), .ZN(G1337gat));
  XOR2_X1   g562(.A(KEYINPUT109), .B(G99gat), .Z(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n751), .B2(new_n499), .ZN(new_n765));
  INV_X1    g564(.A(new_n465), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n766), .A2(new_n764), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n760), .B2(new_n767), .ZN(G1338gat));
  INV_X1    g567(.A(G106gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n756), .A2(new_n769), .A3(new_n468), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  OAI21_X1  g571(.A(G106gat), .B1(new_n751), .B2(new_n413), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n760), .A2(G106gat), .A3(new_n413), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n771), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT53), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(G1339gat));
  NAND3_X1  g577(.A1(new_n610), .A2(new_n645), .A3(new_n735), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n615), .B1(new_n626), .B2(new_n627), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT96), .B1(new_n780), .B2(KEYINPUT18), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n620), .A2(new_n621), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n636), .B(new_n642), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n649), .A2(new_n651), .A3(G230gat), .A4(G233gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n786));
  NAND3_X1  g585(.A1(new_n652), .A2(new_n653), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n659), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n788), .A2(new_n789), .B1(new_n656), .B2(new_n659), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n788), .A2(KEYINPUT112), .A3(new_n789), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n635), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n614), .B1(new_n628), .B2(new_n613), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n639), .A2(new_n641), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND4_X1   g598(.A1(new_n783), .A2(new_n795), .A3(new_n609), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n660), .A3(new_n799), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT113), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n795), .B1(new_n643), .B2(new_n644), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n783), .A2(new_n804), .A3(new_n660), .A4(new_n799), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n800), .B1(new_n806), .B2(new_n685), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n779), .B1(new_n807), .B2(new_n697), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n779), .B(new_n810), .C1(new_n807), .C2(new_n697), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n812), .A2(new_n385), .A3(new_n456), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n666), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n302), .A3(new_n734), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n812), .A2(new_n468), .A3(new_n766), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n688), .A3(new_n666), .ZN(new_n817));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n645), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(G1340gat));
  NAND3_X1  g618(.A1(new_n814), .A2(new_n300), .A3(new_n660), .ZN(new_n820));
  OAI21_X1  g619(.A(G120gat), .B1(new_n817), .B2(new_n735), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1341gat));
  INV_X1    g621(.A(new_n697), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n817), .A2(new_n306), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n814), .A2(new_n544), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT115), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n824), .B1(new_n826), .B2(new_n306), .ZN(G1342gat));
  NAND2_X1  g626(.A1(new_n666), .A2(new_n609), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT116), .Z(new_n829));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n299), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT56), .Z(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n817), .B2(new_n685), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1343gat));
  INV_X1    g632(.A(new_n779), .ZN(new_n834));
  INV_X1    g633(.A(new_n790), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n791), .C1(new_n643), .C2(new_n644), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n801), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n801), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n609), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(new_n800), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n834), .B1(new_n842), .B2(new_n545), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT57), .B1(new_n843), .B2(new_n413), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n809), .A2(new_n468), .A3(new_n811), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n676), .A2(new_n385), .A3(new_n704), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n326), .B1(new_n848), .B2(new_n645), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n676), .A2(new_n413), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n809), .A2(new_n688), .A3(new_n811), .A4(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n666), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n645), .A2(G141gat), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n849), .B(KEYINPUT118), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n848), .B2(new_n735), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n324), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n413), .A2(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n795), .A2(new_n609), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT119), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n783), .A2(new_n799), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n795), .A2(new_n865), .A3(new_n609), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT120), .B1(new_n841), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n840), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT117), .B1(new_n836), .B2(new_n801), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n685), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n867), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n869), .A2(new_n874), .A3(new_n545), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n861), .B1(new_n875), .B2(new_n779), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n660), .A3(new_n847), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n857), .B1(new_n878), .B2(G148gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n660), .A2(new_n324), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n859), .A2(new_n879), .B1(new_n853), .B2(new_n880), .ZN(G1345gat));
  NOR3_X1   g680(.A1(new_n848), .A2(new_n321), .A3(new_n823), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n852), .A2(new_n666), .A3(new_n544), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n321), .B2(new_n883), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n848), .B2(new_n685), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n852), .A2(new_n322), .A3(new_n829), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1347gat));
  NOR2_X1   g686(.A1(new_n688), .A2(new_n666), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n816), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G169gat), .B1(new_n889), .B2(new_n645), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n812), .B2(new_n688), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n809), .A2(KEYINPUT121), .A3(new_n385), .A4(new_n811), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n456), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n704), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n734), .A2(new_n207), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(G1348gat));
  NOR3_X1   g696(.A1(new_n889), .A2(new_n208), .A3(new_n735), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n456), .B(new_n666), .C1(new_n892), .C2(new_n893), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n660), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n900), .B2(new_n208), .ZN(G1349gat));
  INV_X1    g700(.A(new_n214), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n894), .A2(new_n902), .A3(new_n704), .A4(new_n544), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n899), .A2(KEYINPUT122), .A3(new_n902), .A4(new_n544), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G183gat), .B1(new_n889), .B2(new_n823), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  NOR3_X1   g712(.A1(new_n895), .A2(G190gat), .A3(new_n685), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT123), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n917));
  OAI221_X1 g716(.A(G190gat), .B1(new_n916), .B2(new_n917), .C1(new_n889), .C2(new_n685), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n915), .A2(new_n920), .ZN(G1351gat));
  OAI21_X1  g720(.A(KEYINPUT125), .B1(new_n860), .B2(new_n876), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n888), .A2(new_n499), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n845), .A2(KEYINPUT57), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n839), .A2(new_n840), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n868), .B1(new_n927), .B2(new_n685), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n544), .B1(new_n928), .B2(new_n873), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n834), .B1(new_n929), .B2(new_n869), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n925), .B(new_n926), .C1(new_n930), .C2(new_n861), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n922), .A2(new_n924), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n645), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n666), .B1(new_n892), .B2(new_n893), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n934), .A2(new_n850), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n632), .A3(new_n734), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(G1352gat));
  INV_X1    g736(.A(G204gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n938), .A3(new_n660), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n940));
  OAI21_X1  g739(.A(G204gat), .B1(new_n932), .B2(new_n735), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(G1353gat));
  NAND3_X1  g742(.A1(new_n935), .A2(new_n535), .A3(new_n544), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n877), .A2(new_n544), .A3(new_n924), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  NAND2_X1  g747(.A1(new_n932), .A2(KEYINPUT126), .ZN(new_n949));
  INV_X1    g748(.A(G218gat), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n685), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n922), .A2(new_n952), .A3(new_n931), .A4(new_n924), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n609), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n950), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n954), .A2(KEYINPUT127), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1355gat));
endmodule


