

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786;

  XNOR2_X1 U373 ( .A(n731), .B(KEYINPUT91), .ZN(n629) );
  BUF_X1 U374 ( .A(G116), .Z(n351) );
  XNOR2_X2 U375 ( .A(n350), .B(KEYINPUT103), .ZN(n544) );
  NAND2_X1 U376 ( .A1(n629), .A2(n413), .ZN(n350) );
  XNOR2_X2 U377 ( .A(n524), .B(n515), .ZN(n704) );
  BUF_X1 U378 ( .A(G143), .Z(n352) );
  AND2_X2 U379 ( .A1(n404), .A2(n405), .ZN(n387) );
  AND2_X2 U380 ( .A1(n388), .A2(n691), .ZN(n569) );
  NOR2_X2 U381 ( .A1(n446), .A2(KEYINPUT86), .ZN(n440) );
  XNOR2_X2 U382 ( .A(n494), .B(n493), .ZN(n509) );
  XNOR2_X1 U383 ( .A(n560), .B(KEYINPUT1), .ZN(n547) );
  INV_X1 U384 ( .A(KEYINPUT31), .ZN(n357) );
  NAND2_X1 U385 ( .A1(n364), .A2(n373), .ZN(n403) );
  NOR2_X1 U386 ( .A1(n672), .A2(n786), .ZN(n391) );
  NAND2_X1 U387 ( .A1(n356), .A2(n354), .ZN(n676) );
  NAND2_X1 U388 ( .A1(n562), .A2(n561), .ZN(n709) );
  AND2_X1 U389 ( .A1(n562), .A2(n357), .ZN(n355) );
  NAND2_X1 U390 ( .A1(n729), .A2(n562), .ZN(n353) );
  NOR2_X1 U391 ( .A1(n558), .A2(n623), .ZN(n551) );
  NAND2_X1 U392 ( .A1(n437), .A2(n435), .ZN(n434) );
  BUF_X2 U393 ( .A(n547), .Z(n731) );
  XNOR2_X1 U394 ( .A(n736), .B(KEYINPUT6), .ZN(n623) );
  NOR2_X2 U395 ( .A1(n704), .A2(G902), .ZN(n367) );
  XNOR2_X1 U396 ( .A(n360), .B(n458), .ZN(n362) );
  XNOR2_X1 U397 ( .A(n363), .B(n480), .ZN(n360) );
  INV_X1 U398 ( .A(n352), .ZN(n481) );
  NAND2_X1 U399 ( .A1(n353), .A2(KEYINPUT31), .ZN(n356) );
  INV_X1 U400 ( .A(n676), .ZN(n359) );
  NAND2_X1 U401 ( .A1(n729), .A2(n355), .ZN(n354) );
  NAND2_X1 U402 ( .A1(n358), .A2(n565), .ZN(n388) );
  NAND2_X1 U403 ( .A1(n359), .A2(n709), .ZN(n358) );
  XNOR2_X1 U404 ( .A(n456), .B(n455), .ZN(n363) );
  XNOR2_X2 U405 ( .A(n361), .B(n454), .ZN(n678) );
  XNOR2_X2 U406 ( .A(n517), .B(n496), .ZN(n361) );
  XNOR2_X2 U407 ( .A(n678), .B(n362), .ZN(n656) );
  XNOR2_X2 U408 ( .A(n452), .B(n451), .ZN(n517) );
  AND2_X1 U409 ( .A1(n694), .A2(n572), .ZN(n364) );
  BUF_X1 U410 ( .A(n678), .Z(n365) );
  BUF_X1 U411 ( .A(n692), .Z(n366) );
  NOR2_X1 U412 ( .A1(n568), .A2(n543), .ZN(n429) );
  XNOR2_X2 U413 ( .A(n626), .B(n369), .ZN(n389) );
  XNOR2_X2 U414 ( .A(n367), .B(n368), .ZN(n560) );
  XNOR2_X1 U415 ( .A(n516), .B(G469), .ZN(n368) );
  NAND2_X2 U416 ( .A1(n656), .A2(n460), .ZN(n446) );
  XNOR2_X1 U417 ( .A(G113), .B(G104), .ZN(n482) );
  NAND2_X1 U418 ( .A1(n736), .A2(n375), .ZN(n577) );
  NAND2_X1 U419 ( .A1(n612), .A2(n611), .ZN(n416) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n518) );
  XOR2_X1 U421 ( .A(KEYINPUT4), .B(G131), .Z(n449) );
  XNOR2_X1 U422 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n456) );
  XNOR2_X1 U423 ( .A(G146), .B(G125), .ZN(n480) );
  XNOR2_X1 U424 ( .A(KEYINPUT18), .B(KEYINPUT90), .ZN(n457) );
  AND2_X1 U425 ( .A1(n445), .A2(n375), .ZN(n443) );
  NOR2_X1 U426 ( .A1(n436), .A2(n462), .ZN(n435) );
  NOR2_X1 U427 ( .A1(n734), .A2(n423), .ZN(n422) );
  OR2_X1 U428 ( .A1(n651), .A2(G902), .ZN(n525) );
  XNOR2_X1 U429 ( .A(KEYINPUT16), .B(G110), .ZN(n453) );
  XNOR2_X1 U430 ( .A(n484), .B(n394), .ZN(n665) );
  XNOR2_X1 U431 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X1 U432 ( .A(G137), .B(G140), .ZN(n531) );
  XOR2_X1 U433 ( .A(G110), .B(G107), .Z(n512) );
  XNOR2_X1 U434 ( .A(G101), .B(G104), .ZN(n511) );
  NAND2_X1 U435 ( .A1(G953), .A2(G902), .ZN(n579) );
  XNOR2_X1 U436 ( .A(G902), .B(KEYINPUT15), .ZN(n502) );
  NOR2_X1 U437 ( .A1(n417), .A2(n370), .ZN(n392) );
  NAND2_X1 U438 ( .A1(n410), .A2(n570), .ZN(n409) );
  XNOR2_X1 U439 ( .A(n480), .B(KEYINPUT10), .ZN(n532) );
  INV_X1 U440 ( .A(n532), .ZN(n395) );
  XNOR2_X1 U441 ( .A(n483), .B(G122), .ZN(n396) );
  XOR2_X1 U442 ( .A(G131), .B(G140), .Z(n477) );
  XNOR2_X1 U443 ( .A(n401), .B(n571), .ZN(n400) );
  XNOR2_X1 U444 ( .A(n464), .B(KEYINPUT14), .ZN(n728) );
  NOR2_X1 U445 ( .A1(G902), .A2(G237), .ZN(n459) );
  NAND2_X1 U446 ( .A1(n460), .A2(n641), .ZN(n445) );
  INV_X1 U447 ( .A(G902), .ZN(n533) );
  XNOR2_X1 U448 ( .A(G128), .B(KEYINPUT24), .ZN(n527) );
  XNOR2_X1 U449 ( .A(G119), .B(G110), .ZN(n526) );
  XNOR2_X1 U450 ( .A(n488), .B(n487), .ZN(n530) );
  XNOR2_X1 U451 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n487) );
  XNOR2_X1 U452 ( .A(G122), .B(G107), .ZN(n496) );
  INV_X1 U453 ( .A(G134), .ZN(n493) );
  XNOR2_X1 U454 ( .A(n625), .B(KEYINPUT108), .ZN(n633) );
  NOR2_X1 U455 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U456 ( .A(KEYINPUT34), .ZN(n553) );
  AND2_X1 U457 ( .A1(n588), .A2(n587), .ZN(n616) );
  XNOR2_X1 U458 ( .A(n486), .B(G475), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n429), .B(n428), .ZN(n692) );
  INV_X1 U460 ( .A(KEYINPUT104), .ZN(n428) );
  INV_X1 U461 ( .A(G125), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n485), .B(n398), .ZN(n564) );
  INV_X1 U463 ( .A(n564), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n463), .B(KEYINPUT67), .ZN(n369) );
  AND2_X1 U465 ( .A1(n416), .A2(n415), .ZN(n370) );
  XOR2_X1 U466 ( .A(KEYINPUT93), .B(KEYINPUT75), .Z(n371) );
  OR2_X1 U467 ( .A1(n460), .A2(n641), .ZN(n372) );
  AND2_X1 U468 ( .A1(n569), .A2(n410), .ZN(n373) );
  NAND2_X1 U469 ( .A1(n397), .A2(n555), .ZN(n720) );
  INV_X1 U470 ( .A(n720), .ZN(n673) );
  AND2_X1 U471 ( .A1(n444), .A2(n445), .ZN(n374) );
  NAND2_X1 U472 ( .A1(n461), .A2(G214), .ZN(n375) );
  XOR2_X1 U473 ( .A(n546), .B(n545), .Z(n376) );
  XOR2_X1 U474 ( .A(n651), .B(KEYINPUT62), .Z(n377) );
  XNOR2_X1 U475 ( .A(KEYINPUT66), .B(n642), .ZN(n378) );
  XOR2_X1 U476 ( .A(n656), .B(n659), .Z(n379) );
  XNOR2_X1 U477 ( .A(KEYINPUT59), .B(n665), .ZN(n380) );
  XOR2_X1 U478 ( .A(n608), .B(KEYINPUT46), .Z(n381) );
  INV_X1 U479 ( .A(KEYINPUT85), .ZN(n410) );
  AND2_X1 U480 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n382) );
  XOR2_X1 U481 ( .A(n654), .B(KEYINPUT87), .Z(n383) );
  NAND2_X1 U482 ( .A1(n699), .A2(G217), .ZN(n649) );
  XNOR2_X1 U483 ( .A(n427), .B(n376), .ZN(n693) );
  NAND2_X1 U484 ( .A1(n424), .A2(n733), .ZN(n423) );
  INV_X1 U485 ( .A(n595), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n601), .B(n600), .ZN(n414) );
  XNOR2_X1 U487 ( .A(n391), .B(n381), .ZN(n390) );
  NOR2_X2 U488 ( .A1(n385), .A2(n568), .ZN(n427) );
  OR2_X1 U489 ( .A1(n568), .A2(n567), .ZN(n691) );
  NAND2_X1 U490 ( .A1(G237), .A2(G234), .ZN(n464) );
  BUF_X1 U491 ( .A(n759), .Z(n384) );
  XNOR2_X1 U492 ( .A(n551), .B(n450), .ZN(n759) );
  NAND2_X1 U493 ( .A1(n544), .A2(n623), .ZN(n385) );
  XNOR2_X2 U494 ( .A(n508), .B(n507), .ZN(n568) );
  XNOR2_X1 U495 ( .A(n554), .B(n553), .ZN(n426) );
  NAND2_X1 U496 ( .A1(n426), .A2(n618), .ZN(n425) );
  XNOR2_X1 U497 ( .A(n386), .B(n631), .ZN(n636) );
  NAND2_X1 U498 ( .A1(n390), .A2(n392), .ZN(n386) );
  NAND2_X1 U499 ( .A1(n387), .A2(n403), .ZN(n402) );
  NAND2_X1 U500 ( .A1(n389), .A2(n471), .ZN(n473) );
  AND2_X1 U501 ( .A1(n389), .A2(n414), .ZN(n714) );
  XNOR2_X1 U502 ( .A(n418), .B(n393), .ZN(n724) );
  NAND2_X1 U503 ( .A1(n630), .A2(n629), .ZN(n418) );
  NAND2_X1 U504 ( .A1(n402), .A2(n399), .ZN(n574) );
  NAND2_X1 U505 ( .A1(n400), .A2(n572), .ZN(n399) );
  NAND2_X1 U506 ( .A1(n694), .A2(n570), .ZN(n401) );
  NAND2_X1 U507 ( .A1(n411), .A2(n382), .ZN(n404) );
  NAND2_X1 U508 ( .A1(n408), .A2(n407), .ZN(n405) );
  NAND2_X1 U509 ( .A1(n406), .A2(n410), .ZN(n408) );
  INV_X1 U510 ( .A(n569), .ZN(n406) );
  NAND2_X1 U511 ( .A1(n569), .A2(n409), .ZN(n407) );
  NAND2_X1 U512 ( .A1(n572), .A2(n694), .ZN(n411) );
  INV_X1 U513 ( .A(n734), .ZN(n413) );
  NAND2_X1 U514 ( .A1(n414), .A2(n604), .ZN(n607) );
  NAND2_X1 U515 ( .A1(n610), .A2(n609), .ZN(n415) );
  NAND2_X1 U516 ( .A1(n621), .A2(n418), .ZN(n417) );
  XNOR2_X1 U517 ( .A(n419), .B(n774), .ZN(n648) );
  XNOR2_X1 U518 ( .A(n421), .B(n420), .ZN(n419) );
  XNOR2_X1 U519 ( .A(n528), .B(n529), .ZN(n420) );
  NAND2_X1 U520 ( .A1(n530), .A2(G221), .ZN(n421) );
  XNOR2_X1 U521 ( .A(n422), .B(KEYINPUT70), .ZN(n622) );
  XNOR2_X2 U522 ( .A(n540), .B(n539), .ZN(n734) );
  XNOR2_X2 U523 ( .A(n425), .B(n557), .ZN(n694) );
  AND2_X2 U524 ( .A1(n692), .A2(n693), .ZN(n572) );
  AND2_X2 U525 ( .A1(n431), .A2(n430), .ZN(n664) );
  INV_X1 U526 ( .A(n727), .ZN(n430) );
  NAND2_X1 U527 ( .A1(n432), .A2(n378), .ZN(n431) );
  XNOR2_X1 U528 ( .A(n433), .B(KEYINPUT80), .ZN(n432) );
  NAND2_X1 U529 ( .A1(n640), .A2(n639), .ZN(n433) );
  NAND2_X2 U530 ( .A1(n438), .A2(n434), .ZN(n626) );
  INV_X1 U531 ( .A(n446), .ZN(n436) );
  INV_X1 U532 ( .A(n442), .ZN(n437) );
  AND2_X2 U533 ( .A1(n439), .A2(n441), .ZN(n438) );
  INV_X1 U534 ( .A(n440), .ZN(n439) );
  NAND2_X1 U535 ( .A1(n442), .A2(n462), .ZN(n441) );
  NAND2_X1 U536 ( .A1(n374), .A2(n446), .ZN(n589) );
  NAND2_X1 U537 ( .A1(n444), .A2(n443), .ZN(n442) );
  OR2_X2 U538 ( .A1(n656), .A2(n372), .ZN(n444) );
  XNOR2_X1 U539 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U540 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n447) );
  XOR2_X1 U541 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n448) );
  XOR2_X1 U542 ( .A(n550), .B(KEYINPUT33), .Z(n450) );
  NOR2_X1 U543 ( .A1(n777), .A2(G952), .ZN(n707) );
  INV_X1 U544 ( .A(n707), .ZN(n661) );
  INV_X1 U545 ( .A(KEYINPUT68), .ZN(n571) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U547 ( .A(G953), .ZN(n465) );
  INV_X1 U548 ( .A(n695), .ZN(n696) );
  XNOR2_X2 U549 ( .A(G101), .B(G116), .ZN(n452) );
  XNOR2_X2 U550 ( .A(G119), .B(KEYINPUT3), .ZN(n451) );
  XNOR2_X1 U551 ( .A(n482), .B(n453), .ZN(n454) );
  NAND2_X1 U552 ( .A1(n465), .A2(G224), .ZN(n455) );
  XNOR2_X2 U553 ( .A(G128), .B(G143), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(n457), .ZN(n458) );
  INV_X1 U555 ( .A(n502), .ZN(n641) );
  XNOR2_X1 U556 ( .A(KEYINPUT73), .B(n459), .ZN(n461) );
  NAND2_X1 U557 ( .A1(n461), .A2(G210), .ZN(n460) );
  INV_X1 U558 ( .A(KEYINPUT86), .ZN(n462) );
  XNOR2_X1 U559 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n463) );
  BUF_X2 U560 ( .A(n465), .Z(n777) );
  AND2_X1 U561 ( .A1(n777), .A2(G952), .ZN(n583) );
  INV_X1 U562 ( .A(n583), .ZN(n469) );
  INV_X1 U563 ( .A(G898), .ZN(n467) );
  INV_X1 U564 ( .A(n579), .ZN(n466) );
  NAND2_X1 U565 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U566 ( .A1(n469), .A2(n468), .ZN(n470) );
  AND2_X1 U567 ( .A1(n728), .A2(n470), .ZN(n471) );
  INV_X1 U568 ( .A(KEYINPUT0), .ZN(n472) );
  XNOR2_X2 U569 ( .A(n473), .B(n472), .ZN(n552) );
  XNOR2_X1 U570 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n486) );
  XOR2_X1 U571 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n475) );
  XNOR2_X1 U572 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n479) );
  NAND2_X1 U574 ( .A1(G214), .A2(n518), .ZN(n476) );
  XNOR2_X1 U575 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U576 ( .A(n479), .B(n478), .ZN(n484) );
  NOR2_X1 U577 ( .A1(G902), .A2(n665), .ZN(n485) );
  NAND2_X1 U578 ( .A1(n777), .A2(G234), .ZN(n488) );
  NAND2_X1 U579 ( .A1(G217), .A2(n530), .ZN(n492) );
  XOR2_X1 U580 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n490) );
  XNOR2_X1 U581 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U582 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U583 ( .A(n492), .B(n491), .ZN(n499) );
  XNOR2_X1 U584 ( .A(n351), .B(KEYINPUT9), .ZN(n495) );
  XNOR2_X1 U585 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U586 ( .A(n509), .B(n497), .ZN(n498) );
  XNOR2_X1 U587 ( .A(n499), .B(n498), .ZN(n695) );
  NAND2_X1 U588 ( .A1(n695), .A2(n533), .ZN(n501) );
  INV_X1 U589 ( .A(G478), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n501), .B(n500), .ZN(n555) );
  NAND2_X1 U591 ( .A1(n564), .A2(n555), .ZN(n746) );
  NAND2_X1 U592 ( .A1(n502), .A2(G234), .ZN(n503) );
  XNOR2_X1 U593 ( .A(n503), .B(KEYINPUT20), .ZN(n534) );
  AND2_X1 U594 ( .A1(n534), .A2(G221), .ZN(n504) );
  XNOR2_X1 U595 ( .A(n504), .B(KEYINPUT21), .ZN(n733) );
  INV_X1 U596 ( .A(n733), .ZN(n505) );
  NOR2_X1 U597 ( .A1(n746), .A2(n505), .ZN(n506) );
  AND2_X2 U598 ( .A1(n552), .A2(n506), .ZN(n508) );
  INV_X1 U599 ( .A(KEYINPUT22), .ZN(n507) );
  XNOR2_X2 U600 ( .A(n509), .B(n449), .ZN(n775) );
  XNOR2_X2 U601 ( .A(n775), .B(G146), .ZN(n524) );
  NAND2_X1 U602 ( .A1(n777), .A2(G227), .ZN(n510) );
  XNOR2_X1 U603 ( .A(n531), .B(n510), .ZN(n514) );
  XNOR2_X1 U604 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U605 ( .A(n514), .B(n513), .ZN(n515) );
  INV_X1 U606 ( .A(KEYINPUT71), .ZN(n516) );
  INV_X1 U607 ( .A(n731), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n518), .A2(G210), .ZN(n519) );
  XNOR2_X1 U609 ( .A(n519), .B(G113), .ZN(n521) );
  XNOR2_X1 U610 ( .A(KEYINPUT5), .B(G137), .ZN(n520) );
  XNOR2_X1 U611 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U612 ( .A(n517), .B(n522), .ZN(n523) );
  XNOR2_X1 U613 ( .A(n524), .B(n523), .ZN(n651) );
  XNOR2_X2 U614 ( .A(n525), .B(G472), .ZN(n736) );
  XNOR2_X1 U615 ( .A(n526), .B(KEYINPUT23), .ZN(n529) );
  XNOR2_X1 U616 ( .A(n371), .B(n527), .ZN(n528) );
  XNOR2_X1 U617 ( .A(n532), .B(n531), .ZN(n774) );
  NAND2_X1 U618 ( .A1(n648), .A2(n533), .ZN(n540) );
  XNOR2_X1 U619 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n536) );
  AND2_X1 U620 ( .A1(n534), .A2(G217), .ZN(n535) );
  XNOR2_X1 U621 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U622 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n537) );
  XNOR2_X1 U623 ( .A(n538), .B(n537), .ZN(n539) );
  OR2_X1 U624 ( .A1(n736), .A2(n734), .ZN(n541) );
  OR2_X1 U625 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U626 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n546) );
  INV_X1 U627 ( .A(KEYINPUT65), .ZN(n545) );
  NAND2_X1 U628 ( .A1(n734), .A2(n733), .ZN(n730) );
  NOR2_X1 U629 ( .A1(n547), .A2(n730), .ZN(n549) );
  INV_X1 U630 ( .A(KEYINPUT72), .ZN(n548) );
  XNOR2_X1 U631 ( .A(n549), .B(n548), .ZN(n558) );
  INV_X1 U632 ( .A(KEYINPUT89), .ZN(n550) );
  BUF_X2 U633 ( .A(n552), .Z(n562) );
  NAND2_X1 U634 ( .A1(n759), .A2(n562), .ZN(n554) );
  INV_X1 U635 ( .A(n555), .ZN(n563) );
  NAND2_X1 U636 ( .A1(n397), .A2(n563), .ZN(n556) );
  XNOR2_X1 U637 ( .A(n556), .B(KEYINPUT105), .ZN(n618) );
  INV_X1 U638 ( .A(KEYINPUT35), .ZN(n557) );
  INV_X1 U639 ( .A(n558), .ZN(n559) );
  AND2_X1 U640 ( .A1(n559), .A2(n736), .ZN(n729) );
  OR2_X1 U641 ( .A1(n560), .A2(n730), .ZN(n586) );
  NOR2_X1 U642 ( .A1(n586), .A2(n736), .ZN(n561) );
  NAND2_X1 U643 ( .A1(n564), .A2(n563), .ZN(n715) );
  NAND2_X1 U644 ( .A1(n720), .A2(n715), .ZN(n747) );
  INV_X1 U645 ( .A(KEYINPUT79), .ZN(n613) );
  XNOR2_X1 U646 ( .A(n747), .B(n613), .ZN(n565) );
  AND2_X1 U647 ( .A1(n731), .A2(n734), .ZN(n566) );
  NAND2_X1 U648 ( .A1(n566), .A2(n623), .ZN(n567) );
  INV_X1 U649 ( .A(KEYINPUT44), .ZN(n570) );
  XNOR2_X1 U650 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n573) );
  XNOR2_X1 U651 ( .A(n574), .B(n573), .ZN(n643) );
  NAND2_X1 U652 ( .A1(n643), .A2(n641), .ZN(n575) );
  XNOR2_X1 U653 ( .A(n575), .B(KEYINPUT81), .ZN(n640) );
  INV_X1 U654 ( .A(KEYINPUT30), .ZN(n576) );
  XNOR2_X1 U655 ( .A(n577), .B(n576), .ZN(n588) );
  INV_X1 U656 ( .A(n728), .ZN(n578) );
  NOR2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U658 ( .A(KEYINPUT106), .B(n580), .Z(n581) );
  NOR2_X1 U659 ( .A1(G900), .A2(n581), .ZN(n582) );
  XNOR2_X1 U660 ( .A(n582), .B(KEYINPUT107), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n728), .A2(n583), .ZN(n584) );
  AND2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n595) );
  NOR2_X1 U663 ( .A1(n586), .A2(n595), .ZN(n587) );
  XNOR2_X1 U664 ( .A(n589), .B(KEYINPUT38), .ZN(n744) );
  NAND2_X1 U665 ( .A1(n616), .A2(n744), .ZN(n591) );
  INV_X1 U666 ( .A(KEYINPUT39), .ZN(n590) );
  XNOR2_X1 U667 ( .A(n591), .B(n590), .ZN(n638) );
  INV_X1 U668 ( .A(n638), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n592), .A2(n673), .ZN(n594) );
  INV_X1 U670 ( .A(KEYINPUT40), .ZN(n593) );
  XNOR2_X1 U671 ( .A(n594), .B(n593), .ZN(n672) );
  NAND2_X1 U672 ( .A1(n622), .A2(n736), .ZN(n597) );
  INV_X1 U673 ( .A(KEYINPUT28), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n597), .B(n596), .ZN(n599) );
  INV_X1 U675 ( .A(n560), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n601) );
  INV_X1 U677 ( .A(KEYINPUT110), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n744), .A2(n375), .ZN(n748) );
  NOR2_X1 U679 ( .A1(n746), .A2(n748), .ZN(n603) );
  XOR2_X1 U680 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n602) );
  XNOR2_X1 U681 ( .A(n603), .B(n602), .ZN(n760) );
  INV_X1 U682 ( .A(n760), .ZN(n604) );
  INV_X1 U683 ( .A(KEYINPUT112), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n605), .B(KEYINPUT42), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n607), .B(n606), .ZN(n786) );
  INV_X1 U686 ( .A(KEYINPUT64), .ZN(n608) );
  AND2_X1 U687 ( .A1(n714), .A2(n747), .ZN(n610) );
  INV_X1 U688 ( .A(KEYINPUT47), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n613), .A2(n611), .ZN(n609) );
  INV_X1 U690 ( .A(n610), .ZN(n612) );
  NOR2_X1 U691 ( .A1(n747), .A2(n613), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n714), .A2(n614), .ZN(n620) );
  INV_X1 U693 ( .A(n589), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U695 ( .A(n617), .B(KEYINPUT109), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n719) );
  AND2_X1 U697 ( .A1(n620), .A2(n719), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n673), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n633), .A2(n626), .ZN(n628) );
  INV_X1 U700 ( .A(KEYINPUT36), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n630) );
  INV_X1 U702 ( .A(KEYINPUT48), .ZN(n631) );
  AND2_X1 U703 ( .A1(n731), .A2(n375), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n634), .B(KEYINPUT43), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n635), .A2(n589), .ZN(n690) );
  NAND2_X1 U707 ( .A1(n636), .A2(n690), .ZN(n637) );
  XNOR2_X2 U708 ( .A(n637), .B(KEYINPUT83), .ZN(n647) );
  OR2_X1 U709 ( .A1(n638), .A2(n715), .ZN(n670) );
  NAND2_X2 U710 ( .A1(n647), .A2(n670), .ZN(n776) );
  INV_X1 U711 ( .A(n776), .ZN(n639) );
  NAND2_X1 U712 ( .A1(n641), .A2(KEYINPUT2), .ZN(n642) );
  BUF_X1 U713 ( .A(n643), .Z(n644) );
  INV_X1 U714 ( .A(n644), .ZN(n681) );
  NAND2_X1 U715 ( .A1(n670), .A2(KEYINPUT2), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT77), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n767) );
  NOR2_X1 U718 ( .A1(n681), .A2(n767), .ZN(n727) );
  BUF_X2 U719 ( .A(n664), .Z(n699) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n650) );
  AND2_X1 U721 ( .A1(n650), .A2(n661), .ZN(G66) );
  NAND2_X1 U722 ( .A1(n664), .A2(G472), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n652), .B(n377), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n653), .A2(n661), .ZN(n655) );
  XNOR2_X1 U725 ( .A(KEYINPUT92), .B(KEYINPUT63), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n655), .B(n383), .ZN(G57) );
  NAND2_X1 U727 ( .A1(n664), .A2(G210), .ZN(n660) );
  XOR2_X1 U728 ( .A(KEYINPUT78), .B(KEYINPUT88), .Z(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n660), .B(n379), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(n448), .ZN(G51) );
  NAND2_X1 U734 ( .A1(n664), .A2(G475), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n666), .B(n380), .ZN(n667) );
  NAND2_X1 U736 ( .A1(n667), .A2(n661), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n668), .B(n447), .ZN(G60) );
  XNOR2_X1 U738 ( .A(G134), .B(KEYINPUT116), .ZN(n669) );
  XNOR2_X1 U739 ( .A(n670), .B(n669), .ZN(G36) );
  XNOR2_X1 U740 ( .A(G131), .B(KEYINPUT127), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(G33) );
  NAND2_X1 U742 ( .A1(n676), .A2(n673), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n674), .B(G113), .ZN(G15) );
  INV_X1 U744 ( .A(n715), .ZN(n675) );
  NAND2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(n351), .ZN(G18) );
  INV_X1 U747 ( .A(n365), .ZN(n680) );
  OR2_X1 U748 ( .A1(n777), .A2(G898), .ZN(n679) );
  NAND2_X1 U749 ( .A1(n680), .A2(n679), .ZN(n688) );
  NAND2_X1 U750 ( .A1(n644), .A2(n777), .ZN(n686) );
  NAND2_X1 U751 ( .A1(G224), .A2(G953), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n682), .B(KEYINPUT61), .ZN(n683) );
  XNOR2_X1 U753 ( .A(KEYINPUT124), .B(n683), .ZN(n684) );
  NAND2_X1 U754 ( .A1(G898), .A2(n684), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U756 ( .A(n688), .B(n687), .Z(G69) );
  XOR2_X1 U757 ( .A(G140), .B(KEYINPUT117), .Z(n689) );
  XNOR2_X1 U758 ( .A(n690), .B(n689), .ZN(G42) );
  XNOR2_X1 U759 ( .A(n691), .B(G101), .ZN(G3) );
  XNOR2_X1 U760 ( .A(n366), .B(G110), .ZN(G12) );
  XNOR2_X1 U761 ( .A(n693), .B(G119), .ZN(G21) );
  XNOR2_X1 U762 ( .A(n694), .B(G122), .ZN(G24) );
  NAND2_X1 U763 ( .A1(n699), .A2(G478), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n698), .A2(n707), .ZN(G63) );
  NAND2_X1 U765 ( .A1(n699), .A2(G469), .ZN(n706) );
  XNOR2_X1 U766 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(KEYINPUT120), .ZN(n702) );
  XNOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n701) );
  XNOR2_X1 U769 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U770 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U771 ( .A(n706), .B(n705), .ZN(n708) );
  NOR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(G54) );
  NOR2_X1 U773 ( .A1(n709), .A2(n720), .ZN(n710) );
  XOR2_X1 U774 ( .A(G104), .B(n710), .Z(G6) );
  NOR2_X1 U775 ( .A1(n709), .A2(n715), .ZN(n712) );
  XNOR2_X1 U776 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U778 ( .A(G107), .B(n713), .ZN(G9) );
  INV_X1 U779 ( .A(n714), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n721), .A2(n715), .ZN(n717) );
  XNOR2_X1 U781 ( .A(KEYINPUT29), .B(KEYINPUT113), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n717), .B(n716), .ZN(n718) );
  XOR2_X1 U783 ( .A(G128), .B(n718), .Z(G30) );
  XNOR2_X1 U784 ( .A(n352), .B(n719), .ZN(G45) );
  NOR2_X1 U785 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U786 ( .A(KEYINPUT114), .B(n722), .Z(n723) );
  XNOR2_X1 U787 ( .A(G146), .B(n723), .ZN(G48) );
  XOR2_X1 U788 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n725) );
  XNOR2_X1 U789 ( .A(n725), .B(n724), .ZN(G27) );
  INV_X1 U790 ( .A(KEYINPUT2), .ZN(n726) );
  NOR2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n766) );
  NAND2_X1 U792 ( .A1(G952), .A2(n728), .ZN(n757) );
  INV_X1 U793 ( .A(n729), .ZN(n741) );
  NAND2_X1 U794 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U795 ( .A(n732), .B(KEYINPUT50), .ZN(n739) );
  NOR2_X1 U796 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U797 ( .A(KEYINPUT49), .B(n735), .Z(n737) );
  NOR2_X1 U798 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U799 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U800 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U801 ( .A(KEYINPUT51), .B(n742), .ZN(n743) );
  NOR2_X1 U802 ( .A1(n760), .A2(n743), .ZN(n754) );
  NOR2_X1 U803 ( .A1(n744), .A2(n375), .ZN(n745) );
  NOR2_X1 U804 ( .A1(n746), .A2(n745), .ZN(n751) );
  INV_X1 U805 ( .A(n747), .ZN(n749) );
  NOR2_X1 U806 ( .A1(n749), .A2(n748), .ZN(n750) );
  OR2_X1 U807 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U808 ( .A1(n384), .A2(n752), .ZN(n753) );
  NOR2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U810 ( .A(n755), .B(KEYINPUT52), .ZN(n756) );
  NOR2_X1 U811 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U812 ( .A(n758), .B(KEYINPUT118), .ZN(n763) );
  INV_X1 U813 ( .A(n384), .ZN(n761) );
  NOR2_X1 U814 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U815 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U816 ( .A(n764), .B(KEYINPUT119), .ZN(n765) );
  NOR2_X1 U817 ( .A1(n766), .A2(n765), .ZN(n771) );
  INV_X1 U818 ( .A(n767), .ZN(n768) );
  NOR2_X1 U819 ( .A1(n768), .A2(n776), .ZN(n769) );
  NAND2_X1 U820 ( .A1(n769), .A2(n644), .ZN(n770) );
  NAND2_X1 U821 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U822 ( .A1(n772), .A2(G953), .ZN(n773) );
  XNOR2_X1 U823 ( .A(n773), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U824 ( .A(n775), .B(n774), .Z(n779) );
  XNOR2_X1 U825 ( .A(n776), .B(n779), .ZN(n778) );
  NAND2_X1 U826 ( .A1(n778), .A2(n777), .ZN(n784) );
  XOR2_X1 U827 ( .A(G227), .B(n779), .Z(n780) );
  XNOR2_X1 U828 ( .A(n780), .B(KEYINPUT125), .ZN(n781) );
  NAND2_X1 U829 ( .A1(n781), .A2(G900), .ZN(n782) );
  NAND2_X1 U830 ( .A1(n782), .A2(G953), .ZN(n783) );
  NAND2_X1 U831 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U832 ( .A(KEYINPUT126), .B(n785), .ZN(G72) );
  XOR2_X1 U833 ( .A(G137), .B(n786), .Z(G39) );
endmodule

