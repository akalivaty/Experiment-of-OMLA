//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT23), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT64), .A4(new_n208), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n211), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(KEYINPUT65), .A3(new_n221), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  OAI221_X1 g025(.A(new_n207), .B1(new_n226), .B2(new_n203), .C1(new_n204), .C2(KEYINPUT66), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT25), .A3(new_n218), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT68), .B(G113gat), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G120gat), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G113gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT1), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  INV_X1    g037(.A(new_n233), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n232), .A2(G113gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n234), .A2(new_n235), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT27), .B(G183gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n206), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n244), .B(KEYINPUT28), .Z(new_n245));
  AOI21_X1  g044(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(G169gat), .B2(G176gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT26), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .A4(new_n202), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n242), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n229), .A2(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n235), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n241), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n229), .A2(KEYINPUT69), .A3(new_n242), .A4(new_n249), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n252), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT32), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT33), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G15gat), .B(G43gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G71gat), .B(G99gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT32), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n270), .B1(new_n259), .B2(new_n261), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT33), .B1(new_n259), .B2(new_n261), .ZN(new_n272));
  INV_X1    g071(.A(new_n268), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n252), .A2(new_n257), .A3(new_n260), .A4(new_n258), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT34), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n269), .A2(new_n277), .A3(new_n274), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n253), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G226gat), .ZN(new_n284));
  INV_X1    g083(.A(G233gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(KEYINPUT73), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT29), .B1(new_n229), .B2(new_n249), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n253), .A2(new_n286), .ZN(new_n292));
  OR2_X1    g091(.A1(KEYINPUT71), .A2(KEYINPUT22), .ZN(new_n293));
  NAND2_X1  g092(.A1(KEYINPUT71), .A2(KEYINPUT22), .ZN(new_n294));
  INV_X1    g093(.A(G211gat), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n299), .B(KEYINPUT72), .Z(new_n300));
  XOR2_X1   g099(.A(G211gat), .B(G218gat), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n300), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n291), .A3(new_n292), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n292), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n286), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT74), .B(G64gat), .Z(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT75), .B(G92gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT30), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT77), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n305), .A2(new_n308), .A3(KEYINPUT30), .A4(new_n314), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n308), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n313), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(KEYINPUT76), .A3(new_n313), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n322), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n303), .B2(KEYINPUT29), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G141gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G141gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT78), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G141gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n335), .B1(new_n340), .B2(G148gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n332), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n345), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n342), .B1(new_n348), .B2(KEYINPUT2), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n333), .B1(new_n337), .B2(new_n339), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n349), .B(KEYINPUT79), .C1(new_n350), .C2(new_n335), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n336), .A2(G148gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g153(.A(new_n345), .B(new_n343), .C1(new_n354), .C2(new_n344), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n331), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n347), .B2(new_n351), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n359), .A2(new_n360), .A3(new_n330), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n359), .B2(new_n330), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT29), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n358), .B1(new_n364), .B2(new_n304), .ZN(new_n365));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n366), .B(G22gat), .Z(new_n367));
  AND2_X1   g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n358), .B(new_n369), .C1(new_n364), .C2(new_n304), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(G50gat), .ZN(new_n374));
  XOR2_X1   g173(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n376), .A2(KEYINPUT84), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n376), .A2(KEYINPUT84), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n367), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(new_n370), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n281), .A2(new_n329), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n256), .B(new_n387), .C1(new_n361), .C2(new_n362), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n242), .A2(new_n359), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT4), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n242), .A2(new_n359), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n388), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n357), .A2(new_n256), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n390), .ZN(new_n397));
  INV_X1    g196(.A(new_n389), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT5), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G1gat), .B(G29gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(G85gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT0), .B(G57gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n388), .A2(KEYINPUT5), .A3(new_n389), .A4(new_n394), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n407), .A2(new_n408), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT88), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n401), .A2(new_n406), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n405), .B(KEYINPUT85), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  INV_X1    g214(.A(new_n405), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n395), .A2(new_n400), .ZN(new_n417));
  INV_X1    g216(.A(new_n406), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n412), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n405), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n408), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n411), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT35), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n386), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT70), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n431));
  AOI221_X4 g230(.A(new_n270), .B1(KEYINPUT33), .B2(new_n268), .C1(new_n259), .C2(new_n261), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n277), .B1(new_n269), .B2(new_n274), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n277), .A2(new_n433), .B1(new_n434), .B2(new_n430), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n429), .B1(new_n435), .B2(new_n385), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n401), .A2(new_n405), .A3(new_n406), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n415), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n421), .A3(new_n423), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n321), .A2(new_n439), .A3(new_n328), .A4(new_n322), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT82), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n315), .A2(new_n319), .A3(new_n316), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n319), .B1(new_n315), .B2(new_n316), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT76), .B1(new_n323), .B2(new_n313), .ZN(new_n445));
  AOI211_X1 g244(.A(new_n325), .B(new_n314), .C1(new_n305), .C2(new_n308), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n322), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT82), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n439), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n383), .B1(new_n372), .B2(new_n377), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n278), .B1(new_n275), .B2(new_n430), .ZN(new_n452));
  AOI211_X1 g251(.A(KEYINPUT70), .B(new_n277), .C1(new_n269), .C2(new_n274), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(KEYINPUT91), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n436), .A2(new_n441), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT35), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n428), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n389), .B1(new_n388), .B2(new_n394), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT39), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n397), .A2(new_n398), .ZN(new_n462));
  OR3_X1    g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n413), .B1(new_n460), .B2(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT40), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n466), .B(new_n414), .C1(new_n444), .C2(new_n447), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n329), .A2(KEYINPUT86), .A3(new_n414), .A4(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n305), .A2(new_n472), .A3(new_n308), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n288), .A2(new_n291), .A3(new_n292), .A4(new_n303), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(KEYINPUT37), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT38), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n473), .A2(new_n476), .A3(new_n477), .A4(new_n313), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n315), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n478), .A2(new_n479), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n425), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n323), .A2(KEYINPUT37), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n313), .A3(new_n473), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT38), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n489), .A3(new_n451), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n435), .A2(KEYINPUT36), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(KEYINPUT36), .B2(new_n281), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n441), .A2(new_n450), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n385), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n385), .B1(new_n483), .B2(new_n488), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT90), .A3(new_n471), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n492), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n459), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n501), .A2(KEYINPUT96), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(KEYINPUT96), .ZN(new_n503));
  OR3_X1    g302(.A1(new_n502), .A2(new_n503), .A3(G1gat), .ZN(new_n504));
  AOI21_X1  g303(.A(G8gat), .B1(new_n504), .B2(KEYINPUT97), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT16), .ZN(new_n506));
  OAI22_X1  g305(.A1(new_n502), .A2(new_n503), .B1(new_n506), .B2(G1gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n505), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(KEYINPUT94), .Z(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(KEYINPUT15), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  OR3_X1    g313(.A1(new_n514), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT95), .B(G36gat), .Z(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n515), .B(new_n516), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n520), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n509), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n526), .A2(new_n509), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT18), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n509), .B(new_n524), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n530), .B(KEYINPUT13), .Z(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(KEYINPUT93), .B(KEYINPUT11), .Z(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G169gat), .B(G197gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n541), .B(KEYINPUT12), .Z(new_n542));
  OR2_X1    g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n536), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT7), .ZN(new_n548));
  INV_X1    g347(.A(G99gat), .ZN(new_n549));
  INV_X1    g348(.A(G106gat), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT101), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT101), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(G99gat), .A3(G106gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(KEYINPUT8), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT102), .B(G85gat), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n548), .B(new_n554), .C1(G92gat), .C2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G99gat), .B(G106gat), .Z(new_n557));
  OR2_X1    g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT10), .ZN(new_n561));
  XOR2_X1   g360(.A(G57gat), .B(G64gat), .Z(new_n562));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563));
  INV_X1    g362(.A(G71gat), .ZN(new_n564));
  INV_X1    g363(.A(G78gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n560), .A2(new_n561), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT105), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n558), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n560), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n571), .B1(new_n574), .B2(new_n561), .ZN(new_n575));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n576), .B2(new_n574), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT106), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n581), .B(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n546), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n509), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n205), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT19), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G211gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT20), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n600), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n560), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT103), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n528), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT17), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n521), .B2(new_n523), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G134gat), .B(G162gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT104), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n612), .B(new_n616), .ZN(new_n617));
  AND4_X1   g416(.A1(new_n500), .A2(new_n587), .A3(new_n603), .A4(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n439), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n329), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G8gat), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(KEYINPUT107), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(KEYINPUT107), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT16), .B(G8gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT42), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n622), .A2(KEYINPUT42), .A3(new_n626), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n624), .A2(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT108), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT108), .ZN(new_n633));
  OAI221_X1 g432(.A(new_n633), .B1(new_n629), .B2(new_n630), .C1(new_n624), .C2(new_n625), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(G1325gat));
  INV_X1    g434(.A(new_n281), .ZN(new_n636));
  AOI21_X1  g435(.A(G15gat), .B1(new_n618), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n618), .A2(new_n494), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(G15gat), .B2(new_n638), .ZN(G1326gat));
  NAND2_X1  g438(.A1(new_n618), .A2(new_n385), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G22gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  AOI21_X1  g442(.A(new_n617), .B1(new_n459), .B2(new_n499), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n601), .A2(new_n602), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n645), .A2(new_n587), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n519), .A3(new_n619), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT110), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT45), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n612), .B(new_n616), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT113), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT113), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n617), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(KEYINPUT44), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n459), .A2(KEYINPUT112), .A3(new_n499), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT112), .B1(new_n459), .B2(new_n499), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT114), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT92), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT35), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n665), .A2(new_n666), .B1(new_n386), .B2(new_n427), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n497), .A2(KEYINPUT90), .A3(new_n471), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT90), .B1(new_n497), .B2(new_n471), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n495), .A2(new_n385), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n281), .A2(KEYINPUT36), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(KEYINPUT36), .B2(new_n435), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n654), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT44), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT114), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n677), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n646), .B(KEYINPUT111), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n679), .A2(new_n619), .A3(new_n680), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n652), .B(new_n653), .C1(new_n519), .C2(new_n681), .ZN(G1328gat));
  NAND3_X1  g481(.A1(new_n648), .A2(new_n329), .A3(new_n518), .ZN(new_n683));
  AND2_X1   g482(.A1(KEYINPUT115), .A2(KEYINPUT46), .ZN(new_n684));
  NOR2_X1   g483(.A1(KEYINPUT115), .A2(KEYINPUT46), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n679), .A2(new_n329), .A3(new_n680), .ZN(new_n687));
  OAI221_X1 g486(.A(new_n686), .B1(new_n684), .B2(new_n683), .C1(new_n687), .C2(new_n518), .ZN(G1329gat));
  NOR3_X1   g487(.A1(new_n647), .A2(G43gat), .A3(new_n281), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n679), .A2(new_n494), .A3(new_n680), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(G43gat), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI211_X1 g492(.A(KEYINPUT47), .B(new_n689), .C1(new_n690), .C2(G43gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(G1330gat));
  NOR3_X1   g494(.A1(new_n647), .A2(G50gat), .A3(new_n451), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n679), .A2(new_n385), .A3(new_n680), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(G50gat), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI211_X1 g499(.A(KEYINPUT48), .B(new_n696), .C1(new_n697), .C2(G50gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(G1331gat));
  NOR2_X1   g501(.A1(new_n660), .A2(new_n661), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n603), .A2(new_n617), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n586), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n545), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n439), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT116), .B(G57gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  INV_X1    g510(.A(new_n708), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT49), .B(G64gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n329), .A3(new_n713), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n708), .A2(new_n448), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT117), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1333gat));
  NAND3_X1  g517(.A1(new_n712), .A2(new_n564), .A3(new_n636), .ZN(new_n719));
  OAI21_X1  g518(.A(G71gat), .B1(new_n708), .B2(new_n672), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1334gat));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n451), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(new_n565), .ZN(G1335gat));
  NAND2_X1  g524(.A1(new_n675), .A2(KEYINPUT118), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n603), .A2(new_n545), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT118), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n644), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n728), .B1(new_n500), .B2(new_n654), .ZN(new_n733));
  AOI211_X1 g532(.A(KEYINPUT118), .B(new_n617), .C1(new_n459), .C2(new_n499), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(KEYINPUT51), .A3(new_n727), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n706), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n555), .B1(new_n737), .B2(new_n619), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n645), .A2(new_n707), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n679), .A2(new_n619), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n738), .B1(new_n555), .B2(new_n740), .ZN(G1336gat));
  NAND3_X1  g540(.A1(new_n679), .A2(new_n329), .A3(new_n739), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G92gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n448), .A2(G92gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT119), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT51), .B1(new_n735), .B2(new_n727), .ZN(new_n749));
  AND4_X1   g548(.A1(KEYINPUT51), .A2(new_n726), .A3(new_n727), .A4(new_n729), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n732), .A2(KEYINPUT119), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n744), .A2(new_n586), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n753), .A2(new_n754), .B1(G92gat), .B2(new_n742), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n747), .B1(new_n755), .B2(new_n746), .ZN(G1337gat));
  NAND3_X1  g555(.A1(new_n737), .A2(new_n549), .A3(new_n636), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n679), .A2(new_n494), .A3(new_n739), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n549), .B2(new_n758), .ZN(G1338gat));
  NAND3_X1  g558(.A1(new_n679), .A2(new_n385), .A3(new_n739), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G106gat), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n706), .A2(G106gat), .A3(new_n451), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n749), .B2(new_n750), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n753), .A2(new_n762), .B1(G106gat), .B2(new_n760), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(G1339gat));
  NAND4_X1  g567(.A1(new_n603), .A2(new_n546), .A3(new_n706), .A4(new_n617), .ZN(new_n769));
  INV_X1    g568(.A(new_n658), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n584), .B1(new_n578), .B2(KEYINPUT54), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n575), .B2(new_n577), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n578), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT55), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n579), .A2(new_n584), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n545), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n529), .A2(new_n530), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n533), .A2(new_n534), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n541), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n543), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n586), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n770), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n777), .A2(new_n782), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(new_n658), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n645), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n769), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n439), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n386), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(KEYINPUT121), .A3(new_n386), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G113gat), .B1(new_n794), .B2(new_n546), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n436), .A2(new_n454), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n789), .A2(new_n448), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n230), .A3(new_n545), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1340gat));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n232), .A3(new_n586), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n792), .A2(new_n586), .A3(new_n793), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT122), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n802), .A2(new_n803), .A3(G120gat), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n802), .B2(G120gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(G1341gat));
  NAND4_X1  g605(.A1(new_n792), .A2(G127gat), .A3(new_n603), .A4(new_n793), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(KEYINPUT123), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(KEYINPUT123), .ZN(new_n809));
  AOI21_X1  g608(.A(G127gat), .B1(new_n798), .B2(new_n603), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(G1342gat));
  NOR3_X1   g610(.A1(new_n797), .A2(G134gat), .A3(new_n617), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT56), .ZN(new_n813));
  OAI21_X1  g612(.A(G134gat), .B1(new_n794), .B2(new_n617), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1343gat));
  NOR2_X1   g614(.A1(new_n788), .A2(new_n451), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n778), .A2(new_n783), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n778), .A2(new_n783), .A3(KEYINPUT124), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n617), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n786), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n603), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n769), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n385), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT57), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n494), .A2(new_n439), .A3(new_n329), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n818), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n340), .B1(new_n830), .B2(new_n545), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n829), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n545), .A2(new_n336), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT58), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n828), .A3(new_n829), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n337), .B(new_n339), .C1(new_n836), .C2(new_n546), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n837), .B(new_n838), .C1(new_n832), .C2(new_n833), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(G1344gat));
  INV_X1    g639(.A(new_n832), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n333), .A3(new_n586), .ZN(new_n842));
  AOI211_X1 g641(.A(KEYINPUT59), .B(new_n333), .C1(new_n830), .C2(new_n586), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT57), .B1(new_n788), .B2(new_n451), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n777), .A2(new_n782), .A3(new_n654), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n603), .B1(new_n823), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n817), .B(new_n385), .C1(new_n847), .C2(new_n826), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n845), .A2(new_n848), .A3(new_n586), .A4(new_n829), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n849), .B2(G148gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n842), .B1(new_n843), .B2(new_n850), .ZN(G1345gat));
  AOI21_X1  g650(.A(G155gat), .B1(new_n841), .B2(new_n603), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n830), .A2(G155gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n603), .ZN(G1346gat));
  NAND3_X1  g653(.A1(new_n830), .A2(KEYINPUT125), .A3(new_n770), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n836), .B2(new_n658), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(G162gat), .A3(new_n857), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n832), .A2(G162gat), .A3(new_n617), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1347gat));
  NOR2_X1   g659(.A1(new_n788), .A2(new_n619), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n861), .A2(new_n329), .A3(new_n796), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n212), .A3(new_n545), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n281), .A2(new_n385), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(new_n329), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G169gat), .B1(new_n865), .B2(new_n546), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n866), .ZN(G1348gat));
  AOI21_X1  g666(.A(G176gat), .B1(new_n862), .B2(new_n586), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n865), .A2(new_n213), .A3(new_n706), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(G1349gat));
  OAI21_X1  g669(.A(G183gat), .B1(new_n865), .B2(new_n645), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n862), .A2(new_n243), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n645), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g673(.A1(new_n862), .A2(new_n206), .A3(new_n770), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n876));
  INV_X1    g675(.A(new_n865), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n654), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(G190gat), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT61), .B(new_n206), .C1(new_n877), .C2(new_n654), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(G1351gat));
  NOR2_X1   g680(.A1(new_n494), .A2(new_n448), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n845), .A2(new_n848), .A3(new_n439), .A4(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G197gat), .B1(new_n883), .B2(new_n546), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n861), .A2(new_n385), .A3(new_n882), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n885), .A2(G197gat), .A3(new_n546), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(KEYINPUT126), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(KEYINPUT126), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(G1352gat));
  OR3_X1    g688(.A1(new_n883), .A2(KEYINPUT127), .A3(new_n706), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT127), .B1(new_n883), .B2(new_n706), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(G204gat), .A3(new_n891), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n885), .A2(G204gat), .A3(new_n706), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT62), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(KEYINPUT62), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(G1353gat));
  INV_X1    g695(.A(new_n885), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n295), .A3(new_n603), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n883), .A2(new_n645), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT63), .B1(new_n899), .B2(G211gat), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT63), .B(G211gat), .C1(new_n883), .C2(new_n645), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(G1354gat));
  OAI21_X1  g702(.A(G218gat), .B1(new_n883), .B2(new_n617), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n897), .A2(new_n296), .A3(new_n770), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1355gat));
endmodule


