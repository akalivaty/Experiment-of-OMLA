//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT87), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT77), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT3), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G107), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G104), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n196), .A2(new_n198), .B1(new_n193), .B2(KEYINPUT3), .ZN(new_n199));
  OAI21_X1  g013(.A(G101), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n194), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n198), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n197), .A2(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n194), .B1(new_n203), .B2(new_n190), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(new_n206), .A3(KEYINPUT4), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT70), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n209));
  INV_X1    g023(.A(G113), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(KEYINPUT70), .A2(KEYINPUT2), .A3(G113), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G116), .ZN(new_n217));
  INV_X1    g031(.A(G116), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G119), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n211), .A2(new_n212), .B1(new_n209), .B2(new_n210), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n226), .B(G101), .C1(new_n195), .C2(new_n199), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n207), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n203), .B2(new_n190), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n206), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n220), .A2(KEYINPUT5), .ZN(new_n231));
  OAI21_X1  g045(.A(G113), .B1(new_n217), .B2(KEYINPUT5), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n231), .A2(new_n233), .B1(new_n223), .B2(new_n220), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G110), .B(G122), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n228), .A2(new_n235), .A3(new_n237), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT6), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n236), .A2(new_n242), .A3(new_n238), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g060(.A(G128), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n244), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT65), .A2(G143), .ZN(new_n250));
  AOI21_X1  g064(.A(G146), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n247), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G125), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(G146), .A3(new_n250), .ZN(new_n256));
  INV_X1    g070(.A(new_n245), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n254), .A2(new_n255), .A3(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n251), .B2(new_n253), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n256), .A2(new_n262), .A3(new_n257), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n255), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n268), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n241), .A2(new_n243), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n241), .A2(KEYINPUT84), .A3(new_n243), .A4(new_n271), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT65), .B(G143), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n253), .B1(new_n277), .B2(new_n252), .ZN(new_n278));
  INV_X1    g092(.A(new_n264), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n266), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G125), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n254), .A2(new_n255), .A3(new_n260), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n270), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n261), .B2(new_n267), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n237), .B(KEYINPUT8), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n231), .A2(new_n233), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n224), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n230), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n206), .A2(new_n229), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n232), .A2(KEYINPUT85), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n232), .A2(KEYINPUT85), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n231), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n290), .B1(new_n293), .B2(new_n224), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n283), .B(new_n285), .C1(new_n289), .C2(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n228), .A2(new_n235), .A3(new_n237), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n276), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT86), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT86), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n299), .B(new_n276), .C1(new_n295), .C2(new_n296), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n275), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n188), .B1(new_n274), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n298), .A2(new_n300), .ZN(new_n303));
  INV_X1    g117(.A(new_n188), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n272), .A2(new_n273), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n275), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G478), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT15), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G122), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G116), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n218), .A2(G122), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n197), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT94), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n313), .A2(KEYINPUT14), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(KEYINPUT14), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n312), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G107), .ZN(new_n320));
  AND2_X1   g134(.A1(KEYINPUT65), .A2(G143), .ZN(new_n321));
  NOR2_X1   g135(.A1(KEYINPUT65), .A2(G143), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G128), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n258), .A2(G143), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n316), .B(new_n320), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n312), .A2(new_n313), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G107), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n314), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT13), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(KEYINPUT93), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n324), .A2(new_n326), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT93), .B(KEYINPUT13), .Z(new_n337));
  OAI21_X1  g151(.A(G134), .B1(new_n324), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n327), .B(new_n333), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT9), .B(G234), .ZN(new_n341));
  INV_X1    g155(.A(G217), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n341), .A2(new_n342), .A3(G953), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n330), .A2(new_n339), .A3(new_n343), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT71), .B(G902), .Z(new_n348));
  AOI21_X1  g162(.A(new_n310), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  AOI211_X1 g164(.A(new_n350), .B(new_n309), .C1(new_n345), .C2(new_n346), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G237), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(new_n269), .A3(G143), .A4(G214), .ZN(new_n354));
  INV_X1    g168(.A(G214), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n355), .A2(G237), .A3(G953), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n354), .B1(new_n277), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G131), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT17), .ZN(new_n359));
  INV_X1    g173(.A(G131), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n360), .B(new_n354), .C1(new_n277), .C2(new_n356), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT91), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n255), .A2(G140), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT16), .ZN(new_n368));
  OR3_X1    g182(.A1(new_n255), .A2(KEYINPUT16), .A3(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n252), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(G146), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(KEYINPUT72), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT72), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n374), .A3(new_n252), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n357), .A2(KEYINPUT17), .A3(G131), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n358), .A2(KEYINPUT91), .A3(new_n359), .A4(new_n361), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n364), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(G113), .B(G122), .Z(new_n380));
  XOR2_X1   g194(.A(KEYINPUT89), .B(G104), .Z(new_n381));
  XOR2_X1   g195(.A(new_n380), .B(new_n381), .Z(new_n382));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n366), .A2(new_n367), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(G146), .ZN(new_n385));
  XNOR2_X1  g199(.A(G125), .B(G140), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT74), .A3(new_n252), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(G146), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT18), .A2(G131), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n357), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n391), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(new_n354), .C1(new_n277), .C2(new_n356), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n379), .A2(new_n382), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n382), .B1(new_n379), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n276), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT92), .B(G475), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n364), .A2(new_n378), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n368), .A2(G146), .A3(new_n369), .ZN(new_n403));
  AOI21_X1  g217(.A(G146), .B1(new_n368), .B2(new_n369), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(new_n374), .ZN(new_n405));
  INV_X1    g219(.A(new_n375), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n377), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n396), .B(new_n382), .C1(new_n402), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT19), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n409), .B1(new_n384), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n386), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n403), .B1(new_n413), .B2(new_n252), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n358), .A2(new_n361), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n414), .A2(new_n415), .B1(new_n390), .B2(new_n395), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT90), .B1(new_n416), .B2(new_n382), .ZN(new_n417));
  INV_X1    g231(.A(new_n412), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT19), .B1(new_n386), .B2(KEYINPUT88), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n252), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n372), .ZN(new_n421));
  INV_X1    g235(.A(new_n415), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n396), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n424));
  INV_X1    g238(.A(new_n382), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n408), .A2(new_n417), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  NOR2_X1   g242(.A1(G475), .A2(G902), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n352), .B(new_n401), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G952), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G953), .ZN(new_n434));
  INV_X1    g248(.A(G234), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n353), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(new_n269), .B(new_n348), .C1(G234), .C2(G237), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(G898), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT83), .Z(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n307), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G472), .ZN(new_n446));
  INV_X1    g260(.A(new_n225), .ZN(new_n447));
  INV_X1    g261(.A(G137), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G134), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT11), .B1(new_n325), .B2(G137), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT11), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n448), .A3(G134), .ZN(new_n452));
  AOI211_X1 g266(.A(G131), .B(new_n449), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT68), .B1(new_n448), .B2(G134), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n325), .A3(G137), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n448), .A2(G134), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n360), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n254), .A2(new_n260), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n449), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n451), .B1(G134), .B2(new_n448), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n325), .A2(KEYINPUT11), .A3(G137), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT67), .A2(G131), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n449), .B1(new_n450), .B2(new_n452), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(new_n467), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n265), .B(new_n266), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n447), .A2(new_n462), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT28), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT28), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n447), .A2(new_n462), .A3(new_n472), .A4(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n280), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n265), .A2(KEYINPUT66), .A3(new_n266), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n466), .A2(new_n468), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n470), .A2(new_n467), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n245), .B1(new_n323), .B2(G146), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n252), .B1(new_n321), .B2(new_n322), .ZN(new_n485));
  INV_X1    g299(.A(new_n253), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n484), .A2(new_n259), .B1(new_n487), .B2(new_n247), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n360), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n454), .A2(new_n456), .B1(G134), .B2(new_n448), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n489), .B1(new_n360), .B2(new_n490), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT69), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n460), .B2(new_n461), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n483), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n474), .A2(new_n476), .B1(new_n495), .B2(new_n225), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n353), .A2(new_n269), .A3(G210), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT27), .Z(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT26), .B(G101), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n498), .B(new_n499), .Z(new_n500));
  AOI21_X1  g314(.A(KEYINPUT29), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n473), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n462), .A2(new_n472), .A3(KEYINPUT30), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n505), .B2(new_n225), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n501), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n462), .A2(new_n472), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n225), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n474), .B2(new_n476), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n500), .A2(KEYINPUT29), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n350), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n446), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n496), .A2(new_n500), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT31), .B1(new_n506), .B2(new_n500), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n462), .A2(new_n472), .A3(KEYINPUT30), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT69), .B1(new_n488), .B2(new_n491), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n460), .A2(new_n493), .A3(new_n461), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n280), .A2(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n479), .ZN(new_n524));
  INV_X1    g338(.A(new_n504), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n225), .B(new_n520), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n526), .A2(KEYINPUT31), .A3(new_n473), .A4(new_n500), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n518), .B1(new_n519), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(G472), .A2(G902), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n516), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n526), .A2(new_n473), .A3(new_n500), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n517), .B1(new_n534), .B2(new_n527), .ZN(new_n535));
  INV_X1    g349(.A(new_n530), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n515), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n342), .B1(new_n348), .B2(G234), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT22), .B(G137), .ZN(new_n541));
  INV_X1    g355(.A(G221), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n542), .A2(new_n435), .A3(G953), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n541), .B(new_n543), .Z(new_n544));
  NAND2_X1  g358(.A1(new_n258), .A2(G119), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n216), .A2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT24), .B(G110), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT23), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n258), .A2(KEYINPUT23), .A3(G119), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n549), .B1(G110), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n373), .A2(new_n375), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n548), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT73), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G110), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n551), .A2(new_n552), .A3(new_n559), .A4(new_n546), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT73), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n372), .A3(new_n388), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n555), .A2(KEYINPUT75), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT75), .B1(new_n555), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n544), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n544), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n555), .A2(new_n563), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n566), .A2(new_n348), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT25), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n540), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT25), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n539), .A2(G902), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n566), .A2(new_n570), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n341), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n542), .B1(new_n581), .B2(new_n276), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n207), .A2(new_n265), .A3(new_n266), .A4(new_n227), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n230), .A2(KEYINPUT10), .A3(new_n461), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n586));
  INV_X1    g400(.A(new_n260), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT78), .B1(new_n251), .B2(new_n246), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT78), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n485), .A2(new_n589), .A3(KEYINPUT1), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(G128), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n256), .A2(new_n257), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n586), .B1(new_n593), .B2(new_n290), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n585), .A2(new_n594), .B1(new_n480), .B2(new_n481), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT79), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n482), .B(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n594), .A2(new_n583), .A3(new_n584), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(G110), .B(G140), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n269), .A2(G227), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n595), .B1(new_n603), .B2(KEYINPUT80), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n598), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n488), .A2(new_n290), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n593), .B2(new_n290), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(KEYINPUT12), .A3(new_n482), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT12), .B1(new_n608), .B2(new_n482), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n598), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n604), .A2(new_n606), .B1(new_n612), .B2(new_n601), .ZN(new_n613));
  OAI21_X1  g427(.A(G469), .B1(new_n613), .B2(G902), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n603), .A2(KEYINPUT82), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n608), .A2(new_n482), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT12), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n609), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT82), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n598), .A2(new_n620), .A3(new_n602), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n594), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n583), .A2(new_n584), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n482), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n602), .B1(new_n625), .B2(new_n598), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT81), .B(G469), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n348), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n582), .B1(new_n614), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n445), .A2(new_n538), .A3(new_n580), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  INV_X1    g448(.A(new_n440), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n427), .A2(new_n429), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT20), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT95), .B(G478), .Z(new_n640));
  INV_X1    g454(.A(new_n347), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n350), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n347), .A2(KEYINPUT33), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n345), .A2(new_n644), .A3(new_n346), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n350), .A2(new_n308), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n639), .A2(new_n401), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n307), .A2(new_n442), .A3(new_n635), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n582), .ZN(new_n654));
  INV_X1    g468(.A(G469), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n604), .A2(new_n606), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n612), .A2(new_n601), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n655), .B1(new_n658), .B2(new_n276), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n603), .A2(KEYINPUT82), .B1(new_n618), .B2(new_n609), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n626), .B1(new_n660), .B2(new_n621), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n661), .A2(new_n350), .A3(new_n629), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n654), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n580), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n535), .B2(new_n350), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n529), .A2(new_n530), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n663), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n653), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT34), .B(G104), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  INV_X1    g485(.A(new_n442), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n302), .B2(new_n306), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n637), .A2(new_n638), .B1(new_n399), .B2(new_n400), .ZN(new_n674));
  INV_X1    g488(.A(new_n352), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n673), .A2(new_n635), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT35), .B(G107), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  NOR2_X1   g496(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n568), .B(new_n683), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n667), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n632), .A3(new_n445), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  NAND3_X1  g503(.A1(new_n529), .A2(new_n516), .A3(new_n530), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT32), .B1(new_n535), .B2(new_n536), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n514), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(G900), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n437), .B1(new_n438), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n677), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n692), .A2(new_n696), .A3(new_n685), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n614), .A2(new_n631), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n673), .A3(new_n654), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G128), .ZN(G30));
  XOR2_X1   g516(.A(new_n307), .B(KEYINPUT38), .Z(new_n703));
  NOR2_X1   g517(.A1(new_n674), .A2(new_n352), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n685), .A3(new_n442), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n694), .B(KEYINPUT39), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n632), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n690), .A2(new_n691), .ZN(new_n711));
  INV_X1    g525(.A(new_n500), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n506), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n509), .A2(new_n712), .A3(new_n473), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n276), .ZN(new_n715));
  OAI21_X1  g529(.A(G472), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n706), .A2(new_n709), .A3(new_n710), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n277), .ZN(G45));
  OAI21_X1  g533(.A(new_n401), .B1(new_n430), .B2(new_n431), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n648), .A2(new_n642), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n695), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n685), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n538), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT97), .B1(new_n724), .B2(new_n699), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n720), .A2(new_n721), .A3(new_n695), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n573), .A2(new_n574), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n539), .A3(new_n576), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n684), .A2(new_n577), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n692), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT97), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n700), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n725), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  AOI21_X1  g550(.A(new_n664), .B1(new_n711), .B2(new_n515), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n661), .B2(new_n350), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT98), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n631), .A3(new_n739), .A4(new_n654), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n631), .A3(new_n654), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT98), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n737), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n653), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT99), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT41), .B(G113), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NOR2_X1   g562(.A1(new_n743), .A2(new_n678), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n218), .ZN(G18));
  NAND3_X1  g564(.A1(new_n742), .A2(new_n673), .A3(new_n740), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n538), .A2(new_n441), .A3(new_n730), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n216), .ZN(G21));
  OAI22_X1  g568(.A1(new_n519), .A2(new_n528), .B1(new_n500), .B2(new_n511), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n530), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n580), .A2(new_n756), .A3(new_n665), .A4(new_n635), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n307), .A2(new_n442), .A3(new_n704), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n742), .A3(new_n758), .A4(new_n740), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT100), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  NAND2_X1  g576(.A1(new_n756), .A2(new_n665), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n685), .A3(new_n722), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n673), .A3(new_n740), .A4(new_n742), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  INV_X1    g580(.A(KEYINPUT103), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(KEYINPUT102), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n655), .A2(new_n276), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n350), .B1(new_n622), .B2(new_n627), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n630), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n604), .A2(KEYINPUT101), .A3(new_n606), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT101), .B1(new_n604), .B2(new_n606), .ZN(new_n774));
  OAI211_X1 g588(.A(G469), .B(new_n657), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n582), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n307), .A2(new_n672), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n538), .A2(new_n776), .A3(new_n580), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n722), .B1(new_n767), .B2(new_n768), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n769), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n776), .A2(new_n777), .ZN(new_n782));
  INV_X1    g596(.A(new_n769), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n737), .A3(new_n783), .A4(new_n779), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT104), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n781), .A2(new_n784), .A3(KEYINPUT104), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n360), .ZN(G33));
  NOR2_X1   g604(.A1(new_n778), .A2(new_n696), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n325), .ZN(G36));
  OAI211_X1 g606(.A(KEYINPUT45), .B(new_n657), .C1(new_n773), .C2(new_n774), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n655), .B1(new_n658), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n795), .A3(KEYINPUT105), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT105), .B1(new_n793), .B2(new_n795), .ZN(new_n798));
  OAI22_X1  g612(.A1(new_n797), .A2(new_n798), .B1(new_n655), .B2(new_n276), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n662), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI221_X1 g615(.A(KEYINPUT46), .B1(new_n655), .B2(new_n276), .C1(new_n797), .C2(new_n798), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n582), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n721), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT43), .B1(new_n648), .B2(new_n642), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n806), .A2(KEYINPUT43), .B1(new_n674), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n685), .B1(new_n666), .B2(new_n665), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(KEYINPUT44), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT44), .B1(new_n808), .B2(new_n809), .ZN(new_n811));
  INV_X1    g625(.A(new_n777), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n803), .A2(new_n707), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT107), .B(G137), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(G39));
  XNOR2_X1  g630(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n803), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT108), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT47), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n803), .A2(new_n820), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n812), .A2(new_n538), .A3(new_n580), .A4(new_n722), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n818), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G140), .ZN(G42));
  NAND2_X1  g638(.A1(new_n433), .A2(new_n269), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n808), .A2(new_n437), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n763), .A2(new_n664), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n742), .A2(new_n740), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n672), .A3(new_n703), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n828), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n829), .B1(new_n828), .B2(new_n832), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n437), .A2(new_n831), .A3(new_n777), .A4(new_n808), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n763), .A2(new_n685), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n777), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n711), .A2(new_n580), .A3(new_n437), .A4(new_n716), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n674), .A2(new_n642), .A3(new_n648), .ZN(new_n841));
  OR3_X1    g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n835), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n738), .A2(new_n631), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n582), .ZN(new_n847));
  INV_X1    g661(.A(new_n821), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n803), .A2(new_n817), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n826), .A2(new_n827), .A3(new_n777), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT113), .Z(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n844), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT51), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n828), .A2(new_n751), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n720), .A2(new_n721), .ZN(new_n857));
  OR3_X1    g671(.A1(new_n839), .A2(new_n857), .A3(new_n840), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n434), .A3(new_n858), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n859), .A2(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(KEYINPUT115), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n836), .A2(new_n737), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT48), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n862), .A2(KEYINPUT48), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n860), .A2(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n835), .A2(new_n843), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n818), .A2(new_n821), .B1(new_n582), .B2(new_n846), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n868), .B2(new_n852), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n854), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n855), .B(new_n865), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n307), .A2(new_n441), .A3(new_n444), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n663), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n737), .B2(new_n686), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n665), .A2(new_n666), .A3(new_n580), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n443), .B1(new_n302), .B2(new_n306), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n440), .B1(new_n676), .B2(new_n857), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n632), .A4(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n876), .B(new_n880), .C1(new_n652), .C2(new_n743), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n743), .A2(new_n678), .B1(new_n751), .B2(new_n752), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n837), .A2(new_n776), .A3(new_n726), .A4(new_n777), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n674), .A2(KEYINPUT110), .A3(new_n352), .A4(new_n695), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT110), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n432), .B2(new_n694), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n886), .A2(new_n888), .A3(new_n730), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n538), .A3(new_n632), .A4(new_n777), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n885), .B(new_n890), .C1(new_n778), .C2(new_n696), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n882), .A2(new_n761), .A3(new_n884), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n789), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n733), .B1(new_n732), .B2(new_n700), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n699), .A2(new_n692), .A3(KEYINPUT97), .A4(new_n731), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n701), .B(new_n765), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n685), .A2(new_n695), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT111), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n717), .A2(new_n758), .ZN(new_n901));
  INV_X1    g715(.A(new_n776), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n895), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n725), .A2(new_n734), .B1(new_n700), .B2(new_n697), .ZN(new_n905));
  OR3_X1    g719(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(KEYINPUT52), .A3(new_n906), .A4(new_n765), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n894), .A2(KEYINPUT53), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT53), .B1(new_n894), .B2(new_n908), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT112), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI211_X1 g726(.A(KEYINPUT112), .B(KEYINPUT53), .C1(new_n894), .C2(new_n908), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT54), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n787), .A2(new_n788), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n759), .B(KEYINPUT100), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n916), .A2(new_n881), .A3(new_n883), .A4(new_n891), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n908), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT53), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n881), .A2(new_n883), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n761), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n892), .A2(KEYINPUT53), .A3(new_n781), .A4(new_n784), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n908), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n920), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n914), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n825), .B1(new_n873), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n703), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n806), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n845), .A2(KEYINPUT49), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n717), .B1(KEYINPUT49), .B2(new_n845), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n580), .A2(new_n654), .A3(new_n444), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT109), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n929), .A2(new_n936), .ZN(G75));
  NOR2_X1   g751(.A1(new_n269), .A2(G952), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT119), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n241), .A2(new_n243), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n271), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT55), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n920), .A2(new_n926), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n350), .A3(new_n188), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT56), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n945), .A2(KEYINPUT116), .A3(new_n350), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT116), .ZN(new_n950));
  AOI22_X1  g764(.A1(new_n918), .A2(new_n919), .B1(new_n908), .B2(new_n925), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(new_n348), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n952), .A3(new_n188), .ZN(new_n953));
  XNOR2_X1  g767(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT118), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n944), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n955), .B2(new_n944), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n940), .B(new_n948), .C1(new_n953), .C2(new_n957), .ZN(G51));
  INV_X1    g772(.A(new_n923), .ZN(new_n959));
  INV_X1    g773(.A(new_n924), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n959), .A2(new_n908), .A3(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n910), .A2(new_n961), .A3(KEYINPUT54), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n921), .B1(new_n920), .B2(new_n926), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n770), .B(KEYINPUT57), .Z(new_n965));
  OAI21_X1  g779(.A(new_n628), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n797), .A2(new_n798), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n949), .A2(new_n952), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n938), .B1(new_n966), .B2(new_n968), .ZN(G54));
  AND2_X1   g783(.A1(KEYINPUT58), .A2(G475), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n949), .A2(new_n952), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n427), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n938), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n949), .A2(new_n952), .A3(new_n427), .A4(new_n970), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(G60));
  XOR2_X1   g789(.A(new_n646), .B(KEYINPUT120), .Z(new_n976));
  NAND2_X1  g790(.A1(G478), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT59), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n962), .B2(new_n963), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT121), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n982), .A3(new_n939), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT54), .B1(new_n910), .B2(new_n961), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n984), .B2(new_n927), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT121), .B1(new_n985), .B2(new_n940), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n976), .B1(new_n928), .B2(new_n978), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(G63));
  NAND2_X1  g803(.A1(G217), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT122), .Z(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT60), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n951), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n940), .B1(new_n993), .B2(new_n684), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT123), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n993), .B2(new_n684), .ZN(new_n996));
  OAI221_X1 g810(.A(new_n994), .B1(new_n579), .B2(new_n993), .C1(new_n996), .C2(KEYINPUT61), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n993), .A2(new_n684), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n998), .B(new_n939), .C1(new_n579), .C2(new_n993), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT61), .B1(new_n998), .B2(KEYINPUT123), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n997), .A2(new_n1001), .ZN(G66));
  NAND2_X1  g816(.A1(G224), .A2(G953), .ZN(new_n1003));
  OAI22_X1  g817(.A1(new_n923), .A2(G953), .B1(new_n439), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n941), .B1(G898), .B2(new_n269), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT124), .Z(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G69));
  INV_X1    g821(.A(new_n823), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n803), .A2(new_n737), .A3(new_n707), .A4(new_n758), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n898), .A2(new_n791), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n915), .A2(new_n814), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT126), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n915), .A2(new_n814), .A3(new_n1010), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n1014), .A3(new_n823), .A4(new_n1009), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1012), .A2(new_n1015), .A3(new_n269), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n505), .B(new_n413), .Z(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(G900), .B2(G953), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n898), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n718), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT62), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1020), .A2(KEYINPUT62), .A3(new_n718), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n676), .A2(new_n857), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT125), .Z(new_n1027));
  NOR2_X1   g841(.A1(new_n1027), .A2(new_n812), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1028), .A2(new_n737), .A3(new_n632), .A4(new_n707), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1025), .A2(new_n823), .A3(new_n814), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n269), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT127), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n1033));
  AOI22_X1  g847(.A1(new_n1031), .A2(new_n1017), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n1033), .A2(new_n1032), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n1019), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1035), .B1(new_n1019), .B2(new_n1034), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1036), .A2(new_n1037), .ZN(G72));
  NAND3_X1  g852(.A1(new_n526), .A2(new_n473), .A3(new_n712), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1012), .A2(new_n1015), .A3(new_n959), .ZN(new_n1040));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT63), .Z(new_n1042));
  AOI21_X1  g856(.A(new_n1039), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n912), .A2(new_n913), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n506), .A2(new_n500), .ZN(new_n1045));
  INV_X1    g859(.A(new_n532), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1042), .B1(new_n1030), .B2(new_n923), .ZN(new_n1049));
  AND2_X1   g863(.A1(new_n1049), .A2(new_n713), .ZN(new_n1050));
  NOR4_X1   g864(.A1(new_n1043), .A2(new_n1048), .A3(new_n1050), .A4(new_n938), .ZN(G57));
endmodule


