//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n203), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n214), .B1(new_n217), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT64), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  OAI21_X1  g0048(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n209), .A2(G33), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  OAI21_X1  g0051(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR3_X1   g0053(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G150), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n249), .B1(new_n250), .B2(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n215), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n258), .A2(new_n215), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n242), .B1(new_n208), .B2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n262), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n264), .A2(new_n265), .B1(new_n242), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G223), .A3(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n274), .A2(G77), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n276), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT66), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n271), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n285), .B2(new_n284), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(new_n271), .A3(G274), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT65), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n290), .A2(new_n271), .A3(KEYINPUT65), .A4(G274), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n271), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n290), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n296), .B1(G226), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n269), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(G179), .B2(new_n300), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(G200), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n268), .B(KEYINPUT9), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n287), .A2(G190), .A3(new_n299), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND4_X1   g0109(.A1(new_n304), .A2(new_n305), .A3(new_n308), .A4(new_n306), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g0111(.A(KEYINPUT8), .B(G58), .Z(new_n312));
  NAND2_X1  g0112(.A1(new_n208), .A2(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n314), .A2(new_n263), .B1(new_n262), .B2(new_n312), .ZN(new_n315));
  XOR2_X1   g0115(.A(new_n315), .B(KEYINPUT73), .Z(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT7), .B1(new_n274), .B2(new_n209), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n280), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G68), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT70), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n279), .A2(new_n209), .A3(new_n280), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT7), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n318), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(G68), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(G159), .B1(new_n253), .B2(new_n254), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G58), .A2(G68), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n203), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G20), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT71), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G159), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT67), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(new_n209), .A3(new_n278), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n335), .B1(new_n337), .B2(new_n252), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n209), .B1(new_n203), .B2(new_n330), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT71), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(new_n340), .A3(KEYINPUT16), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n261), .B1(new_n328), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n333), .B1(new_n329), .B2(new_n332), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT71), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n324), .A2(KEYINPUT72), .A3(new_n318), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n322), .A2(new_n348), .A3(new_n323), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(G68), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n316), .B1(new_n343), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G226), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G1698), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G223), .B2(G1698), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n357), .A2(new_n274), .B1(new_n278), .B2(new_n221), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n297), .B1(new_n298), .B2(G232), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n301), .B1(new_n359), .B2(new_n295), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n295), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(G179), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT18), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(KEYINPUT74), .A2(G190), .ZN(new_n364));
  NOR2_X1   g0164(.A1(KEYINPUT74), .A2(G190), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(new_n295), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n361), .B2(G200), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n315), .B(KEYINPUT73), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n326), .B1(new_n325), .B2(G68), .ZN(new_n370));
  AOI211_X1 g0170(.A(KEYINPUT70), .B(new_n202), .C1(new_n324), .C2(new_n318), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n259), .B1(new_n372), .B2(new_n341), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT16), .B1(new_n346), .B2(new_n350), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n368), .B(new_n369), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT18), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n361), .A2(G179), .ZN(new_n379));
  INV_X1    g0179(.A(new_n360), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n341), .B1(new_n321), .B2(new_n327), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n382), .A2(new_n374), .A3(new_n261), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n378), .B(new_n381), .C1(new_n383), .C2(new_n316), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n328), .A2(new_n342), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n353), .A3(new_n259), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n369), .A4(new_n368), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n363), .A2(new_n377), .A3(new_n384), .A4(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n311), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n255), .A2(new_n242), .ZN(new_n390));
  INV_X1    g0190(.A(G77), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n250), .A2(new_n391), .B1(new_n209), .B2(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n259), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT11), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT12), .B1(new_n262), .B2(G68), .ZN(new_n397));
  OR3_X1    g0197(.A1(new_n262), .A2(KEYINPUT12), .A3(G68), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n264), .A2(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n393), .B2(new_n394), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n293), .A2(new_n294), .B1(new_n298), .B2(G238), .ZN(new_n403));
  INV_X1    g0203(.A(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n355), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G232), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n407), .C1(new_n272), .C2(new_n273), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT69), .B1(new_n410), .B2(new_n297), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT69), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n412), .B(new_n271), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n403), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT13), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n403), .B(new_n416), .C1(new_n411), .C2(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(G169), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(G179), .A3(new_n417), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n419), .B1(new_n418), .B2(G169), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n402), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G190), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n401), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G200), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n415), .B2(new_n417), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G20), .A2(G77), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n431), .B1(new_n250), .B2(new_n432), .C1(new_n255), .C2(new_n251), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n259), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n313), .A2(G77), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n434), .B1(G77), .B2(new_n262), .C1(new_n263), .C2(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n293), .A2(new_n294), .B1(new_n298), .B2(G244), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n438));
  INV_X1    g0238(.A(G107), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n281), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n275), .A2(G232), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT68), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT68), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n275), .A2(new_n443), .A3(G232), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n437), .B1(new_n445), .B2(new_n271), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n436), .B1(new_n447), .B2(G190), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(G200), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n301), .ZN(new_n451));
  INV_X1    g0251(.A(G179), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n437), .B(new_n452), .C1(new_n445), .C2(new_n271), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n436), .A3(new_n453), .ZN(new_n454));
  AND4_X1   g0254(.A1(new_n424), .A2(new_n430), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n389), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(G257), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n458));
  OAI211_X1 g0258(.A(G250), .B(new_n404), .C1(new_n272), .C2(new_n273), .ZN(new_n459));
  INV_X1    g0259(.A(G294), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n458), .B(new_n459), .C1(new_n278), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n297), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT76), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(new_n288), .A3(KEYINPUT5), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(KEYINPUT76), .B2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n289), .A2(G1), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G264), .A3(new_n271), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n271), .A2(G274), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n462), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n427), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n468), .A2(new_n271), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n297), .A2(new_n461), .B1(new_n475), .B2(G264), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(new_n425), .A3(new_n472), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n209), .B2(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n439), .A2(KEYINPUT23), .A3(G20), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G116), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G20), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n209), .A2(KEYINPUT82), .A3(G33), .A4(G116), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n482), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n209), .B(G87), .C1(new_n272), .C2(new_n273), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(KEYINPUT81), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n281), .A2(new_n491), .A3(new_n209), .A4(G87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT24), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT24), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n487), .A2(new_n495), .A3(new_n490), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n259), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n261), .B(new_n262), .C1(G1), .C2(new_n278), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT25), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n262), .B2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n262), .A2(new_n500), .A3(G107), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n499), .A2(new_n439), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n478), .A2(new_n498), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n473), .A2(G169), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n476), .A2(G179), .A3(new_n472), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT83), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n476), .A2(KEYINPUT83), .A3(G179), .A4(new_n472), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n261), .B1(new_n494), .B2(new_n496), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n506), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(G244), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n515));
  OAI211_X1 g0315(.A(G238), .B(new_n404), .C1(new_n272), .C2(new_n273), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n484), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n297), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n467), .A2(new_n222), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n471), .A2(new_n467), .B1(new_n519), .B2(new_n271), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT78), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n452), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT19), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n209), .B1(new_n409), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(G87), .B2(new_n206), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n209), .B(G68), .C1(new_n272), .C2(new_n273), .ZN(new_n528));
  INV_X1    g0328(.A(G97), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n525), .B1(new_n250), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT79), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n527), .A2(KEYINPUT79), .A3(new_n528), .A4(new_n530), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n259), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n432), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n262), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n499), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n536), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT78), .B1(new_n521), .B2(G179), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n521), .A2(new_n301), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n524), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n261), .B1(new_n531), .B2(new_n532), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n537), .B1(new_n545), .B2(new_n534), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n539), .A2(G87), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n521), .A2(G190), .ZN(new_n548));
  AOI21_X1  g0348(.A(G200), .B1(new_n518), .B2(new_n520), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n514), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G244), .B(new_n404), .C1(new_n272), .C2(new_n273), .ZN(new_n553));
  XOR2_X1   g0353(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n558), .C1(new_n553), .C2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n297), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n468), .A2(G257), .A3(new_n271), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n472), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n301), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n472), .A2(new_n562), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n404), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n555), .A2(new_n567), .A3(new_n557), .A4(new_n558), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n566), .B1(new_n297), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n452), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n347), .A2(G107), .A3(new_n349), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n439), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  XOR2_X1   g0372(.A(G97), .B(G107), .Z(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(KEYINPUT6), .ZN(new_n574));
  INV_X1    g0374(.A(new_n255), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n574), .A2(G20), .B1(new_n575), .B2(G77), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n261), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n262), .A2(G97), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n539), .B2(G97), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n565), .B(new_n570), .C1(new_n577), .C2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT77), .B1(new_n569), .B2(new_n427), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT77), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n564), .A2(new_n583), .A3(G200), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n569), .A2(G190), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n571), .A2(new_n576), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n259), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n588), .A3(new_n579), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n581), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(G20), .B1(G33), .B2(G283), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(G33), .B2(new_n529), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G116), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n258), .A2(new_n215), .B1(G20), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n591), .B(KEYINPUT80), .C1(G33), .C2(new_n529), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n594), .A2(new_n596), .A3(KEYINPUT20), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n499), .A2(G116), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n262), .A2(new_n595), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n600), .A2(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(G264), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n606));
  OAI211_X1 g0406(.A(G257), .B(new_n404), .C1(new_n272), .C2(new_n273), .ZN(new_n607));
  INV_X1    g0407(.A(G303), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n606), .B(new_n607), .C1(new_n608), .C2(new_n281), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n297), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n468), .A2(G270), .A3(new_n271), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n472), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n605), .A2(KEYINPUT21), .A3(G169), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(G169), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n604), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n472), .A2(new_n611), .ZN(new_n617));
  INV_X1    g0417(.A(new_n366), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(new_n610), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n610), .A2(new_n472), .A3(new_n611), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n604), .B(new_n619), .C1(new_n620), .C2(new_n427), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n617), .A2(G179), .A3(new_n610), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n605), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n613), .A2(new_n616), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n590), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n457), .A2(new_n552), .A3(new_n625), .ZN(G372));
  OR2_X1    g0426(.A1(new_n309), .A2(new_n310), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n377), .A2(new_n387), .ZN(new_n628));
  INV_X1    g0428(.A(new_n454), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n430), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(new_n424), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n363), .A2(new_n384), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n627), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n303), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n522), .A2(new_n452), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n541), .A2(new_n635), .A3(new_n543), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n585), .A2(new_n589), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n636), .A2(new_n550), .A3(KEYINPUT84), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT84), .B1(new_n636), .B2(new_n550), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n637), .B(new_n581), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n513), .A2(new_n510), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n613), .A2(new_n616), .A3(new_n623), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n506), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n636), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n551), .A2(new_n645), .A3(new_n581), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n581), .A2(KEYINPUT85), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n588), .A2(new_n579), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT85), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n565), .A4(new_n570), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n647), .B(new_n650), .C1(new_n638), .C2(new_n639), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n651), .B2(new_n645), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n634), .B1(new_n457), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT86), .ZN(G369));
  INV_X1    g0455(.A(G13), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n656), .A2(G1), .A3(G20), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(G213), .B1(new_n658), .B2(KEYINPUT27), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT27), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n657), .A2(KEYINPUT87), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT87), .B1(new_n657), .B2(new_n660), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n604), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n624), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n642), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G330), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n665), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n512), .B2(new_n504), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  INV_X1    g0475(.A(new_n514), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n641), .A2(new_n673), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT89), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n641), .A2(new_n665), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n642), .A2(new_n665), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(new_n675), .A3(new_n676), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n212), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n218), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n653), .A2(new_n693), .A3(new_n665), .ZN(new_n694));
  INV_X1    g0494(.A(new_n636), .ZN(new_n695));
  INV_X1    g0495(.A(new_n639), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n636), .A2(new_n550), .A3(KEYINPUT84), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n590), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n642), .A2(new_n506), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n513), .A2(new_n510), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n695), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n551), .A2(KEYINPUT26), .A3(new_n581), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n651), .B2(KEYINPUT26), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n673), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n694), .B1(new_n693), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n552), .A2(new_n625), .A3(new_n665), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n569), .A2(new_n522), .A3(new_n476), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n620), .A2(G179), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n612), .A2(new_n452), .A3(new_n521), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n476), .A2(new_n472), .B1(new_n561), .B2(new_n563), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND4_X1   g0515(.A1(new_n518), .A2(new_n462), .A3(new_n520), .A4(new_n469), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n622), .A2(new_n716), .A3(KEYINPUT30), .A4(new_n569), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n673), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n622), .A2(new_n716), .A3(new_n569), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n722), .A2(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n665), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT31), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n708), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n707), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n692), .B1(new_n729), .B2(G1), .ZN(G364));
  NOR2_X1   g0530(.A1(new_n656), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n208), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n687), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n686), .A2(new_n274), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n736), .A2(G355), .B1(new_n595), .B2(new_n686), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n686), .A2(new_n281), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G45), .B2(new_n218), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n247), .A2(new_n289), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT91), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n215), .B1(G20), .B2(new_n301), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n735), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n425), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n209), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n274), .B1(new_n751), .B2(new_n460), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n209), .A2(new_n452), .A3(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n618), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n209), .A2(new_n425), .A3(new_n427), .A4(G179), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n755), .A2(G322), .B1(G303), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G311), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n753), .A2(new_n425), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n209), .A2(new_n452), .A3(new_n427), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT92), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT92), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n762), .A2(new_n618), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT95), .Z(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT96), .B(G326), .Z(new_n767));
  AOI211_X1 g0567(.A(new_n752), .B(new_n760), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n452), .A2(new_n425), .A3(new_n427), .A4(G20), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n209), .A2(new_n427), .A3(G179), .A4(G190), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n773), .A2(G329), .B1(G283), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n762), .A2(new_n425), .A3(new_n763), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT94), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n762), .A2(KEYINPUT94), .A3(new_n425), .A4(new_n763), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(KEYINPUT33), .B(G317), .Z(new_n782));
  OAI211_X1 g0582(.A(new_n768), .B(new_n776), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n781), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G68), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n281), .B1(new_n754), .B2(new_n201), .ZN(new_n786));
  INV_X1    g0586(.A(new_n756), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n787), .A2(new_n221), .B1(new_n391), .B2(new_n759), .ZN(new_n788));
  INV_X1    g0588(.A(new_n774), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n439), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n751), .A2(new_n529), .ZN(new_n791));
  NOR4_X1   g0591(.A1(new_n786), .A2(new_n788), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n773), .A2(G159), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT32), .ZN(new_n794));
  INV_X1    g0594(.A(new_n764), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(KEYINPUT32), .B1(new_n795), .B2(G50), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n785), .A2(new_n792), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n783), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n747), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n749), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT98), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n669), .B2(new_n745), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n670), .A2(new_n671), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT90), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n804), .B(new_n735), .C1(new_n671), .C2(new_n670), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  OAI221_X1 g0607(.A(new_n274), .B1(new_n529), .B2(new_n751), .C1(new_n772), .C2(new_n758), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n756), .A2(G107), .B1(new_n774), .B2(G87), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n809), .B1(new_n595), .B2(new_n759), .C1(new_n460), .C2(new_n754), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n808), .B(new_n810), .C1(G303), .C2(new_n795), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n781), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT100), .ZN(new_n814));
  INV_X1    g0614(.A(new_n759), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n755), .A2(G143), .B1(G159), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n817), .B2(new_n764), .C1(new_n781), .C2(new_n256), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n274), .B1(new_n774), .B2(G68), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n822), .B1(new_n201), .B2(new_n751), .C1(new_n242), .C2(new_n787), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G132), .B2(new_n773), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n747), .B1(new_n814), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n747), .A2(new_n742), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT99), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n735), .B1(new_n829), .B2(new_n391), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT101), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n629), .A2(new_n665), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n448), .A2(new_n449), .B1(new_n436), .B2(new_n673), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n629), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n833), .B(new_n834), .C1(new_n742), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n653), .A2(new_n665), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n837), .ZN(new_n840));
  INV_X1    g0640(.A(new_n837), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n665), .B(new_n841), .C1(new_n644), .C2(new_n652), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n843), .A2(new_n727), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n734), .B1(new_n843), .B2(new_n727), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  NOR2_X1   g0647(.A1(new_n731), .A2(new_n208), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n346), .B1(new_n370), .B2(new_n371), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n352), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n315), .B1(new_n343), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n664), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n375), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n851), .A2(new_n362), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n383), .A2(new_n316), .B1(new_n381), .B2(new_n664), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n375), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n851), .A2(new_n852), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n388), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n861), .A3(KEYINPUT38), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT39), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n354), .A2(new_n852), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n857), .B1(new_n856), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n375), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n386), .A2(new_n369), .B1(new_n362), .B2(new_n852), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n388), .A2(new_n865), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n869), .B2(KEYINPUT104), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n868), .B2(new_n869), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT105), .B1(new_n864), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n388), .A2(new_n865), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n867), .A2(new_n870), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT105), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(new_n863), .A4(new_n862), .ZN(new_n882));
  INV_X1    g0682(.A(new_n862), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n859), .B2(new_n861), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT39), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n875), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n417), .ZN(new_n887));
  NOR2_X1   g0687(.A1(G226), .A2(G1698), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n406), .B2(G1698), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n889), .A2(new_n281), .B1(G33), .B2(G97), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n412), .B1(new_n890), .B2(new_n271), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n410), .A2(KEYINPUT69), .A3(new_n297), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n416), .B1(new_n893), .B2(new_n403), .ZN(new_n894));
  OAI21_X1  g0694(.A(G169), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT14), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n421), .A3(new_n420), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n402), .A3(new_n665), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n886), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n402), .A2(new_n673), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n424), .A2(new_n430), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n402), .B(new_n673), .C1(new_n897), .C2(new_n429), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n842), .B2(new_n835), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n859), .A2(new_n861), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n879), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n862), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n906), .A2(new_n909), .B1(new_n632), .B2(new_n852), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n900), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n634), .B1(new_n706), .B2(new_n457), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n911), .B(new_n912), .Z(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT106), .B1(new_n724), .B2(KEYINPUT31), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT106), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n719), .A2(new_n915), .A3(new_n720), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n708), .A2(new_n914), .A3(new_n725), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n837), .B1(new_n902), .B2(new_n903), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n917), .B(new_n918), .C1(new_n883), .C2(new_n884), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n880), .A2(new_n862), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n918), .A2(KEYINPUT40), .A3(new_n917), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n919), .A2(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n457), .A2(new_n917), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(new_n457), .A3(new_n917), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(G330), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n848), .B1(new_n913), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n913), .B2(new_n927), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT102), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n243), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n242), .A2(KEYINPUT102), .A3(G68), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n330), .A2(G77), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n931), .B(new_n932), .C1(new_n218), .C2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(G1), .A3(new_n656), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT103), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n595), .B(new_n217), .C1(new_n574), .C2(KEYINPUT35), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(KEYINPUT35), .B2(new_n574), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT36), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n938), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n929), .A2(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n648), .A2(new_n673), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n637), .A2(new_n581), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n581), .A2(new_n665), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n684), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n581), .B1(new_n944), .B2(new_n700), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n949), .A2(KEYINPUT42), .B1(new_n665), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n546), .A2(new_n547), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n673), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n638), .B2(new_n639), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n636), .B2(new_n954), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n950), .A2(new_n952), .B1(KEYINPUT43), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n680), .B(KEYINPUT89), .Z(new_n959));
  INV_X1    g0759(.A(KEYINPUT107), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n960), .A3(new_n946), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT107), .B1(new_n681), .B2(new_n947), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n958), .A3(new_n962), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n957), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n961), .A2(new_n958), .A3(new_n962), .ZN(new_n967));
  INV_X1    g0767(.A(new_n957), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n967), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n687), .B(KEYINPUT41), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n684), .A2(new_n682), .ZN(new_n972));
  OR3_X1    g0772(.A1(new_n972), .A2(new_n947), .A3(KEYINPUT108), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT108), .B1(new_n972), .B2(new_n947), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n946), .B1(new_n684), .B2(new_n682), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT44), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(new_n959), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n684), .B1(new_n679), .B2(new_n683), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n672), .A2(KEYINPUT110), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n672), .A2(KEYINPUT110), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n985), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n728), .A2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n981), .A2(new_n983), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n984), .B(new_n990), .C1(new_n991), .C2(new_n959), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n971), .B1(new_n992), .B2(new_n729), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n970), .B1(new_n993), .B2(new_n733), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n748), .B1(new_n212), .B2(new_n432), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n738), .A2(new_n232), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n734), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(G317), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n274), .B1(new_n529), .B2(new_n789), .C1(new_n772), .C2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n787), .A2(new_n595), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT46), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT111), .B1(new_n1000), .B2(KEYINPUT46), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n1000), .A2(KEYINPUT111), .A3(KEYINPUT46), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n751), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n755), .A2(G303), .B1(G107), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n812), .B2(new_n759), .ZN(new_n1007));
  NOR4_X1   g0807(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1007), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n460), .B2(new_n781), .C1(new_n758), .C2(new_n765), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n784), .A2(G159), .B1(G50), .B2(new_n815), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n756), .A2(G58), .B1(new_n774), .B2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n256), .B2(new_n754), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n281), .B1(new_n202), .B2(new_n751), .C1(new_n772), .C2(new_n817), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n766), .C2(G143), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1009), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n997), .B1(new_n1019), .B2(new_n747), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n745), .B2(new_n956), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n994), .A2(new_n1021), .ZN(G387));
  NOR2_X1   g0822(.A1(new_n989), .A2(new_n732), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n754), .A2(new_n998), .B1(new_n608), .B2(new_n759), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT116), .Z(new_n1025));
  INV_X1    g0825(.A(G322), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1025), .B1(new_n758), .B2(new_n781), .C1(new_n765), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1005), .A2(G283), .B1(G294), .B2(new_n756), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n274), .B1(new_n789), .B2(new_n595), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n773), .B2(new_n767), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n756), .A2(G77), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n772), .B2(new_n256), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT114), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n281), .B1(new_n529), .B2(new_n789), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT115), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G68), .A2(new_n815), .B1(new_n1005), .B2(new_n536), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n242), .B2(new_n754), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G159), .B2(new_n795), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1044), .B(new_n1047), .C1(new_n251), .C2(new_n781), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n799), .B1(new_n1038), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n251), .A2(G50), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT50), .Z(new_n1051));
  OAI211_X1 g0851(.A(new_n689), .B(new_n289), .C1(new_n202), .C2(new_n391), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n738), .B1(new_n1051), .B2(new_n1052), .C1(new_n237), .C2(new_n289), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n212), .A2(new_n281), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1053), .B1(G107), .B2(new_n212), .C1(new_n689), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT113), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n746), .B(new_n747), .C1(new_n1056), .C2(KEYINPUT113), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n735), .B(new_n1049), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT117), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n679), .A2(new_n745), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1023), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n990), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n728), .A2(new_n989), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n687), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1064), .A2(new_n1067), .ZN(G393));
  NOR2_X1   g0868(.A1(new_n981), .A2(new_n959), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n982), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n992), .B(new_n687), .C1(new_n990), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n947), .A2(new_n746), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n748), .B1(new_n529), .B2(new_n212), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n241), .A2(new_n686), .A3(new_n281), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n734), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n787), .A2(new_n812), .B1(new_n460), .B2(new_n759), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n274), .B1(new_n439), .B2(new_n789), .C1(new_n772), .C2(new_n1026), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G116), .C2(new_n1005), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n764), .A2(new_n998), .B1(new_n754), .B2(new_n758), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n608), .C2(new_n781), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n281), .B1(new_n789), .B2(new_n221), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n751), .A2(new_n391), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G68), .B2(new_n756), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n251), .B2(new_n759), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1082), .B(new_n1085), .C1(G143), .C2(new_n773), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n781), .B2(new_n242), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n764), .A2(new_n256), .B1(new_n754), .B2(new_n335), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1081), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1075), .B1(new_n1091), .B2(new_n747), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1070), .A2(new_n733), .B1(new_n1072), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1071), .A2(new_n1093), .ZN(G390));
  NAND2_X1  g0894(.A1(new_n436), .A2(new_n673), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n629), .B1(new_n450), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n705), .A2(new_n1097), .B1(new_n629), .B2(new_n665), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n898), .B(new_n921), .C1(new_n1098), .C2(new_n905), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n906), .A2(new_n899), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n886), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n837), .A2(new_n671), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n917), .A2(new_n904), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n726), .A2(new_n1102), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1106), .A2(new_n905), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1099), .B(new_n1108), .C1(new_n886), .C2(new_n1100), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1105), .A2(KEYINPUT119), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT119), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1101), .A2(new_n1111), .A3(new_n1104), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n389), .A2(G330), .A3(new_n455), .A4(new_n917), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT120), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n904), .B1(new_n917), .B2(new_n1102), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1116), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1106), .A2(new_n905), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1118), .A2(new_n1103), .B1(new_n835), .B2(new_n842), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n912), .B(new_n1114), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1110), .A2(new_n1112), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1110), .A2(KEYINPUT121), .A3(new_n1112), .A4(new_n1120), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1120), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n688), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n733), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n734), .B1(new_n828), .B2(new_n312), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n274), .B1(new_n221), .B2(new_n787), .C1(new_n772), .C2(new_n460), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n789), .A2(new_n202), .B1(new_n751), .B2(new_n391), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n754), .A2(new_n595), .B1(new_n529), .B2(new_n759), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n812), .B2(new_n764), .C1(new_n439), .C2(new_n781), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n787), .A2(new_n256), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT53), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n274), .B(new_n1139), .C1(G50), .C2(new_n774), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n751), .A2(new_n335), .ZN(new_n1141));
  INV_X1    g0941(.A(G132), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n754), .A2(new_n1142), .B1(new_n759), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1141), .B(new_n1144), .C1(new_n795), .C2(G128), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n773), .A2(G125), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1140), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n781), .A2(new_n817), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1136), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1131), .B1(new_n1149), .B2(new_n747), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n886), .B2(new_n743), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1130), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1129), .A2(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(KEYINPUT57), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n912), .A2(new_n1114), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n921), .A2(new_n922), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n918), .A2(new_n917), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n862), .B2(new_n908), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(G330), .C1(new_n1160), .C2(KEYINPUT40), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT124), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n923), .A2(KEYINPUT124), .A3(G330), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n269), .A2(new_n852), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n311), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n311), .A2(new_n1165), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1163), .A2(new_n1164), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1173), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1175), .A2(new_n923), .A3(KEYINPUT124), .A4(G330), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n911), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n911), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1174), .A2(new_n1176), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1155), .B1(new_n1157), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1156), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1174), .A2(new_n1179), .A3(new_n1176), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1179), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n1155), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1182), .A2(new_n1189), .A3(new_n687), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1175), .A2(new_n742), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n734), .B1(new_n828), .B2(G50), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n789), .A2(new_n201), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n281), .A2(G41), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1039), .A2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G283), .C2(new_n773), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT122), .Z(new_n1198));
  AOI22_X1  g0998(.A1(new_n536), .A2(new_n815), .B1(new_n1005), .B2(G68), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n439), .B2(new_n754), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G116), .B2(new_n795), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(new_n529), .C2(new_n781), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT123), .Z(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(G33), .A2(G41), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1195), .A2(G50), .A3(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n755), .A2(G128), .B1(G137), .B2(new_n815), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n256), .B2(new_n751), .C1(new_n787), .C2(new_n1143), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G125), .B2(new_n795), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1142), .B2(new_n781), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1212));
  INV_X1    g1012(.A(G124), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1206), .B1(new_n335), .B2(new_n789), .C1(new_n772), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1211), .B2(KEYINPUT59), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1207), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1204), .A2(new_n1205), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1193), .B1(new_n1217), .B2(new_n747), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1191), .A2(new_n733), .B1(new_n1192), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1190), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n905), .A2(new_n742), .ZN(new_n1221));
  INV_X1    g1021(.A(G128), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n281), .B1(new_n201), .B2(new_n789), .C1(new_n772), .C2(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n754), .A2(new_n817), .B1(new_n256), .B2(new_n759), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n787), .A2(new_n335), .B1(new_n242), .B2(new_n751), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n1142), .B2(new_n764), .C1(new_n781), .C2(new_n1143), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n274), .B1(new_n789), .B2(new_n391), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n764), .A2(new_n460), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1229), .B2(new_n1228), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n787), .A2(new_n529), .B1(new_n439), .B2(new_n759), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n754), .A2(new_n812), .B1(new_n432), .B2(new_n751), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(G303), .C2(new_n773), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1231), .B(new_n1234), .C1(new_n595), .C2(new_n781), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n799), .B1(new_n1227), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n735), .B(new_n1236), .C1(new_n202), .C2(new_n829), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1221), .A2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1238), .B1(new_n1239), .B2(new_n732), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1127), .A2(new_n971), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1156), .A2(new_n1239), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G381));
  INV_X1    g1044(.A(G390), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(G393), .A2(G396), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1245), .A2(new_n846), .A3(new_n1243), .A4(new_n1246), .ZN(new_n1247));
  OR4_X1    g1047(.A1(G387), .A2(G375), .A3(new_n1247), .A4(G378), .ZN(G407));
  AOI21_X1  g1048(.A(new_n1152), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1249));
  INV_X1    g1049(.A(G343), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(G213), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G375), .C2(new_n1253), .ZN(G409));
  NAND2_X1  g1054(.A1(G387), .A2(new_n1245), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(G393), .B(new_n806), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n994), .A2(new_n1021), .A3(G390), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1190), .A2(G378), .A3(new_n1219), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1219), .B1(new_n1263), .B2(new_n971), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1249), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1252), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1156), .A2(new_n1239), .A3(KEYINPUT60), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1267), .A2(new_n687), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1120), .A2(KEYINPUT60), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1242), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1240), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G384), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n846), .B(new_n1240), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1252), .A2(G2897), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1273), .A2(new_n1274), .A3(KEYINPUT126), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1240), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(G384), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT126), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1276), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1261), .B1(new_n1266), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1266), .B2(new_n1278), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1252), .B(new_n1282), .C1(new_n1262), .C2(new_n1265), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1286), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1260), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1278), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1292), .B(new_n1261), .C1(new_n1266), .C2(new_n1284), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1260), .B1(new_n1289), .B2(KEYINPUT63), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(KEYINPUT127), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1266), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1284), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1266), .A2(new_n1278), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT62), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1301), .A3(new_n1290), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1260), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1300), .A2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1299), .A2(new_n1307), .A3(new_n1260), .A4(new_n1292), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1304), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1296), .A2(new_n1309), .ZN(G405));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1249), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1262), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(new_n1282), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1313), .B(new_n1260), .ZN(G402));
endmodule


