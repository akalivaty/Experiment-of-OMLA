

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786;

  XNOR2_X1 U373 ( .A(n424), .B(n423), .ZN(n746) );
  NOR2_X1 U374 ( .A1(n729), .A2(n490), .ZN(n652) );
  XNOR2_X1 U375 ( .A(n386), .B(KEYINPUT109), .ZN(n651) );
  NOR2_X1 U376 ( .A1(n635), .A2(n700), .ZN(n618) );
  XNOR2_X1 U377 ( .A(n484), .B(n507), .ZN(n742) );
  OR2_X1 U378 ( .A1(n607), .A2(n358), .ZN(n475) );
  XNOR2_X1 U379 ( .A(n585), .B(n549), .ZN(n769) );
  XNOR2_X2 U380 ( .A(n521), .B(n520), .ZN(n782) );
  NAND2_X1 U381 ( .A1(n355), .A2(n382), .ZN(n387) );
  NAND2_X1 U382 ( .A1(n380), .A2(n381), .ZN(n355) );
  INV_X1 U383 ( .A(n637), .ZN(n381) );
  INV_X1 U384 ( .A(G953), .ZN(n774) );
  XNOR2_X2 U385 ( .A(n526), .B(KEYINPUT104), .ZN(n400) );
  AND2_X2 U386 ( .A1(n414), .A2(n419), .ZN(n416) );
  XNOR2_X2 U387 ( .A(KEYINPUT68), .B(G131), .ZN(n580) );
  OR2_X2 U388 ( .A1(n772), .A2(G101), .ZN(n546) );
  AND2_X2 U389 ( .A1(n435), .A2(n456), .ZN(n628) );
  XNOR2_X2 U390 ( .A(n491), .B(n650), .ZN(n729) );
  NOR2_X2 U391 ( .A1(n718), .A2(n716), .ZN(n491) );
  INV_X2 U392 ( .A(G128), .ZN(n544) );
  XNOR2_X1 U393 ( .A(n484), .B(n548), .ZN(n607) );
  XNOR2_X2 U394 ( .A(n592), .B(KEYINPUT4), .ZN(n772) );
  XNOR2_X2 U395 ( .A(n544), .B(G143), .ZN(n592) );
  INV_X2 U396 ( .A(G125), .ZN(n510) );
  INV_X1 U397 ( .A(KEYINPUT32), .ZN(n528) );
  XNOR2_X1 U398 ( .A(n652), .B(n513), .ZN(n378) );
  XNOR2_X1 U399 ( .A(n667), .B(KEYINPUT108), .ZN(n783) );
  NAND2_X1 U400 ( .A1(n546), .A2(n545), .ZN(n377) );
  XNOR2_X1 U401 ( .A(G134), .B(n580), .ZN(n770) );
  XNOR2_X1 U402 ( .A(n524), .B(G110), .ZN(n762) );
  XNOR2_X1 U403 ( .A(n373), .B(n370), .ZN(n356) );
  XNOR2_X1 U404 ( .A(n373), .B(n370), .ZN(n735) );
  OR2_X2 U405 ( .A1(n748), .A2(G902), .ZN(n431) );
  NOR2_X2 U406 ( .A1(n742), .A2(G902), .ZN(n406) );
  INV_X1 U407 ( .A(KEYINPUT30), .ZN(n472) );
  XNOR2_X1 U408 ( .A(n437), .B(n502), .ZN(n397) );
  INV_X1 U409 ( .A(KEYINPUT48), .ZN(n502) );
  NOR2_X1 U410 ( .A1(n428), .A2(n427), .ZN(n426) );
  XNOR2_X1 U411 ( .A(n425), .B(KEYINPUT66), .ZN(n444) );
  NOR2_X1 U412 ( .A1(n782), .A2(KEYINPUT44), .ZN(n425) );
  XNOR2_X1 U413 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n553) );
  XNOR2_X1 U414 ( .A(n485), .B(n533), .ZN(n585) );
  INV_X1 U415 ( .A(KEYINPUT10), .ZN(n533) );
  AND2_X1 U416 ( .A1(n418), .A2(n417), .ZN(n414) );
  INV_X1 U417 ( .A(n670), .ZN(n417) );
  INV_X1 U418 ( .A(G469), .ZN(n405) );
  XNOR2_X1 U419 ( .A(n762), .B(KEYINPUT73), .ZN(n606) );
  XNOR2_X1 U420 ( .A(n770), .B(G146), .ZN(n547) );
  NAND2_X1 U421 ( .A1(n487), .A2(n529), .ZN(n428) );
  XNOR2_X1 U422 ( .A(n661), .B(KEYINPUT78), .ZN(n487) );
  INV_X1 U423 ( .A(KEYINPUT102), .ZN(n505) );
  NOR2_X1 U424 ( .A1(G953), .A2(G237), .ZN(n573) );
  XNOR2_X1 U425 ( .A(n557), .B(KEYINPUT25), .ZN(n534) );
  XNOR2_X1 U426 ( .A(n508), .B(KEYINPUT77), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n509), .B(KEYINPUT76), .ZN(n508) );
  INV_X1 U428 ( .A(KEYINPUT18), .ZN(n509) );
  XNOR2_X1 U429 ( .A(n560), .B(n606), .ZN(n374) );
  XOR2_X1 U430 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n559) );
  NAND2_X1 U431 ( .A1(n714), .A2(n713), .ZN(n718) );
  NAND2_X1 U432 ( .A1(n469), .A2(n468), .ZN(n467) );
  AND2_X1 U433 ( .A1(n473), .A2(n357), .ZN(n470) );
  NAND2_X1 U434 ( .A1(n474), .A2(n477), .ZN(n473) );
  AND2_X1 U435 ( .A1(n475), .A2(KEYINPUT30), .ZN(n474) );
  NAND2_X1 U436 ( .A1(n477), .A2(n475), .ZN(n704) );
  XNOR2_X1 U437 ( .A(n704), .B(n518), .ZN(n658) );
  INV_X1 U438 ( .A(KEYINPUT6), .ZN(n518) );
  XNOR2_X1 U439 ( .A(n503), .B(n457), .ZN(n435) );
  INV_X1 U440 ( .A(KEYINPUT22), .ZN(n457) );
  NAND2_X2 U441 ( .A1(n390), .A2(n388), .ZN(n773) );
  NAND2_X1 U442 ( .A1(n389), .A2(n393), .ZN(n388) );
  AND2_X1 U443 ( .A1(n395), .A2(n391), .ZN(n390) );
  NAND2_X1 U444 ( .A1(n402), .A2(n403), .ZN(n376) );
  INV_X1 U445 ( .A(KEYINPUT45), .ZN(n458) );
  XOR2_X1 U446 ( .A(KEYINPUT90), .B(KEYINPUT72), .Z(n551) );
  XNOR2_X1 U447 ( .A(G119), .B(KEYINPUT79), .ZN(n550) );
  XNOR2_X1 U448 ( .A(n450), .B(n449), .ZN(n448) );
  XNOR2_X1 U449 ( .A(G128), .B(G110), .ZN(n449) );
  XNOR2_X1 U450 ( .A(n451), .B(KEYINPUT23), .ZN(n450) );
  XNOR2_X1 U451 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n451) );
  NOR2_X1 U452 ( .A1(n654), .A2(n653), .ZN(n655) );
  AND2_X1 U453 ( .A1(n453), .A2(n452), .ZN(n662) );
  NOR2_X1 U454 ( .A1(n690), .A2(n565), .ZN(n452) );
  XNOR2_X1 U455 ( .A(n455), .B(n454), .ZN(n453) );
  INV_X1 U456 ( .A(KEYINPUT106), .ZN(n454) );
  AND2_X1 U457 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U458 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n523) );
  XNOR2_X1 U459 ( .A(n596), .B(n407), .ZN(n747) );
  XNOR2_X1 U460 ( .A(n597), .B(n595), .ZN(n407) );
  XNOR2_X1 U461 ( .A(n605), .B(n606), .ZN(n507) );
  XNOR2_X1 U462 ( .A(n462), .B(n603), .ZN(n605) );
  XNOR2_X1 U463 ( .A(n604), .B(n463), .ZN(n462) );
  XNOR2_X1 U464 ( .A(KEYINPUT20), .B(KEYINPUT92), .ZN(n555) );
  NAND2_X1 U465 ( .A1(n713), .A2(n472), .ZN(n471) );
  INV_X1 U466 ( .A(KEYINPUT28), .ZN(n385) );
  OR2_X1 U467 ( .A1(G237), .A2(G902), .ZN(n564) );
  XNOR2_X1 U468 ( .A(G902), .B(KEYINPUT15), .ZN(n670) );
  INV_X1 U469 ( .A(G902), .ZN(n476) );
  AND2_X1 U470 ( .A1(n479), .A2(n478), .ZN(n477) );
  NAND2_X1 U471 ( .A1(G472), .A2(G902), .ZN(n478) );
  INV_X1 U472 ( .A(KEYINPUT5), .ZN(n539) );
  INV_X1 U473 ( .A(KEYINPUT81), .ZN(n393) );
  AND2_X1 U474 ( .A1(n392), .A2(n785), .ZN(n391) );
  NAND2_X1 U475 ( .A1(n394), .A2(n393), .ZN(n392) );
  INV_X1 U476 ( .A(n783), .ZN(n394) );
  INV_X1 U477 ( .A(KEYINPUT71), .ZN(n497) );
  INV_X1 U478 ( .A(n400), .ZN(n511) );
  INV_X1 U479 ( .A(KEYINPUT84), .ZN(n459) );
  XOR2_X1 U480 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n575) );
  XNOR2_X1 U481 ( .A(G113), .B(G143), .ZN(n576) );
  XOR2_X1 U482 ( .A(G140), .B(KEYINPUT12), .Z(n577) );
  XOR2_X1 U483 ( .A(G122), .B(G104), .Z(n581) );
  INV_X1 U484 ( .A(KEYINPUT64), .ZN(n423) );
  NAND2_X1 U485 ( .A1(G234), .A2(G237), .ZN(n566) );
  XOR2_X1 U486 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n567) );
  NAND2_X1 U487 ( .A1(n773), .A2(n422), .ZN(n418) );
  INV_X1 U488 ( .A(KEYINPUT38), .ZN(n649) );
  NAND2_X1 U489 ( .A1(n658), .A2(n517), .ZN(n455) );
  XNOR2_X1 U490 ( .A(n614), .B(n364), .ZN(n493) );
  INV_X1 U491 ( .A(KEYINPUT105), .ZN(n612) );
  NAND2_X1 U492 ( .A1(n659), .A2(n385), .ZN(n383) );
  NAND2_X1 U493 ( .A1(n637), .A2(n385), .ZN(n384) );
  NOR2_X1 U494 ( .A1(n659), .A2(n385), .ZN(n380) );
  INV_X1 U495 ( .A(G107), .ZN(n524) );
  XNOR2_X1 U496 ( .A(G116), .B(G107), .ZN(n408) );
  XNOR2_X1 U497 ( .A(G122), .B(KEYINPUT7), .ZN(n590) );
  XOR2_X1 U498 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n591) );
  INV_X1 U499 ( .A(G104), .ZN(n463) );
  XNOR2_X1 U500 ( .A(n377), .B(n371), .ZN(n370) );
  XNOR2_X1 U501 ( .A(n485), .B(n372), .ZN(n371) );
  NAND2_X1 U502 ( .A1(n421), .A2(n420), .ZN(n415) );
  NOR2_X1 U503 ( .A1(n773), .A2(n422), .ZN(n421) );
  INV_X1 U504 ( .A(n404), .ZN(n486) );
  BUF_X1 U505 ( .A(n493), .Z(n404) );
  NAND2_X1 U506 ( .A1(n470), .A2(n465), .ZN(n643) );
  AND2_X1 U507 ( .A1(n467), .A2(n466), .ZN(n465) );
  INV_X1 U508 ( .A(KEYINPUT19), .ZN(n525) );
  NOR2_X1 U509 ( .A1(n608), .A2(n381), .ZN(n527) );
  INV_X1 U510 ( .A(n658), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n483), .B(n482), .ZN(n748) );
  XNOR2_X1 U512 ( .A(n536), .B(n552), .ZN(n482) );
  XNOR2_X1 U513 ( .A(n769), .B(n448), .ZN(n483) );
  NOR2_X1 U514 ( .A1(n729), .A2(n486), .ZN(n730) );
  INV_X1 U515 ( .A(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U516 ( .A(n464), .B(KEYINPUT40), .ZN(n784) );
  INV_X1 U517 ( .A(n690), .ZN(n438) );
  XNOR2_X1 U518 ( .A(n516), .B(n515), .ZN(n514) );
  INV_X1 U519 ( .A(KEYINPUT36), .ZN(n515) );
  XNOR2_X1 U520 ( .A(KEYINPUT35), .B(KEYINPUT80), .ZN(n520) );
  INV_X1 U521 ( .A(n647), .ZN(n616) );
  INV_X1 U522 ( .A(KEYINPUT31), .ZN(n460) );
  INV_X1 U523 ( .A(n709), .ZN(n492) );
  NAND2_X1 U524 ( .A1(n623), .A2(n622), .ZN(n694) );
  NAND2_X1 U525 ( .A1(n531), .A2(n500), .ZN(n530) );
  NAND2_X1 U526 ( .A1(n504), .A2(n500), .ZN(n498) );
  XNOR2_X1 U527 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U528 ( .A(n497), .B(G116), .ZN(n496) );
  OR2_X1 U529 ( .A1(n477), .A2(n471), .ZN(n357) );
  NAND2_X1 U530 ( .A1(n519), .A2(n476), .ZN(n358) );
  AND2_X1 U531 ( .A1(n419), .A2(n418), .ZN(n359) );
  AND2_X1 U532 ( .A1(n511), .A2(n512), .ZN(n360) );
  XOR2_X1 U533 ( .A(n611), .B(KEYINPUT88), .Z(n657) );
  NOR2_X1 U534 ( .A1(n722), .A2(n486), .ZN(n361) );
  INV_X1 U535 ( .A(G472), .ZN(n519) );
  AND2_X1 U536 ( .A1(n527), .A2(n611), .ZN(n362) );
  XOR2_X1 U537 ( .A(KEYINPUT0), .B(KEYINPUT86), .Z(n363) );
  XOR2_X1 U538 ( .A(n613), .B(n612), .Z(n364) );
  XOR2_X1 U539 ( .A(n747), .B(KEYINPUT122), .Z(n365) );
  XNOR2_X1 U540 ( .A(n674), .B(KEYINPUT59), .ZN(n366) );
  XOR2_X1 U541 ( .A(n607), .B(KEYINPUT62), .Z(n367) );
  XOR2_X1 U542 ( .A(n676), .B(KEYINPUT60), .Z(n368) );
  NOR2_X1 U543 ( .A1(G952), .A2(n774), .ZN(n753) );
  INV_X1 U544 ( .A(n753), .ZN(n500) );
  INV_X1 U545 ( .A(n561), .ZN(n401) );
  XNOR2_X2 U546 ( .A(n369), .B(n496), .ZN(n561) );
  XNOR2_X2 U547 ( .A(n495), .B(n494), .ZN(n369) );
  XNOR2_X2 U548 ( .A(n761), .B(n374), .ZN(n373) );
  NAND2_X2 U549 ( .A1(n376), .A2(n375), .ZN(n761) );
  NAND2_X1 U550 ( .A1(n561), .A2(n489), .ZN(n375) );
  XNOR2_X2 U551 ( .A(n377), .B(n547), .ZN(n484) );
  NAND2_X1 U552 ( .A1(n378), .A2(n784), .ZN(n430) );
  XNOR2_X1 U553 ( .A(n378), .B(G137), .ZN(G39) );
  NAND2_X1 U554 ( .A1(n387), .A2(n638), .ZN(n386) );
  INV_X1 U555 ( .A(n397), .ZN(n389) );
  NAND2_X1 U556 ( .A1(n397), .A2(n396), .ZN(n395) );
  AND2_X1 U557 ( .A1(n783), .A2(KEYINPUT81), .ZN(n396) );
  INV_X1 U558 ( .A(n660), .ZN(n398) );
  XNOR2_X1 U559 ( .A(n424), .B(n423), .ZN(n399) );
  AND2_X1 U560 ( .A1(n435), .A2(n362), .ZN(n526) );
  INV_X1 U561 ( .A(n561), .ZN(n402) );
  INV_X1 U562 ( .A(n489), .ZN(n403) );
  XNOR2_X1 U563 ( .A(n581), .B(KEYINPUT16), .ZN(n489) );
  XNOR2_X1 U564 ( .A(n675), .B(n366), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n532), .B(n365), .ZN(n531) );
  NAND2_X1 U566 ( .A1(n635), .A2(n636), .ZN(n659) );
  INV_X1 U567 ( .A(n659), .ZN(n517) );
  INV_X1 U568 ( .A(n757), .ZN(n420) );
  NOR2_X1 U569 ( .A1(n716), .A2(n700), .ZN(n601) );
  AND2_X2 U570 ( .A1(n628), .A2(n610), .ZN(n446) );
  XNOR2_X2 U571 ( .A(n406), .B(n405), .ZN(n638) );
  NAND2_X1 U572 ( .A1(n757), .A2(n422), .ZN(n419) );
  XNOR2_X2 U573 ( .A(n442), .B(n458), .ZN(n757) );
  NAND2_X1 U574 ( .A1(n429), .A2(n426), .ZN(n437) );
  XNOR2_X1 U575 ( .A(n430), .B(n656), .ZN(n429) );
  XNOR2_X1 U576 ( .A(n411), .B(n505), .ZN(n410) );
  NAND2_X1 U577 ( .A1(n488), .A2(n687), .ZN(n427) );
  XNOR2_X1 U578 ( .A(n592), .B(n408), .ZN(n593) );
  INV_X2 U579 ( .A(n666), .ZN(n660) );
  XNOR2_X1 U580 ( .A(n409), .B(n459), .ZN(n445) );
  NAND2_X1 U581 ( .A1(n412), .A2(n410), .ZN(n409) );
  NAND2_X1 U582 ( .A1(n434), .A2(n677), .ZN(n411) );
  NAND2_X1 U583 ( .A1(n413), .A2(KEYINPUT44), .ZN(n412) );
  NAND2_X1 U584 ( .A1(n436), .A2(n447), .ZN(n413) );
  NAND2_X1 U585 ( .A1(n415), .A2(n359), .ZN(n432) );
  NAND2_X2 U586 ( .A1(n416), .A2(n415), .ZN(n424) );
  INV_X1 U587 ( .A(KEYINPUT2), .ZN(n422) );
  XNOR2_X2 U588 ( .A(n431), .B(n534), .ZN(n635) );
  NAND2_X1 U589 ( .A1(n432), .A2(n728), .ZN(n731) );
  NAND2_X1 U590 ( .A1(n433), .A2(n717), .ZN(n434) );
  XNOR2_X1 U591 ( .A(n621), .B(KEYINPUT96), .ZN(n433) );
  NOR2_X1 U592 ( .A1(n782), .A2(n400), .ZN(n436) );
  XNOR2_X2 U593 ( .A(n446), .B(n528), .ZN(n447) );
  NAND2_X1 U594 ( .A1(n440), .A2(n438), .ZN(n464) );
  AND2_X1 U595 ( .A1(n440), .A2(n439), .ZN(n669) );
  INV_X1 U596 ( .A(n668), .ZN(n439) );
  XNOR2_X1 U597 ( .A(n655), .B(n441), .ZN(n440) );
  INV_X1 U598 ( .A(KEYINPUT39), .ZN(n441) );
  NAND2_X1 U599 ( .A1(n445), .A2(n443), .ZN(n442) );
  NAND2_X1 U600 ( .A1(n444), .A2(n360), .ZN(n443) );
  INV_X1 U601 ( .A(n447), .ZN(n781) );
  XNOR2_X2 U602 ( .A(n510), .B(G146), .ZN(n485) );
  NAND2_X1 U603 ( .A1(n735), .A2(n670), .ZN(n562) );
  XNOR2_X2 U604 ( .A(n461), .B(n460), .ZN(n693) );
  NAND2_X1 U605 ( .A1(n602), .A2(n492), .ZN(n461) );
  NAND2_X1 U606 ( .A1(n607), .A2(G472), .ZN(n479) );
  OR2_X1 U607 ( .A1(n713), .A2(n472), .ZN(n466) );
  INV_X1 U608 ( .A(n471), .ZN(n468) );
  INV_X1 U609 ( .A(n475), .ZN(n469) );
  XNOR2_X2 U610 ( .A(n480), .B(n363), .ZN(n602) );
  NAND2_X1 U611 ( .A1(n639), .A2(n572), .ZN(n480) );
  XNOR2_X1 U612 ( .A(n481), .B(n525), .ZN(n639) );
  NOR2_X2 U613 ( .A1(n666), .A2(n565), .ZN(n481) );
  NAND2_X1 U614 ( .A1(n641), .A2(n642), .ZN(n488) );
  INV_X1 U615 ( .A(n651), .ZN(n490) );
  AND2_X1 U616 ( .A1(n602), .A2(n493), .ZN(n615) );
  AND2_X1 U617 ( .A1(n602), .A2(n637), .ZN(n619) );
  XNOR2_X2 U618 ( .A(G119), .B(KEYINPUT70), .ZN(n494) );
  XNOR2_X2 U619 ( .A(KEYINPUT3), .B(G113), .ZN(n495) );
  XNOR2_X1 U620 ( .A(n498), .B(n368), .ZN(G60) );
  AND2_X2 U621 ( .A1(n746), .A2(G210), .ZN(n737) );
  NAND2_X1 U622 ( .A1(n602), .A2(n601), .ZN(n503) );
  INV_X1 U623 ( .A(n499), .ZN(n506) );
  NAND2_X1 U624 ( .A1(n501), .A2(n500), .ZN(n499) );
  XNOR2_X1 U625 ( .A(n671), .B(n367), .ZN(n501) );
  XNOR2_X1 U626 ( .A(n615), .B(KEYINPUT34), .ZN(n522) );
  NAND2_X1 U627 ( .A1(n746), .A2(G472), .ZN(n671) );
  NAND2_X1 U628 ( .A1(n617), .A2(n658), .ZN(n614) );
  XNOR2_X1 U629 ( .A(n506), .B(n673), .ZN(G57) );
  NAND2_X1 U630 ( .A1(n522), .A2(n616), .ZN(n521) );
  INV_X1 U631 ( .A(n781), .ZN(n512) );
  NAND2_X1 U632 ( .A1(n514), .A2(n657), .ZN(n529) );
  NAND2_X1 U633 ( .A1(n662), .A2(n660), .ZN(n516) );
  XNOR2_X2 U634 ( .A(n638), .B(n523), .ZN(n611) );
  NOR2_X2 U635 ( .A1(n611), .A2(n698), .ZN(n617) );
  XNOR2_X2 U636 ( .A(n562), .B(n563), .ZN(n666) );
  INV_X1 U637 ( .A(n529), .ZN(n696) );
  XNOR2_X1 U638 ( .A(n530), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U639 ( .A1(n399), .A2(G478), .ZN(n532) );
  XOR2_X1 U640 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n535) );
  AND2_X1 U641 ( .A1(n589), .A2(G221), .ZN(n536) );
  XNOR2_X1 U642 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U643 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U644 ( .A(n543), .B(n401), .ZN(n548) );
  BUF_X1 U645 ( .A(n399), .Z(n749) );
  XNOR2_X1 U646 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U647 ( .A(n672), .B(KEYINPUT85), .ZN(n673) );
  XOR2_X1 U648 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n538) );
  NAND2_X1 U649 ( .A1(n573), .A2(G210), .ZN(n537) );
  XNOR2_X1 U650 ( .A(n538), .B(n537), .ZN(n542) );
  XNOR2_X1 U651 ( .A(G137), .B(KEYINPUT93), .ZN(n540) );
  NAND2_X1 U652 ( .A1(G101), .A2(n772), .ZN(n545) );
  XOR2_X1 U653 ( .A(G137), .B(G140), .Z(n603) );
  INV_X1 U654 ( .A(n603), .ZN(n549) );
  XNOR2_X1 U655 ( .A(n551), .B(n550), .ZN(n552) );
  NAND2_X1 U656 ( .A1(n774), .A2(G234), .ZN(n554) );
  XNOR2_X1 U657 ( .A(n554), .B(n553), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n670), .A2(G234), .ZN(n556) );
  XNOR2_X1 U659 ( .A(n556), .B(n555), .ZN(n599) );
  NAND2_X1 U660 ( .A1(G217), .A2(n599), .ZN(n557) );
  INV_X1 U661 ( .A(n635), .ZN(n608) );
  NAND2_X1 U662 ( .A1(n564), .A2(G210), .ZN(n563) );
  NAND2_X1 U663 ( .A1(G224), .A2(n774), .ZN(n558) );
  XNOR2_X1 U664 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U665 ( .A1(G214), .A2(n564), .ZN(n713) );
  INV_X1 U666 ( .A(n713), .ZN(n565) );
  XNOR2_X1 U667 ( .A(n567), .B(n566), .ZN(n569) );
  NAND2_X1 U668 ( .A1(G952), .A2(n569), .ZN(n726) );
  NOR2_X1 U669 ( .A1(G953), .A2(n726), .ZN(n568) );
  XNOR2_X1 U670 ( .A(KEYINPUT89), .B(n568), .ZN(n632) );
  NAND2_X1 U671 ( .A1(G902), .A2(n569), .ZN(n629) );
  INV_X1 U672 ( .A(n629), .ZN(n570) );
  NOR2_X1 U673 ( .A1(G898), .A2(n774), .ZN(n766) );
  NAND2_X1 U674 ( .A1(n570), .A2(n766), .ZN(n571) );
  NAND2_X1 U675 ( .A1(n632), .A2(n571), .ZN(n572) );
  XNOR2_X1 U676 ( .A(KEYINPUT13), .B(G475), .ZN(n588) );
  NAND2_X1 U677 ( .A1(G214), .A2(n573), .ZN(n574) );
  XNOR2_X1 U678 ( .A(n575), .B(n574), .ZN(n579) );
  XNOR2_X1 U679 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U680 ( .A(n579), .B(n578), .Z(n584) );
  INV_X1 U681 ( .A(n580), .ZN(n582) );
  XNOR2_X1 U682 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U683 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U684 ( .A(n585), .B(n586), .Z(n674) );
  NOR2_X1 U685 ( .A1(G902), .A2(n674), .ZN(n587) );
  XNOR2_X1 U686 ( .A(n588), .B(n587), .ZN(n625) );
  INV_X1 U687 ( .A(n625), .ZN(n623) );
  NAND2_X1 U688 ( .A1(n589), .A2(G217), .ZN(n597) );
  XNOR2_X1 U689 ( .A(n591), .B(n590), .ZN(n594) );
  XOR2_X1 U690 ( .A(n594), .B(n593), .Z(n596) );
  XNOR2_X1 U691 ( .A(G134), .B(KEYINPUT9), .ZN(n595) );
  NOR2_X1 U692 ( .A1(n747), .A2(G902), .ZN(n598) );
  XNOR2_X1 U693 ( .A(n598), .B(G478), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n623), .A2(n624), .ZN(n716) );
  NAND2_X1 U695 ( .A1(n599), .A2(G221), .ZN(n600) );
  XOR2_X1 U696 ( .A(KEYINPUT21), .B(n600), .Z(n633) );
  INV_X1 U697 ( .A(n633), .ZN(n700) );
  NAND2_X1 U698 ( .A1(G227), .A2(n774), .ZN(n604) );
  INV_X1 U699 ( .A(n611), .ZN(n626) );
  INV_X1 U700 ( .A(n704), .ZN(n637) );
  XNOR2_X1 U701 ( .A(KEYINPUT101), .B(n608), .ZN(n701) );
  NAND2_X1 U702 ( .A1(n657), .A2(n701), .ZN(n609) );
  XNOR2_X1 U703 ( .A(KEYINPUT103), .B(n609), .ZN(n610) );
  INV_X1 U704 ( .A(n618), .ZN(n698) );
  XOR2_X1 U705 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n613) );
  INV_X1 U706 ( .A(n624), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n625), .A2(n622), .ZN(n647) );
  NAND2_X1 U708 ( .A1(n381), .A2(n617), .ZN(n709) );
  NAND2_X1 U709 ( .A1(n638), .A2(n618), .ZN(n644) );
  INV_X1 U710 ( .A(n644), .ZN(n620) );
  NAND2_X1 U711 ( .A1(n620), .A2(n619), .ZN(n682) );
  NAND2_X1 U712 ( .A1(n693), .A2(n682), .ZN(n621) );
  XNOR2_X1 U713 ( .A(KEYINPUT100), .B(n694), .ZN(n668) );
  NAND2_X1 U714 ( .A1(n625), .A2(n624), .ZN(n690) );
  NAND2_X1 U715 ( .A1(n668), .A2(n690), .ZN(n717) );
  NOR2_X1 U716 ( .A1(n701), .A2(n626), .ZN(n627) );
  NAND2_X1 U717 ( .A1(n628), .A2(n627), .ZN(n677) );
  INV_X1 U718 ( .A(KEYINPUT47), .ZN(n640) );
  XNOR2_X1 U719 ( .A(n640), .B(n717), .ZN(n642) );
  NOR2_X1 U720 ( .A1(G900), .A2(n629), .ZN(n630) );
  NAND2_X1 U721 ( .A1(G953), .A2(n630), .ZN(n631) );
  NAND2_X1 U722 ( .A1(n632), .A2(n631), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n645), .A2(n633), .ZN(n634) );
  XNOR2_X1 U724 ( .A(KEYINPUT69), .B(n634), .ZN(n636) );
  NAND2_X1 U725 ( .A1(n651), .A2(n639), .ZN(n688) );
  NAND2_X1 U726 ( .A1(n640), .A2(n688), .ZN(n641) );
  NOR2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n654), .A2(n647), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n660), .A2(n648), .ZN(n687) );
  XNOR2_X1 U731 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n656) );
  XNOR2_X2 U732 ( .A(n660), .B(n649), .ZN(n714) );
  XNOR2_X1 U733 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n650) );
  INV_X1 U734 ( .A(n714), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n688), .A2(KEYINPUT47), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n664) );
  NAND2_X1 U737 ( .A1(n662), .A2(n611), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U739 ( .A1(n398), .A2(n665), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n669), .B(KEYINPUT111), .ZN(n785) );
  XNOR2_X1 U741 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n672) );
  NAND2_X1 U742 ( .A1(G475), .A2(n399), .ZN(n675) );
  INV_X1 U743 ( .A(KEYINPUT121), .ZN(n676) );
  XNOR2_X1 U744 ( .A(G101), .B(n677), .ZN(G3) );
  NOR2_X1 U745 ( .A1(n690), .A2(n682), .ZN(n679) );
  XNOR2_X1 U746 ( .A(G104), .B(KEYINPUT113), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(G6) );
  XOR2_X1 U748 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n681) );
  XNOR2_X1 U749 ( .A(G107), .B(KEYINPUT27), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n681), .B(n680), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n694), .A2(n682), .ZN(n683) );
  XOR2_X1 U752 ( .A(n684), .B(n683), .Z(G9) );
  NOR2_X1 U753 ( .A1(n694), .A2(n688), .ZN(n686) );
  XNOR2_X1 U754 ( .A(G128), .B(KEYINPUT29), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n686), .B(n685), .ZN(G30) );
  XNOR2_X1 U756 ( .A(G143), .B(n687), .ZN(G45) );
  NOR2_X1 U757 ( .A1(n690), .A2(n688), .ZN(n689) );
  XOR2_X1 U758 ( .A(G146), .B(n689), .Z(G48) );
  NOR2_X1 U759 ( .A1(n690), .A2(n693), .ZN(n692) );
  XNOR2_X1 U760 ( .A(G113), .B(KEYINPUT115), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n692), .B(n691), .ZN(G15) );
  NOR2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U763 ( .A(G116), .B(n695), .Z(G18) );
  XNOR2_X1 U764 ( .A(G125), .B(n696), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n697), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U766 ( .A1(n611), .A2(n698), .ZN(n699) );
  XNOR2_X1 U767 ( .A(KEYINPUT50), .B(n699), .ZN(n707) );
  XOR2_X1 U768 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n703) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n703), .B(n702), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U774 ( .A(n710), .B(KEYINPUT118), .ZN(n711) );
  XNOR2_X1 U775 ( .A(KEYINPUT51), .B(n711), .ZN(n712) );
  NOR2_X1 U776 ( .A1(n729), .A2(n712), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n721) );
  INV_X1 U779 ( .A(n717), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U781 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U782 ( .A1(n723), .A2(n361), .ZN(n724) );
  XNOR2_X1 U783 ( .A(n724), .B(KEYINPUT52), .ZN(n725) );
  NOR2_X1 U784 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U785 ( .A(n727), .B(KEYINPUT119), .ZN(n728) );
  NOR2_X1 U786 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U787 ( .A(KEYINPUT120), .B(n732), .Z(n733) );
  NOR2_X1 U788 ( .A1(G953), .A2(n733), .ZN(n734) );
  XNOR2_X1 U789 ( .A(KEYINPUT53), .B(n734), .ZN(G75) );
  XNOR2_X1 U790 ( .A(n356), .B(n535), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U792 ( .A1(n738), .A2(n753), .ZN(n740) );
  XNOR2_X1 U793 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n739) );
  XNOR2_X1 U794 ( .A(n740), .B(n739), .ZN(G51) );
  NAND2_X1 U795 ( .A1(G469), .A2(n749), .ZN(n744) );
  XOR2_X1 U796 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n741) );
  NOR2_X1 U797 ( .A1(n753), .A2(n745), .ZN(G54) );
  XNOR2_X1 U798 ( .A(n748), .B(KEYINPUT124), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n749), .A2(G217), .ZN(n750) );
  XNOR2_X1 U800 ( .A(n751), .B(n750), .ZN(n752) );
  NOR2_X1 U801 ( .A1(n753), .A2(n752), .ZN(G66) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n754) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n754), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n755), .A2(G898), .ZN(n756) );
  XNOR2_X1 U805 ( .A(n756), .B(KEYINPUT125), .ZN(n759) );
  NOR2_X1 U806 ( .A1(n757), .A2(G953), .ZN(n758) );
  NOR2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U808 ( .A(n760), .B(KEYINPUT127), .ZN(n768) );
  XNOR2_X1 U809 ( .A(n761), .B(n762), .ZN(n763) );
  XNOR2_X1 U810 ( .A(n763), .B(KEYINPUT126), .ZN(n764) );
  XNOR2_X1 U811 ( .A(n764), .B(G101), .ZN(n765) );
  NOR2_X1 U812 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U813 ( .A(n768), .B(n767), .ZN(G69) );
  XNOR2_X1 U814 ( .A(n769), .B(n770), .ZN(n771) );
  XNOR2_X1 U815 ( .A(n772), .B(n771), .ZN(n776) );
  XNOR2_X1 U816 ( .A(n776), .B(n773), .ZN(n775) );
  NAND2_X1 U817 ( .A1(n775), .A2(n774), .ZN(n780) );
  XNOR2_X1 U818 ( .A(G227), .B(n776), .ZN(n777) );
  NAND2_X1 U819 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U820 ( .A1(G953), .A2(n778), .ZN(n779) );
  NAND2_X1 U821 ( .A1(n780), .A2(n779), .ZN(G72) );
  XOR2_X1 U822 ( .A(n781), .B(G119), .Z(G21) );
  XOR2_X1 U823 ( .A(n400), .B(G110), .Z(G12) );
  XOR2_X1 U824 ( .A(n782), .B(G122), .Z(G24) );
  XNOR2_X1 U825 ( .A(G140), .B(n783), .ZN(G42) );
  XNOR2_X1 U826 ( .A(n784), .B(G131), .ZN(G33) );
  XNOR2_X1 U827 ( .A(G134), .B(KEYINPUT116), .ZN(n786) );
  XNOR2_X1 U828 ( .A(n786), .B(n785), .ZN(G36) );
endmodule

