

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754;

  NOR2_X1 U375 ( .A1(n626), .A2(n723), .ZN(n627) );
  NOR2_X1 U376 ( .A1(n633), .A2(n723), .ZN(n635) );
  NOR2_X1 U377 ( .A1(n641), .A2(n723), .ZN(n643) );
  AND2_X2 U378 ( .A1(n355), .A2(n354), .ZN(n644) );
  NOR2_X1 U379 ( .A1(n593), .A2(n592), .ZN(n596) );
  XNOR2_X1 U380 ( .A(n582), .B(n581), .ZN(n708) );
  XNOR2_X1 U381 ( .A(n493), .B(n353), .ZN(n512) );
  INV_X1 U382 ( .A(n492), .ZN(n353) );
  XNOR2_X1 U383 ( .A(n405), .B(KEYINPUT97), .ZN(n490) );
  NAND2_X1 U384 ( .A1(n521), .A2(n518), .ZN(n403) );
  OR2_X1 U385 ( .A1(n645), .A2(G902), .ZN(n396) );
  XNOR2_X1 U386 ( .A(n394), .B(KEYINPUT25), .ZN(n395) );
  XNOR2_X1 U387 ( .A(n732), .B(n412), .ZN(n454) );
  XNOR2_X1 U388 ( .A(G902), .B(KEYINPUT92), .ZN(n390) );
  XNOR2_X1 U389 ( .A(KEYINPUT93), .B(G104), .ZN(n367) );
  INV_X1 U390 ( .A(G953), .ZN(n748) );
  XNOR2_X1 U391 ( .A(n607), .B(KEYINPUT73), .ZN(n563) );
  NAND2_X1 U392 ( .A1(n562), .A2(n609), .ZN(n607) );
  INV_X1 U393 ( .A(n715), .ZN(n354) );
  NAND2_X1 U394 ( .A1(n606), .A2(n366), .ZN(n355) );
  NAND2_X1 U395 ( .A1(n638), .A2(n440), .ZN(n417) );
  XNOR2_X1 U396 ( .A(n415), .B(n416), .ZN(n638) );
  NOR2_X1 U397 ( .A1(G953), .A2(G237), .ZN(n428) );
  XNOR2_X1 U398 ( .A(n417), .B(G472), .ZN(n496) );
  XNOR2_X1 U399 ( .A(n367), .B(G110), .ZN(n461) );
  INV_X1 U400 ( .A(KEYINPUT22), .ZN(n356) );
  BUF_X1 U401 ( .A(n618), .Z(n724) );
  NOR2_X1 U402 ( .A1(n601), .A2(n618), .ZN(n603) );
  INV_X1 U403 ( .A(n564), .ZN(n583) );
  BUF_X2 U404 ( .A(n496), .Z(n685) );
  XNOR2_X1 U405 ( .A(n375), .B(G469), .ZN(n526) );
  OR2_X1 U406 ( .A1(n650), .A2(G902), .ZN(n375) );
  INV_X2 U407 ( .A(KEYINPUT3), .ZN(n411) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n495) );
  NOR2_X1 U409 ( .A1(n564), .A2(n483), .ZN(n357) );
  INV_X1 U410 ( .A(n583), .ZN(n358) );
  XNOR2_X1 U411 ( .A(G143), .B(G128), .ZN(n359) );
  XNOR2_X1 U412 ( .A(G143), .B(G128), .ZN(n452) );
  XNOR2_X1 U413 ( .A(G125), .B(G146), .ZN(n360) );
  XNOR2_X1 U414 ( .A(G125), .B(G146), .ZN(n453) );
  XNOR2_X2 U415 ( .A(KEYINPUT4), .B(G101), .ZN(n412) );
  XNOR2_X1 U416 ( .A(n600), .B(n599), .ZN(n618) );
  XNOR2_X1 U417 ( .A(n568), .B(n497), .ZN(n578) );
  INV_X1 U418 ( .A(n496), .ZN(n568) );
  XNOR2_X1 U419 ( .A(n401), .B(n400), .ZN(n518) );
  OR2_X1 U420 ( .A1(n399), .A2(n398), .ZN(n401) );
  XNOR2_X1 U421 ( .A(n554), .B(n553), .ZN(n609) );
  NOR2_X1 U422 ( .A1(n628), .A2(n604), .ZN(n468) );
  INV_X1 U423 ( .A(KEYINPUT19), .ZN(n475) );
  NAND2_X1 U424 ( .A1(n526), .A2(n404), .ZN(n405) );
  AND2_X1 U425 ( .A1(n397), .A2(G217), .ZN(n394) );
  NAND2_X1 U426 ( .A1(n498), .A2(n578), .ZN(n504) );
  AND2_X1 U427 ( .A1(n625), .A2(G953), .ZN(n723) );
  NOR2_X1 U428 ( .A1(n358), .A2(n569), .ZN(n361) );
  NOR2_X1 U429 ( .A1(n521), .A2(n520), .ZN(n362) );
  XOR2_X1 U430 ( .A(n453), .B(n452), .Z(n363) );
  OR2_X1 U431 ( .A1(n478), .A2(n477), .ZN(n364) );
  NAND2_X1 U432 ( .A1(n467), .A2(G210), .ZN(n365) );
  BUF_X1 U433 ( .A(n576), .Z(n508) );
  BUF_X1 U434 ( .A(n644), .Z(n719) );
  XNOR2_X1 U435 ( .A(n468), .B(n365), .ZN(n472) );
  NAND2_X1 U436 ( .A1(n605), .A2(KEYINPUT2), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n363), .B(n454), .ZN(n459) );
  BUF_X1 U438 ( .A(n454), .Z(n413) );
  INV_X1 U439 ( .A(KEYINPUT80), .ZN(n602) );
  XNOR2_X1 U440 ( .A(n413), .B(G146), .ZN(n414) );
  NAND2_X1 U441 ( .A1(n472), .A2(n692), .ZN(n474) );
  XNOR2_X1 U442 ( .A(n412), .B(n741), .ZN(n372) );
  BUF_X1 U443 ( .A(n577), .Z(n679) );
  XNOR2_X1 U444 ( .A(n360), .B(n376), .ZN(n742) );
  XNOR2_X1 U445 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U446 ( .A(n526), .B(n484), .ZN(n580) );
  XNOR2_X1 U447 ( .A(n480), .B(KEYINPUT0), .ZN(n564) );
  BUF_X1 U448 ( .A(n607), .Z(n747) );
  XNOR2_X1 U449 ( .A(n374), .B(n373), .ZN(n650) );
  BUF_X1 U450 ( .A(n636), .Z(n637) );
  XNOR2_X1 U451 ( .A(n359), .B(G134), .ZN(n448) );
  XOR2_X1 U452 ( .A(KEYINPUT69), .B(G131), .Z(n437) );
  XNOR2_X1 U453 ( .A(n448), .B(n437), .ZN(n739) );
  XNOR2_X1 U454 ( .A(n739), .B(G146), .ZN(n374) );
  XNOR2_X1 U455 ( .A(G140), .B(G137), .ZN(n382) );
  XNOR2_X1 U456 ( .A(n382), .B(KEYINPUT95), .ZN(n741) );
  INV_X1 U457 ( .A(n461), .ZN(n370) );
  NAND2_X1 U458 ( .A1(G227), .A2(n748), .ZN(n368) );
  XNOR2_X1 U459 ( .A(n368), .B(G107), .ZN(n369) );
  XNOR2_X1 U460 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U461 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n376) );
  INV_X1 U462 ( .A(n742), .ZN(n380) );
  NAND2_X1 U463 ( .A1(n748), .A2(G234), .ZN(n378) );
  XNOR2_X1 U464 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n377) );
  XNOR2_X1 U465 ( .A(n378), .B(n377), .ZN(n443) );
  NAND2_X1 U466 ( .A1(n443), .A2(G221), .ZN(n379) );
  XNOR2_X1 U467 ( .A(n380), .B(n379), .ZN(n388) );
  XNOR2_X1 U468 ( .A(KEYINPUT24), .B(KEYINPUT71), .ZN(n381) );
  XNOR2_X1 U469 ( .A(n382), .B(n381), .ZN(n386) );
  XNOR2_X1 U470 ( .A(G119), .B(G128), .ZN(n384) );
  XNOR2_X1 U471 ( .A(G110), .B(KEYINPUT23), .ZN(n383) );
  XNOR2_X1 U472 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U473 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U474 ( .A(n388), .B(n387), .ZN(n645) );
  INV_X1 U475 ( .A(KEYINPUT15), .ZN(n389) );
  XNOR2_X2 U476 ( .A(n390), .B(n389), .ZN(n604) );
  INV_X1 U477 ( .A(n604), .ZN(n391) );
  NAND2_X1 U478 ( .A1(n391), .A2(G234), .ZN(n393) );
  XNOR2_X1 U479 ( .A(KEYINPUT20), .B(KEYINPUT96), .ZN(n392) );
  XNOR2_X1 U480 ( .A(n393), .B(n392), .ZN(n397) );
  XNOR2_X2 U481 ( .A(n395), .B(n396), .ZN(n521) );
  INV_X1 U482 ( .A(n397), .ZN(n399) );
  INV_X1 U483 ( .A(G221), .ZN(n398) );
  INV_X1 U484 ( .A(KEYINPUT21), .ZN(n400) );
  INV_X1 U485 ( .A(KEYINPUT67), .ZN(n402) );
  XNOR2_X2 U486 ( .A(n403), .B(n402), .ZN(n577) );
  INV_X1 U487 ( .A(n577), .ZN(n404) );
  XOR2_X1 U488 ( .A(G137), .B(KEYINPUT98), .Z(n407) );
  NAND2_X1 U489 ( .A1(n428), .A2(G210), .ZN(n406) );
  XNOR2_X1 U490 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U491 ( .A(n408), .B(KEYINPUT5), .Z(n410) );
  XNOR2_X1 U492 ( .A(G116), .B(G113), .ZN(n409) );
  XNOR2_X1 U493 ( .A(n410), .B(n409), .ZN(n416) );
  XNOR2_X2 U494 ( .A(n411), .B(G119), .ZN(n732) );
  XNOR2_X1 U495 ( .A(n739), .B(n414), .ZN(n415) );
  INV_X1 U496 ( .A(G902), .ZN(n440) );
  INV_X1 U497 ( .A(G237), .ZN(n418) );
  NAND2_X1 U498 ( .A1(n440), .A2(n418), .ZN(n467) );
  NAND2_X1 U499 ( .A1(n467), .A2(G214), .ZN(n692) );
  AND2_X1 U500 ( .A1(n685), .A2(n692), .ZN(n420) );
  INV_X1 U501 ( .A(KEYINPUT30), .ZN(n419) );
  XNOR2_X1 U502 ( .A(n420), .B(n419), .ZN(n489) );
  NAND2_X1 U503 ( .A1(G234), .A2(G237), .ZN(n421) );
  XNOR2_X1 U504 ( .A(n421), .B(KEYINPUT14), .ZN(n424) );
  NAND2_X1 U505 ( .A1(G902), .A2(n424), .ZN(n422) );
  XOR2_X1 U506 ( .A(KEYINPUT94), .B(n422), .Z(n423) );
  NAND2_X1 U507 ( .A1(G953), .A2(n423), .ZN(n476) );
  NOR2_X1 U508 ( .A1(G900), .A2(n476), .ZN(n425) );
  NAND2_X1 U509 ( .A1(G952), .A2(n424), .ZN(n707) );
  NOR2_X1 U510 ( .A1(n707), .A2(G953), .ZN(n477) );
  OR2_X1 U511 ( .A1(n425), .A2(n477), .ZN(n426) );
  XNOR2_X1 U512 ( .A(n426), .B(KEYINPUT77), .ZN(n487) );
  NOR2_X1 U513 ( .A1(n489), .A2(n487), .ZN(n427) );
  AND2_X1 U514 ( .A1(n490), .A2(n427), .ZN(n470) );
  XOR2_X1 U515 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n430) );
  NAND2_X1 U516 ( .A1(G214), .A2(n428), .ZN(n429) );
  XNOR2_X1 U517 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U518 ( .A(KEYINPUT100), .B(G140), .Z(n432) );
  XNOR2_X1 U519 ( .A(G143), .B(G104), .ZN(n431) );
  XNOR2_X1 U520 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U521 ( .A(n434), .B(n433), .Z(n435) );
  XNOR2_X1 U522 ( .A(n435), .B(n742), .ZN(n439) );
  INV_X1 U523 ( .A(G122), .ZN(n436) );
  XNOR2_X1 U524 ( .A(n436), .B(G113), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n437), .B(n462), .ZN(n438) );
  XNOR2_X1 U526 ( .A(n439), .B(n438), .ZN(n622) );
  NAND2_X1 U527 ( .A1(n622), .A2(n440), .ZN(n442) );
  XOR2_X1 U528 ( .A(KEYINPUT13), .B(G475), .Z(n441) );
  XNOR2_X1 U529 ( .A(n442), .B(n441), .ZN(n511) );
  XOR2_X1 U530 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n445) );
  NAND2_X1 U531 ( .A1(G217), .A2(n443), .ZN(n444) );
  XNOR2_X1 U532 ( .A(n445), .B(n444), .ZN(n450) );
  XOR2_X1 U533 ( .A(KEYINPUT101), .B(G122), .Z(n446) );
  XNOR2_X1 U534 ( .A(G116), .B(G107), .ZN(n460) );
  XNOR2_X1 U535 ( .A(n446), .B(n460), .ZN(n447) );
  XOR2_X1 U536 ( .A(n448), .B(n447), .Z(n449) );
  XNOR2_X1 U537 ( .A(n450), .B(n449), .ZN(n720) );
  NOR2_X1 U538 ( .A1(G902), .A2(n720), .ZN(n451) );
  XNOR2_X1 U539 ( .A(G478), .B(n451), .ZN(n510) );
  INV_X1 U540 ( .A(n510), .ZN(n481) );
  NAND2_X1 U541 ( .A1(n511), .A2(n481), .ZN(n585) );
  XOR2_X1 U542 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n457) );
  NAND2_X1 U543 ( .A1(G224), .A2(n748), .ZN(n455) );
  XNOR2_X1 U544 ( .A(n455), .B(KEYINPUT74), .ZN(n456) );
  XNOR2_X1 U545 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U546 ( .A(n459), .B(n458), .ZN(n466) );
  XNOR2_X1 U547 ( .A(n461), .B(n460), .ZN(n465) );
  INV_X1 U548 ( .A(n462), .ZN(n463) );
  XNOR2_X1 U549 ( .A(n463), .B(KEYINPUT16), .ZN(n464) );
  XNOR2_X1 U550 ( .A(n465), .B(n464), .ZN(n734) );
  XNOR2_X1 U551 ( .A(n466), .B(n734), .ZN(n628) );
  INV_X1 U552 ( .A(n472), .ZN(n558) );
  NOR2_X1 U553 ( .A1(n585), .A2(n558), .ZN(n469) );
  NAND2_X1 U554 ( .A1(n470), .A2(n469), .ZN(n542) );
  XNOR2_X1 U555 ( .A(G143), .B(KEYINPUT116), .ZN(n471) );
  XNOR2_X1 U556 ( .A(n542), .B(n471), .ZN(G45) );
  INV_X1 U557 ( .A(KEYINPUT89), .ZN(n473) );
  XNOR2_X2 U558 ( .A(n474), .B(n473), .ZN(n535) );
  XNOR2_X1 U559 ( .A(n535), .B(n475), .ZN(n543) );
  INV_X1 U560 ( .A(n543), .ZN(n479) );
  NOR2_X1 U561 ( .A1(n476), .A2(G898), .ZN(n478) );
  NAND2_X1 U562 ( .A1(n479), .A2(n364), .ZN(n480) );
  OR2_X1 U563 ( .A1(n511), .A2(n481), .ZN(n696) );
  INV_X1 U564 ( .A(n518), .ZN(n674) );
  NOR2_X1 U565 ( .A1(n696), .A2(n674), .ZN(n482) );
  XNOR2_X1 U566 ( .A(n482), .B(KEYINPUT103), .ZN(n483) );
  XNOR2_X1 U567 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n484) );
  INV_X1 U568 ( .A(n580), .ZN(n678) );
  NOR2_X1 U569 ( .A1(n685), .A2(n521), .ZN(n485) );
  NAND2_X1 U570 ( .A1(n678), .A2(n485), .ZN(n486) );
  OR2_X1 U571 ( .A1(n495), .A2(n486), .ZN(n591) );
  XNOR2_X1 U572 ( .A(n591), .B(G110), .ZN(G12) );
  INV_X1 U573 ( .A(n487), .ZN(n519) );
  XNOR2_X1 U574 ( .A(n558), .B(KEYINPUT38), .ZN(n693) );
  NAND2_X1 U575 ( .A1(n519), .A2(n693), .ZN(n488) );
  NOR2_X1 U576 ( .A1(n489), .A2(n488), .ZN(n491) );
  NAND2_X1 U577 ( .A1(n491), .A2(n490), .ZN(n493) );
  XNOR2_X1 U578 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n492) );
  OR2_X1 U579 ( .A1(n511), .A2(n510), .ZN(n659) );
  XNOR2_X1 U580 ( .A(n659), .B(KEYINPUT102), .ZN(n546) );
  INV_X1 U581 ( .A(n546), .ZN(n494) );
  AND2_X1 U582 ( .A1(n512), .A2(n494), .ZN(n610) );
  XOR2_X1 U583 ( .A(G134), .B(n610), .Z(G36) );
  INV_X1 U584 ( .A(n495), .ZN(n498) );
  INV_X1 U585 ( .A(KEYINPUT6), .ZN(n497) );
  INV_X1 U586 ( .A(KEYINPUT91), .ZN(n499) );
  XNOR2_X1 U587 ( .A(n580), .B(n499), .ZN(n540) );
  INV_X1 U588 ( .A(n521), .ZN(n675) );
  NAND2_X1 U589 ( .A1(n540), .A2(n675), .ZN(n500) );
  NOR2_X1 U590 ( .A1(n504), .A2(n500), .ZN(n502) );
  XNOR2_X1 U591 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n501) );
  XNOR2_X1 U592 ( .A(n502), .B(n501), .ZN(n593) );
  XOR2_X1 U593 ( .A(n593), .B(G119), .Z(G21) );
  INV_X1 U594 ( .A(KEYINPUT86), .ZN(n503) );
  XNOR2_X1 U595 ( .A(n504), .B(n503), .ZN(n505) );
  NAND2_X1 U596 ( .A1(n505), .A2(n678), .ZN(n506) );
  XNOR2_X1 U597 ( .A(n506), .B(KEYINPUT87), .ZN(n507) );
  NAND2_X1 U598 ( .A1(n507), .A2(n521), .ZN(n576) );
  XNOR2_X1 U599 ( .A(n508), .B(G101), .ZN(G3) );
  AND2_X1 U600 ( .A1(n511), .A2(n510), .ZN(n666) );
  NAND2_X1 U601 ( .A1(n512), .A2(n666), .ZN(n515) );
  INV_X1 U602 ( .A(KEYINPUT109), .ZN(n513) );
  XNOR2_X1 U603 ( .A(n513), .B(KEYINPUT40), .ZN(n514) );
  XNOR2_X1 U604 ( .A(n515), .B(n514), .ZN(n636) );
  NAND2_X1 U605 ( .A1(n693), .A2(n692), .ZN(n699) );
  NOR2_X1 U606 ( .A1(n696), .A2(n699), .ZN(n517) );
  XNOR2_X1 U607 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U608 ( .A(n517), .B(n516), .ZN(n709) );
  NAND2_X1 U609 ( .A1(n519), .A2(n518), .ZN(n520) );
  AND2_X1 U610 ( .A1(n685), .A2(n362), .ZN(n524) );
  XOR2_X1 U611 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n522) );
  XNOR2_X1 U612 ( .A(KEYINPUT28), .B(n522), .ZN(n523) );
  XNOR2_X1 U613 ( .A(n524), .B(n523), .ZN(n525) );
  NAND2_X1 U614 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U615 ( .A(KEYINPUT108), .B(n527), .ZN(n544) );
  NOR2_X1 U616 ( .A1(n709), .A2(n544), .ZN(n529) );
  INV_X1 U617 ( .A(KEYINPUT42), .ZN(n528) );
  XNOR2_X1 U618 ( .A(n529), .B(n528), .ZN(n753) );
  NAND2_X1 U619 ( .A1(n636), .A2(n753), .ZN(n532) );
  XNOR2_X1 U620 ( .A(KEYINPUT84), .B(KEYINPUT46), .ZN(n530) );
  XOR2_X1 U621 ( .A(n530), .B(KEYINPUT64), .Z(n531) );
  XNOR2_X1 U622 ( .A(n532), .B(n531), .ZN(n551) );
  INV_X1 U623 ( .A(n666), .ZN(n545) );
  NOR2_X1 U624 ( .A1(n578), .A2(n545), .ZN(n533) );
  NAND2_X1 U625 ( .A1(n362), .A2(n533), .ZN(n534) );
  XNOR2_X1 U626 ( .A(KEYINPUT104), .B(n534), .ZN(n555) );
  BUF_X1 U627 ( .A(n535), .Z(n536) );
  NOR2_X1 U628 ( .A1(n555), .A2(n536), .ZN(n539) );
  XOR2_X1 U629 ( .A(KEYINPUT88), .B(KEYINPUT111), .Z(n537) );
  XNOR2_X1 U630 ( .A(KEYINPUT36), .B(n537), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n539), .B(n538), .ZN(n541) );
  NAND2_X1 U632 ( .A1(n541), .A2(n540), .ZN(n672) );
  NAND2_X1 U633 ( .A1(n672), .A2(n542), .ZN(n549) );
  NOR2_X1 U634 ( .A1(n544), .A2(n543), .ZN(n664) );
  AND2_X1 U635 ( .A1(n546), .A2(n545), .ZN(n698) );
  INV_X1 U636 ( .A(n698), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n664), .A2(n570), .ZN(n547) );
  XNOR2_X1 U638 ( .A(n547), .B(KEYINPUT47), .ZN(n548) );
  NOR2_X1 U639 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U640 ( .A1(n551), .A2(n550), .ZN(n554) );
  INV_X1 U641 ( .A(KEYINPUT70), .ZN(n552) );
  XNOR2_X1 U642 ( .A(n552), .B(KEYINPUT48), .ZN(n553) );
  NOR2_X1 U643 ( .A1(n580), .A2(n555), .ZN(n556) );
  NAND2_X1 U644 ( .A1(n556), .A2(n692), .ZN(n557) );
  XNOR2_X1 U645 ( .A(n557), .B(KEYINPUT43), .ZN(n559) );
  AND2_X1 U646 ( .A1(n559), .A2(n558), .ZN(n561) );
  INV_X1 U647 ( .A(KEYINPUT105), .ZN(n560) );
  XNOR2_X1 U648 ( .A(n561), .B(n560), .ZN(n752) );
  NOR2_X1 U649 ( .A1(n752), .A2(n610), .ZN(n562) );
  NAND2_X1 U650 ( .A1(n563), .A2(n604), .ZN(n601) );
  NAND2_X1 U651 ( .A1(n580), .A2(n685), .ZN(n565) );
  OR2_X1 U652 ( .A1(n679), .A2(n565), .ZN(n673) );
  OR2_X1 U653 ( .A1(n358), .A2(n673), .ZN(n567) );
  XOR2_X1 U654 ( .A(KEYINPUT31), .B(KEYINPUT99), .Z(n566) );
  XNOR2_X1 U655 ( .A(n567), .B(n566), .ZN(n669) );
  NAND2_X1 U656 ( .A1(n490), .A2(n568), .ZN(n569) );
  OR2_X1 U657 ( .A1(n669), .A2(n361), .ZN(n571) );
  NAND2_X1 U658 ( .A1(n571), .A2(n570), .ZN(n574) );
  INV_X1 U659 ( .A(KEYINPUT72), .ZN(n572) );
  NAND2_X1 U660 ( .A1(n572), .A2(KEYINPUT44), .ZN(n573) );
  AND2_X1 U661 ( .A1(n574), .A2(n573), .ZN(n575) );
  AND2_X1 U662 ( .A1(n576), .A2(n575), .ZN(n598) );
  NOR2_X1 U663 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U664 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U665 ( .A(KEYINPUT33), .ZN(n581) );
  NOR2_X1 U666 ( .A1(n564), .A2(n708), .ZN(n584) );
  XNOR2_X1 U667 ( .A(n584), .B(KEYINPUT34), .ZN(n587) );
  XNOR2_X1 U668 ( .A(KEYINPUT75), .B(n585), .ZN(n586) );
  NAND2_X1 U669 ( .A1(n587), .A2(n586), .ZN(n590) );
  INV_X1 U670 ( .A(KEYINPUT82), .ZN(n588) );
  XNOR2_X1 U671 ( .A(n588), .B(KEYINPUT35), .ZN(n589) );
  XNOR2_X2 U672 ( .A(n590), .B(n589), .ZN(n754) );
  NAND2_X1 U673 ( .A1(n754), .A2(n591), .ZN(n592) );
  INV_X1 U674 ( .A(KEYINPUT44), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n594), .A2(KEYINPUT72), .ZN(n595) );
  XNOR2_X1 U676 ( .A(n596), .B(n595), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X1 U678 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n603), .B(n602), .ZN(n606) );
  XOR2_X1 U680 ( .A(KEYINPUT81), .B(n604), .Z(n605) );
  NAND2_X1 U681 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n747), .A2(n608), .ZN(n617) );
  INV_X1 U683 ( .A(n609), .ZN(n615) );
  NOR2_X1 U684 ( .A1(n752), .A2(KEYINPUT78), .ZN(n613) );
  INV_X1 U685 ( .A(n610), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n611), .A2(KEYINPUT2), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n619) );
  NOR2_X1 U690 ( .A1(n619), .A2(n724), .ZN(n715) );
  NAND2_X1 U691 ( .A1(n644), .A2(G475), .ZN(n624) );
  XOR2_X1 U692 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n624), .B(n623), .ZN(n626) );
  INV_X1 U695 ( .A(G952), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n627), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U697 ( .A1(n644), .A2(G210), .ZN(n632) );
  XOR2_X1 U698 ( .A(KEYINPUT90), .B(KEYINPUT54), .Z(n629) );
  XNOR2_X1 U699 ( .A(n629), .B(KEYINPUT55), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n628), .B(n630), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n633) );
  XOR2_X1 U702 ( .A(KEYINPUT83), .B(KEYINPUT56), .Z(n634) );
  XNOR2_X1 U703 ( .A(n635), .B(n634), .ZN(G51) );
  XNOR2_X1 U704 ( .A(n637), .B(G131), .ZN(G33) );
  NAND2_X1 U705 ( .A1(n644), .A2(G472), .ZN(n640) );
  XOR2_X1 U706 ( .A(KEYINPUT62), .B(n638), .Z(n639) );
  XNOR2_X1 U707 ( .A(n640), .B(n639), .ZN(n641) );
  XOR2_X1 U708 ( .A(KEYINPUT112), .B(KEYINPUT63), .Z(n642) );
  XNOR2_X1 U709 ( .A(n643), .B(n642), .ZN(G57) );
  NAND2_X1 U710 ( .A1(n719), .A2(G217), .ZN(n647) );
  XNOR2_X1 U711 ( .A(n645), .B(KEYINPUT124), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U713 ( .A1(n648), .A2(n723), .ZN(G66) );
  NAND2_X1 U714 ( .A1(n719), .A2(G469), .ZN(n652) );
  XOR2_X1 U715 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n649) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U718 ( .A1(n653), .A2(n723), .ZN(G54) );
  XOR2_X1 U719 ( .A(G104), .B(KEYINPUT113), .Z(n655) );
  NAND2_X1 U720 ( .A1(n361), .A2(n666), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(G6) );
  XOR2_X1 U722 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n657) );
  XNOR2_X1 U723 ( .A(G107), .B(KEYINPUT114), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U725 ( .A(KEYINPUT26), .B(n658), .Z(n661) );
  INV_X1 U726 ( .A(n659), .ZN(n668) );
  NAND2_X1 U727 ( .A1(n361), .A2(n668), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n661), .B(n660), .ZN(G9) );
  XOR2_X1 U729 ( .A(G128), .B(KEYINPUT29), .Z(n663) );
  NAND2_X1 U730 ( .A1(n664), .A2(n668), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(G30) );
  NAND2_X1 U732 ( .A1(n664), .A2(n666), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(G146), .ZN(G48) );
  NAND2_X1 U734 ( .A1(n669), .A2(n666), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(G113), .ZN(G15) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(G116), .ZN(G18) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(G27) );
  INV_X1 U740 ( .A(n673), .ZN(n688) );
  NAND2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U742 ( .A(n676), .B(KEYINPUT49), .ZN(n677) );
  XNOR2_X1 U743 ( .A(KEYINPUT117), .B(n677), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n680), .B(KEYINPUT118), .ZN(n681) );
  XNOR2_X1 U746 ( .A(KEYINPUT50), .B(n681), .ZN(n682) );
  NAND2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U749 ( .A(KEYINPUT119), .B(n686), .Z(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U751 ( .A(KEYINPUT120), .B(n689), .Z(n690) );
  XNOR2_X1 U752 ( .A(n690), .B(KEYINPUT51), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n709), .A2(n691), .ZN(n704) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U755 ( .A(KEYINPUT121), .B(n694), .Z(n695) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U757 ( .A(n697), .B(KEYINPUT122), .ZN(n701) );
  NOR2_X1 U758 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U759 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n702), .A2(n708), .ZN(n703) );
  NOR2_X1 U761 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U762 ( .A(n705), .B(KEYINPUT52), .ZN(n706) );
  NOR2_X1 U763 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U766 ( .A1(n712), .A2(n748), .ZN(n717) );
  NOR2_X1 U767 ( .A1(n724), .A2(n747), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n713), .A2(KEYINPUT2), .ZN(n714) );
  NOR2_X1 U769 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U770 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n718), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U772 ( .A1(n719), .A2(G478), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U774 ( .A1(n723), .A2(n722), .ZN(G63) );
  NOR2_X1 U775 ( .A1(n724), .A2(G953), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n725), .B(KEYINPUT127), .ZN(n731) );
  XOR2_X1 U777 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n727) );
  NAND2_X1 U778 ( .A1(G224), .A2(G953), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U780 ( .A(KEYINPUT125), .B(n728), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n738) );
  XNOR2_X1 U783 ( .A(n732), .B(G101), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(n733), .ZN(n736) );
  NOR2_X1 U785 ( .A1(G898), .A2(n748), .ZN(n735) );
  NOR2_X1 U786 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n738), .B(n737), .ZN(G69) );
  XNOR2_X1 U788 ( .A(KEYINPUT4), .B(n739), .ZN(n740) );
  XNOR2_X1 U789 ( .A(n741), .B(n740), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n743), .B(n742), .ZN(n746) );
  XNOR2_X1 U791 ( .A(G227), .B(n746), .ZN(n744) );
  NAND2_X1 U792 ( .A1(G900), .A2(n744), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G953), .ZN(n751) );
  XNOR2_X1 U794 ( .A(n747), .B(n746), .ZN(n749) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U796 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U797 ( .A(G140), .B(n752), .Z(G42) );
  XNOR2_X1 U798 ( .A(G137), .B(n753), .ZN(G39) );
  XNOR2_X1 U799 ( .A(n754), .B(G122), .ZN(G24) );
endmodule

