

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762;

  AND2_X1 U377 ( .A1(n679), .A2(KEYINPUT2), .ZN(n642) );
  AND2_X1 U378 ( .A1(n570), .A2(n534), .ZN(n544) );
  BUF_X1 U379 ( .A(n539), .Z(n558) );
  NAND2_X1 U380 ( .A1(n408), .A2(n363), .ZN(n411) );
  INV_X2 U381 ( .A(G953), .ZN(n459) );
  OR2_X2 U382 ( .A1(n649), .A2(n580), .ZN(n437) );
  XNOR2_X2 U383 ( .A(n411), .B(n410), .ZN(n643) );
  AND2_X1 U384 ( .A1(n528), .A2(n689), .ZN(n549) );
  XNOR2_X2 U385 ( .A(n592), .B(KEYINPUT1), .ZN(n689) );
  XNOR2_X1 U386 ( .A(n527), .B(KEYINPUT32), .ZN(n531) );
  AND2_X1 U387 ( .A1(n567), .A2(n566), .ZN(n577) );
  AND2_X1 U388 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U389 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U390 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U391 ( .A(n465), .B(n464), .ZN(n552) );
  OR2_X1 U392 ( .A1(n732), .A2(G902), .ZN(n465) );
  XNOR2_X1 U393 ( .A(n726), .B(n725), .ZN(n727) );
  INV_X1 U394 ( .A(G143), .ZN(n663) );
  XNOR2_X1 U395 ( .A(G146), .B(G125), .ZN(n468) );
  XOR2_X1 U396 ( .A(KEYINPUT99), .B(KEYINPUT97), .Z(n454) );
  XNOR2_X1 U397 ( .A(G137), .B(G140), .ZN(n516) );
  NAND2_X1 U398 ( .A1(n409), .A2(n382), .ZN(n408) );
  XNOR2_X1 U399 ( .A(n417), .B(G107), .ZN(n452) );
  INV_X1 U400 ( .A(G122), .ZN(n417) );
  XNOR2_X1 U401 ( .A(n468), .B(KEYINPUT10), .ZN(n748) );
  NOR2_X1 U402 ( .A1(n612), .A2(n664), .ZN(n613) );
  XNOR2_X1 U403 ( .A(n369), .B(KEYINPUT46), .ZN(n368) );
  NOR2_X1 U404 ( .A1(n760), .A2(n762), .ZN(n369) );
  XNOR2_X1 U405 ( .A(n663), .B(G128), .ZN(n451) );
  NAND2_X1 U406 ( .A1(G234), .A2(G237), .ZN(n440) );
  XNOR2_X1 U407 ( .A(n393), .B(n392), .ZN(n598) );
  INV_X1 U408 ( .A(KEYINPUT19), .ZN(n392) );
  XNOR2_X1 U409 ( .A(G116), .B(G101), .ZN(n420) );
  INV_X1 U410 ( .A(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U411 ( .A(n451), .B(n450), .ZN(n488) );
  INV_X1 U412 ( .A(G134), .ZN(n450) );
  XNOR2_X1 U413 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U414 ( .A(KEYINPUT7), .B(n452), .Z(n456) );
  XNOR2_X1 U415 ( .A(KEYINPUT9), .B(KEYINPUT98), .ZN(n453) );
  XNOR2_X1 U416 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n460) );
  XNOR2_X1 U417 ( .A(G143), .B(G122), .ZN(n466) );
  XOR2_X1 U418 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n471) );
  XNOR2_X1 U419 ( .A(n469), .B(G140), .ZN(n396) );
  INV_X1 U420 ( .A(KEYINPUT64), .ZN(n410) );
  AND2_X1 U421 ( .A1(n594), .A2(n593), .ZN(n629) );
  NOR2_X1 U422 ( .A1(n688), .A2(n615), .ZN(n591) );
  XNOR2_X1 U423 ( .A(n376), .B(n374), .ZN(n698) );
  XNOR2_X1 U424 ( .A(n628), .B(n375), .ZN(n374) );
  NAND2_X1 U425 ( .A1(n377), .A2(n483), .ZN(n376) );
  INV_X1 U426 ( .A(KEYINPUT107), .ZN(n375) );
  NAND2_X1 U427 ( .A1(n358), .A2(n668), .ZN(n633) );
  NAND2_X1 U428 ( .A1(n398), .A2(n701), .ZN(n397) );
  INV_X1 U429 ( .A(n615), .ZN(n398) );
  BUF_X1 U430 ( .A(n610), .Z(n373) );
  NAND2_X1 U431 ( .A1(n383), .A2(n387), .ZN(n372) );
  NOR2_X1 U432 ( .A1(n642), .A2(n384), .ZN(n383) );
  INV_X1 U433 ( .A(G472), .ZN(n384) );
  XNOR2_X1 U434 ( .A(n406), .B(n405), .ZN(n736) );
  XNOR2_X1 U435 ( .A(n518), .B(n356), .ZN(n405) );
  XNOR2_X1 U436 ( .A(n519), .B(n407), .ZN(n406) );
  NAND2_X1 U437 ( .A1(n385), .A2(n387), .ZN(n381) );
  NOR2_X1 U438 ( .A1(n642), .A2(n386), .ZN(n385) );
  INV_X1 U439 ( .A(G210), .ZN(n386) );
  INV_X1 U440 ( .A(G237), .ZN(n433) );
  XNOR2_X1 U441 ( .A(n367), .B(n364), .ZN(n400) );
  XOR2_X1 U442 ( .A(n489), .B(n488), .Z(n750) );
  INV_X1 U443 ( .A(G101), .ZN(n501) );
  XNOR2_X1 U444 ( .A(G107), .B(G104), .ZN(n502) );
  INV_X1 U445 ( .A(KEYINPUT70), .ZN(n423) );
  XNOR2_X1 U446 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n426) );
  INV_X1 U447 ( .A(n707), .ZN(n377) );
  XNOR2_X1 U448 ( .A(n610), .B(KEYINPUT38), .ZN(n702) );
  NOR2_X1 U449 ( .A1(n689), .A2(n690), .ZN(n553) );
  XNOR2_X1 U450 ( .A(n391), .B(KEYINPUT0), .ZN(n539) );
  XNOR2_X1 U451 ( .A(G137), .B(G113), .ZN(n493) );
  AND2_X1 U452 ( .A1(n400), .A2(n637), .ZN(n752) );
  XOR2_X1 U453 ( .A(KEYINPUT88), .B(G110), .Z(n512) );
  XNOR2_X1 U454 ( .A(G119), .B(G128), .ZN(n511) );
  XNOR2_X1 U455 ( .A(n515), .B(n514), .ZN(n407) );
  XNOR2_X1 U456 ( .A(n422), .B(n492), .ZN(n738) );
  XNOR2_X1 U457 ( .A(n488), .B(G116), .ZN(n458) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n726) );
  XNOR2_X1 U459 ( .A(n475), .B(n748), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n474), .B(n396), .ZN(n395) );
  NAND2_X1 U461 ( .A1(n390), .A2(n388), .ZN(n728) );
  NOR2_X1 U462 ( .A1(n642), .A2(n389), .ZN(n388) );
  INV_X1 U463 ( .A(G475), .ZN(n389) );
  NAND2_X1 U464 ( .A1(n718), .A2(n359), .ZN(n404) );
  NAND2_X1 U465 ( .A1(n355), .A2(n373), .ZN(n677) );
  NAND2_X1 U466 ( .A1(n629), .A2(n698), .ZN(n630) );
  NOR2_X1 U467 ( .A1(n633), .A2(n373), .ZN(n616) );
  NOR2_X1 U468 ( .A1(n611), .A2(n373), .ZN(n664) );
  XNOR2_X1 U469 ( .A(n372), .B(n360), .ZN(n371) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n381), .B(n361), .ZN(n380) );
  XNOR2_X1 U472 ( .A(n403), .B(n401), .ZN(G75) );
  XNOR2_X1 U473 ( .A(n402), .B(KEYINPUT53), .ZN(n401) );
  OR2_X1 U474 ( .A1(n682), .A2(n404), .ZN(n403) );
  INV_X1 U475 ( .A(KEYINPUT120), .ZN(n402) );
  XNOR2_X1 U476 ( .A(n531), .B(n365), .ZN(G21) );
  AND2_X1 U477 ( .A1(n550), .A2(n399), .ZN(n668) );
  AND2_X1 U478 ( .A1(n637), .A2(n362), .ZN(n354) );
  XOR2_X1 U479 ( .A(n636), .B(KEYINPUT43), .Z(n355) );
  XOR2_X1 U480 ( .A(n512), .B(n511), .Z(n356) );
  AND2_X1 U481 ( .A1(n619), .A2(n618), .ZN(n357) );
  NOR2_X1 U482 ( .A1(n614), .A2(n397), .ZN(n358) );
  OR2_X1 U483 ( .A1(n681), .A2(n680), .ZN(n359) );
  XOR2_X1 U484 ( .A(n644), .B(KEYINPUT62), .Z(n360) );
  XOR2_X1 U485 ( .A(n649), .B(n648), .Z(n361) );
  NAND2_X1 U486 ( .A1(n582), .A2(n581), .ZN(n362) );
  NAND2_X1 U487 ( .A1(n362), .A2(n640), .ZN(n363) );
  XOR2_X1 U488 ( .A(KEYINPUT78), .B(KEYINPUT48), .Z(n364) );
  INV_X1 U489 ( .A(n737), .ZN(n379) );
  XOR2_X1 U490 ( .A(G119), .B(KEYINPUT127), .Z(n365) );
  XOR2_X1 U491 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n366) );
  NAND2_X1 U492 ( .A1(n357), .A2(n368), .ZN(n367) );
  XNOR2_X1 U493 ( .A(n370), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U494 ( .A1(n371), .A2(n379), .ZN(n370) );
  XNOR2_X1 U495 ( .A(n378), .B(n366), .ZN(G51) );
  NAND2_X1 U496 ( .A1(n380), .A2(n379), .ZN(n378) );
  AND2_X1 U497 ( .A1(n752), .A2(n382), .ZN(n679) );
  NAND2_X1 U498 ( .A1(n382), .A2(n459), .ZN(n741) );
  XNOR2_X2 U499 ( .A(n578), .B(KEYINPUT45), .ZN(n382) );
  NOR2_X1 U500 ( .A1(n643), .A2(n642), .ZN(n731) );
  INV_X1 U501 ( .A(n643), .ZN(n387) );
  INV_X1 U502 ( .A(n643), .ZN(n390) );
  NAND2_X1 U503 ( .A1(n731), .A2(G217), .ZN(n414) );
  NAND2_X1 U504 ( .A1(n598), .A2(n449), .ZN(n391) );
  NOR2_X2 U505 ( .A1(n610), .A2(n439), .ZN(n393) );
  XNOR2_X2 U506 ( .A(n437), .B(n436), .ZN(n610) );
  NOR2_X1 U507 ( .A1(n729), .A2(n737), .ZN(n730) );
  XNOR2_X1 U508 ( .A(n508), .B(n496), .ZN(n644) );
  NOR2_X1 U509 ( .A1(n550), .A2(n399), .ZN(n551) );
  INV_X1 U510 ( .A(n552), .ZN(n399) );
  AND2_X1 U511 ( .A1(n400), .A2(n354), .ZN(n409) );
  NOR2_X1 U512 ( .A1(n412), .A2(n737), .ZN(G66) );
  XNOR2_X1 U513 ( .A(n736), .B(n735), .ZN(n413) );
  XOR2_X1 U514 ( .A(n494), .B(n493), .Z(n415) );
  XNOR2_X1 U515 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U516 ( .A(KEYINPUT24), .ZN(n514) );
  XNOR2_X1 U517 ( .A(n504), .B(n503), .ZN(n506) );
  INV_X1 U518 ( .A(KEYINPUT90), .ZN(n556) );
  XNOR2_X1 U519 ( .A(n495), .B(n415), .ZN(n496) );
  XNOR2_X2 U520 ( .A(G113), .B(G104), .ZN(n473) );
  XNOR2_X1 U521 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n416) );
  XNOR2_X1 U522 ( .A(n473), .B(n416), .ZN(n418) );
  XNOR2_X1 U523 ( .A(n418), .B(n452), .ZN(n422) );
  XNOR2_X1 U524 ( .A(n419), .B(G119), .ZN(n421) );
  XNOR2_X1 U525 ( .A(n421), .B(n420), .ZN(n492) );
  XNOR2_X1 U526 ( .A(n423), .B(G110), .ZN(n500) );
  NAND2_X1 U527 ( .A1(n459), .A2(G224), .ZN(n424) );
  XNOR2_X1 U528 ( .A(n424), .B(KEYINPUT4), .ZN(n425) );
  XNOR2_X1 U529 ( .A(n500), .B(n425), .ZN(n429) );
  XNOR2_X1 U530 ( .A(n468), .B(n426), .ZN(n427) );
  XNOR2_X1 U531 ( .A(n427), .B(n451), .ZN(n428) );
  XNOR2_X1 U532 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U533 ( .A(n738), .B(n430), .ZN(n649) );
  XNOR2_X1 U534 ( .A(G902), .B(KEYINPUT83), .ZN(n432) );
  INV_X1 U535 ( .A(KEYINPUT15), .ZN(n431) );
  XNOR2_X1 U536 ( .A(n432), .B(n431), .ZN(n581) );
  INV_X1 U537 ( .A(n581), .ZN(n580) );
  INV_X1 U538 ( .A(G902), .ZN(n434) );
  NAND2_X1 U539 ( .A1(n434), .A2(n433), .ZN(n438) );
  NAND2_X1 U540 ( .A1(n438), .A2(G210), .ZN(n435) );
  XNOR2_X1 U541 ( .A(n435), .B(KEYINPUT84), .ZN(n436) );
  NAND2_X1 U542 ( .A1(n438), .A2(G214), .ZN(n701) );
  INV_X1 U543 ( .A(n701), .ZN(n439) );
  XNOR2_X1 U544 ( .A(n440), .B(KEYINPUT14), .ZN(n683) );
  INV_X1 U545 ( .A(n683), .ZN(n443) );
  NOR2_X1 U546 ( .A1(G898), .A2(n459), .ZN(n441) );
  XOR2_X1 U547 ( .A(KEYINPUT85), .B(n441), .Z(n739) );
  NAND2_X1 U548 ( .A1(G902), .A2(n739), .ZN(n442) );
  NOR2_X1 U549 ( .A1(n443), .A2(n442), .ZN(n445) );
  INV_X1 U550 ( .A(KEYINPUT86), .ZN(n444) );
  XNOR2_X1 U551 ( .A(n445), .B(n444), .ZN(n448) );
  NAND2_X1 U552 ( .A1(G952), .A2(n459), .ZN(n585) );
  INV_X1 U553 ( .A(n585), .ZN(n446) );
  NAND2_X1 U554 ( .A1(n683), .A2(n446), .ZN(n447) );
  NAND2_X1 U555 ( .A1(n448), .A2(n447), .ZN(n449) );
  XOR2_X1 U556 ( .A(n454), .B(n453), .Z(n455) );
  XNOR2_X1 U557 ( .A(n458), .B(n457), .ZN(n463) );
  NAND2_X1 U558 ( .A1(n459), .A2(G234), .ZN(n461) );
  XNOR2_X1 U559 ( .A(n461), .B(n460), .ZN(n513) );
  NAND2_X1 U560 ( .A1(G217), .A2(n513), .ZN(n462) );
  XNOR2_X1 U561 ( .A(n463), .B(n462), .ZN(n732) );
  XNOR2_X1 U562 ( .A(KEYINPUT100), .B(G478), .ZN(n464) );
  XOR2_X1 U563 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n467) );
  XNOR2_X1 U564 ( .A(n467), .B(n466), .ZN(n475) );
  NOR2_X1 U565 ( .A1(G953), .A2(G237), .ZN(n490) );
  NAND2_X1 U566 ( .A1(G214), .A2(n490), .ZN(n469) );
  XNOR2_X1 U567 ( .A(G131), .B(KEYINPUT11), .ZN(n470) );
  XNOR2_X1 U568 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U569 ( .A(n473), .B(n472), .ZN(n474) );
  NOR2_X1 U570 ( .A1(G902), .A2(n726), .ZN(n477) );
  XNOR2_X1 U571 ( .A(KEYINPUT13), .B(G475), .ZN(n476) );
  XNOR2_X1 U572 ( .A(n477), .B(n476), .ZN(n550) );
  NOR2_X1 U573 ( .A1(n552), .A2(n550), .ZN(n478) );
  XNOR2_X1 U574 ( .A(n478), .B(KEYINPUT103), .ZN(n704) );
  INV_X1 U575 ( .A(n704), .ZN(n483) );
  XOR2_X1 U576 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n480) );
  NAND2_X1 U577 ( .A1(G234), .A2(n581), .ZN(n479) );
  XNOR2_X1 U578 ( .A(n480), .B(n479), .ZN(n520) );
  AND2_X1 U579 ( .A1(n520), .A2(G221), .ZN(n482) );
  INV_X1 U580 ( .A(KEYINPUT21), .ZN(n481) );
  XNOR2_X1 U581 ( .A(n482), .B(n481), .ZN(n588) );
  NAND2_X1 U582 ( .A1(n483), .A2(n684), .ZN(n484) );
  NOR2_X2 U583 ( .A1(n539), .A2(n484), .ZN(n487) );
  INV_X1 U584 ( .A(KEYINPUT65), .ZN(n485) );
  XNOR2_X1 U585 ( .A(n485), .B(KEYINPUT22), .ZN(n486) );
  XNOR2_X1 U586 ( .A(n487), .B(n486), .ZN(n528) );
  XNOR2_X1 U587 ( .A(KEYINPUT4), .B(G131), .ZN(n489) );
  XNOR2_X1 U588 ( .A(G146), .B(n750), .ZN(n508) );
  NAND2_X1 U589 ( .A1(n490), .A2(G210), .ZN(n491) );
  XNOR2_X1 U590 ( .A(n492), .B(n491), .ZN(n495) );
  XOR2_X1 U591 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n494) );
  NOR2_X1 U592 ( .A1(G902), .A2(n644), .ZN(n498) );
  XNOR2_X1 U593 ( .A(G472), .B(KEYINPUT93), .ZN(n497) );
  XNOR2_X1 U594 ( .A(n498), .B(n497), .ZN(n603) );
  XNOR2_X1 U595 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n499) );
  XNOR2_X1 U596 ( .A(n603), .B(n499), .ZN(n614) );
  XNOR2_X1 U597 ( .A(KEYINPUT87), .B(n516), .ZN(n749) );
  XOR2_X1 U598 ( .A(n749), .B(n500), .Z(n504) );
  NAND2_X1 U599 ( .A1(G227), .A2(n459), .ZN(n505) );
  XNOR2_X1 U600 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U601 ( .A(n508), .B(n507), .ZN(n719) );
  NOR2_X1 U602 ( .A1(G902), .A2(n719), .ZN(n510) );
  XNOR2_X1 U603 ( .A(KEYINPUT68), .B(G469), .ZN(n509) );
  XNOR2_X2 U604 ( .A(n510), .B(n509), .ZN(n592) );
  NAND2_X1 U605 ( .A1(G221), .A2(n513), .ZN(n515) );
  INV_X1 U606 ( .A(n516), .ZN(n517) );
  XOR2_X1 U607 ( .A(n517), .B(KEYINPUT69), .Z(n518) );
  XNOR2_X1 U608 ( .A(n748), .B(KEYINPUT23), .ZN(n519) );
  NOR2_X1 U609 ( .A1(G902), .A2(n736), .ZN(n524) );
  NAND2_X1 U610 ( .A1(n520), .A2(G217), .ZN(n521) );
  XNOR2_X1 U611 ( .A(KEYINPUT74), .B(n521), .ZN(n522) );
  XNOR2_X1 U612 ( .A(n522), .B(KEYINPUT25), .ZN(n523) );
  XNOR2_X1 U613 ( .A(n524), .B(n523), .ZN(n535) );
  INV_X1 U614 ( .A(n535), .ZN(n589) );
  INV_X1 U615 ( .A(n589), .ZN(n685) );
  NOR2_X1 U616 ( .A1(n689), .A2(n685), .ZN(n525) );
  AND2_X1 U617 ( .A1(n614), .A2(n525), .ZN(n526) );
  NAND2_X1 U618 ( .A1(n528), .A2(n526), .ZN(n527) );
  INV_X1 U619 ( .A(n603), .ZN(n688) );
  INV_X1 U620 ( .A(n688), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n561), .A2(n685), .ZN(n529) );
  AND2_X2 U622 ( .A1(n549), .A2(n529), .ZN(n659) );
  INV_X1 U623 ( .A(n659), .ZN(n530) );
  XNOR2_X2 U624 ( .A(n532), .B(KEYINPUT81), .ZN(n570) );
  INV_X1 U625 ( .A(KEYINPUT71), .ZN(n533) );
  AND2_X1 U626 ( .A1(n533), .A2(KEYINPUT44), .ZN(n534) );
  INV_X1 U627 ( .A(n614), .ZN(n536) );
  INV_X1 U628 ( .A(n588), .ZN(n684) );
  NAND2_X1 U629 ( .A1(n535), .A2(n684), .ZN(n690) );
  NAND2_X1 U630 ( .A1(n536), .A2(n553), .ZN(n538) );
  XOR2_X1 U631 ( .A(KEYINPUT82), .B(KEYINPUT33), .Z(n537) );
  XNOR2_X1 U632 ( .A(n538), .B(n537), .ZN(n680) );
  NOR2_X1 U633 ( .A1(n680), .A2(n558), .ZN(n540) );
  XNOR2_X1 U634 ( .A(n540), .B(KEYINPUT34), .ZN(n541) );
  AND2_X1 U635 ( .A1(n552), .A2(n550), .ZN(n608) );
  NAND2_X1 U636 ( .A1(n541), .A2(n608), .ZN(n542) );
  XNOR2_X2 U637 ( .A(n542), .B(KEYINPUT35), .ZN(n761) );
  NAND2_X1 U638 ( .A1(n761), .A2(KEYINPUT80), .ZN(n543) );
  NAND2_X1 U639 ( .A1(n544), .A2(n543), .ZN(n547) );
  INV_X1 U640 ( .A(KEYINPUT44), .ZN(n545) );
  NAND2_X1 U641 ( .A1(n545), .A2(KEYINPUT80), .ZN(n546) );
  NAND2_X1 U642 ( .A1(n547), .A2(n546), .ZN(n567) );
  AND2_X1 U643 ( .A1(n614), .A2(n685), .ZN(n548) );
  AND2_X1 U644 ( .A1(n549), .A2(n548), .ZN(n650) );
  XNOR2_X1 U645 ( .A(n551), .B(KEYINPUT101), .ZN(n655) );
  INV_X1 U646 ( .A(n668), .ZN(n625) );
  NAND2_X1 U647 ( .A1(n655), .A2(n625), .ZN(n583) );
  INV_X1 U648 ( .A(n583), .ZN(n706) );
  AND2_X1 U649 ( .A1(n553), .A2(n561), .ZN(n694) );
  INV_X1 U650 ( .A(n558), .ZN(n554) );
  NAND2_X1 U651 ( .A1(n694), .A2(n554), .ZN(n555) );
  XNOR2_X1 U652 ( .A(n555), .B(KEYINPUT31), .ZN(n671) );
  NOR2_X1 U653 ( .A1(n592), .A2(n690), .ZN(n557) );
  XNOR2_X1 U654 ( .A(n557), .B(n556), .ZN(n620) );
  NOR2_X1 U655 ( .A1(n620), .A2(n558), .ZN(n559) );
  XNOR2_X1 U656 ( .A(n559), .B(KEYINPUT91), .ZN(n560) );
  NOR2_X1 U657 ( .A1(n561), .A2(n560), .ZN(n656) );
  NOR2_X1 U658 ( .A1(n671), .A2(n656), .ZN(n562) );
  NOR2_X1 U659 ( .A1(n706), .A2(n562), .ZN(n563) );
  OR2_X1 U660 ( .A1(n650), .A2(n563), .ZN(n565) );
  INV_X1 U661 ( .A(KEYINPUT104), .ZN(n564) );
  XNOR2_X1 U662 ( .A(n565), .B(n564), .ZN(n566) );
  INV_X1 U663 ( .A(n761), .ZN(n572) );
  NAND2_X1 U664 ( .A1(n572), .A2(n570), .ZN(n568) );
  NAND2_X1 U665 ( .A1(n568), .A2(KEYINPUT71), .ZN(n575) );
  NOR2_X1 U666 ( .A1(KEYINPUT44), .A2(KEYINPUT71), .ZN(n569) );
  NAND2_X1 U667 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U668 ( .A1(n571), .A2(KEYINPUT80), .ZN(n573) );
  NAND2_X1 U669 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U670 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U671 ( .A1(KEYINPUT2), .A2(KEYINPUT77), .ZN(n579) );
  NOR2_X1 U672 ( .A1(n580), .A2(n579), .ZN(n638) );
  INV_X1 U673 ( .A(n638), .ZN(n582) );
  AND2_X1 U674 ( .A1(n583), .A2(n598), .ZN(n595) );
  NOR2_X1 U675 ( .A1(G900), .A2(n459), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n584), .A2(G902), .ZN(n586) );
  NAND2_X1 U677 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U678 ( .A1(n587), .A2(n683), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n588), .A2(n607), .ZN(n590) );
  NAND2_X1 U680 ( .A1(n590), .A2(n589), .ZN(n615) );
  XNOR2_X1 U681 ( .A(n591), .B(KEYINPUT28), .ZN(n594) );
  INV_X1 U682 ( .A(n592), .ZN(n593) );
  NAND2_X1 U683 ( .A1(n595), .A2(n629), .ZN(n596) );
  NAND2_X1 U684 ( .A1(n596), .A2(KEYINPUT76), .ZN(n597) );
  XNOR2_X1 U685 ( .A(n597), .B(KEYINPUT47), .ZN(n602) );
  INV_X1 U686 ( .A(KEYINPUT76), .ZN(n600) );
  NAND2_X1 U687 ( .A1(n629), .A2(n598), .ZN(n660) );
  NAND2_X1 U688 ( .A1(n660), .A2(n583), .ZN(n599) );
  NAND2_X1 U689 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U690 ( .A1(n602), .A2(n601), .ZN(n612) );
  AND2_X1 U691 ( .A1(n603), .A2(n701), .ZN(n605) );
  INV_X1 U692 ( .A(KEYINPUT30), .ZN(n604) );
  XNOR2_X1 U693 ( .A(n605), .B(n604), .ZN(n606) );
  OR2_X1 U694 ( .A1(n607), .A2(n606), .ZN(n622) );
  NOR2_X1 U695 ( .A1(n622), .A2(n620), .ZN(n609) );
  NAND2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n611) );
  XOR2_X1 U697 ( .A(KEYINPUT73), .B(n613), .Z(n619) );
  INV_X1 U698 ( .A(n689), .ZN(n635) );
  XNOR2_X1 U699 ( .A(n616), .B(KEYINPUT36), .ZN(n617) );
  AND2_X1 U700 ( .A1(n635), .A2(n617), .ZN(n676) );
  XNOR2_X1 U701 ( .A(KEYINPUT79), .B(n676), .ZN(n618) );
  INV_X1 U702 ( .A(n702), .ZN(n621) );
  OR2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n624), .B(KEYINPUT39), .ZN(n631) );
  NOR2_X1 U705 ( .A1(n631), .A2(n625), .ZN(n627) );
  XNOR2_X1 U706 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n626) );
  XNOR2_X1 U707 ( .A(n627), .B(n626), .ZN(n760) );
  NAND2_X1 U708 ( .A1(n702), .A2(n701), .ZN(n707) );
  XNOR2_X1 U709 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n628) );
  XOR2_X1 U710 ( .A(KEYINPUT42), .B(n630), .Z(n762) );
  NOR2_X1 U711 ( .A1(n631), .A2(n655), .ZN(n632) );
  XNOR2_X1 U712 ( .A(n632), .B(KEYINPUT109), .ZN(n759) );
  XOR2_X1 U713 ( .A(KEYINPUT105), .B(n633), .Z(n634) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  AND2_X1 U715 ( .A1(n759), .A2(n677), .ZN(n637) );
  INV_X1 U716 ( .A(KEYINPUT2), .ZN(n641) );
  NOR2_X1 U717 ( .A1(n641), .A2(KEYINPUT77), .ZN(n639) );
  OR2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n640) );
  INV_X1 U719 ( .A(G952), .ZN(n645) );
  AND2_X1 U720 ( .A1(n645), .A2(G953), .ZN(n737) );
  XOR2_X1 U721 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n647) );
  XNOR2_X1 U722 ( .A(KEYINPUT55), .B(KEYINPUT75), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(n648) );
  XOR2_X1 U724 ( .A(G101), .B(n650), .Z(G3) );
  NAND2_X1 U725 ( .A1(n668), .A2(n656), .ZN(n651) );
  XNOR2_X1 U726 ( .A(G104), .B(n651), .ZN(G6) );
  XOR2_X1 U727 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n653) );
  XNOR2_X1 U728 ( .A(G107), .B(KEYINPUT26), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U730 ( .A(KEYINPUT110), .B(n654), .Z(n658) );
  INV_X1 U731 ( .A(n655), .ZN(n670) );
  NAND2_X1 U732 ( .A1(n656), .A2(n670), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n658), .B(n657), .ZN(G9) );
  XOR2_X1 U734 ( .A(n659), .B(G110), .Z(G12) );
  XOR2_X1 U735 ( .A(G128), .B(KEYINPUT29), .Z(n662) );
  INV_X1 U736 ( .A(n660), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n666), .A2(n670), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n662), .B(n661), .ZN(G30) );
  XNOR2_X1 U739 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U740 ( .A(KEYINPUT112), .B(n665), .ZN(G45) );
  NAND2_X1 U741 ( .A1(n666), .A2(n668), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n667), .B(G146), .ZN(G48) );
  NAND2_X1 U743 ( .A1(n671), .A2(n668), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n669), .B(G113), .ZN(G15) );
  NAND2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n672), .B(G116), .ZN(G18) );
  XOR2_X1 U747 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n674) );
  XNOR2_X1 U748 ( .A(G125), .B(KEYINPUT37), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U750 ( .A(n676), .B(n675), .ZN(G27) );
  XOR2_X1 U751 ( .A(G140), .B(n677), .Z(n678) );
  XNOR2_X1 U752 ( .A(n678), .B(KEYINPUT115), .ZN(G42) );
  XOR2_X1 U753 ( .A(KEYINPUT2), .B(n679), .Z(n682) );
  INV_X1 U754 ( .A(n698), .ZN(n681) );
  NAND2_X1 U755 ( .A1(G952), .A2(n683), .ZN(n716) );
  NOR2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT49), .ZN(n687) );
  NAND2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n693) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U760 ( .A(KEYINPUT50), .B(n691), .Z(n692) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n695) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U763 ( .A(n696), .B(KEYINPUT51), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n697), .B(KEYINPUT116), .ZN(n699) );
  NAND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U766 ( .A(n700), .B(KEYINPUT117), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n705), .B(KEYINPUT118), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U772 ( .A1(n680), .A2(n710), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U774 ( .A(KEYINPUT52), .B(n713), .Z(n714) );
  XNOR2_X1 U775 ( .A(KEYINPUT119), .B(n714), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U777 ( .A1(G953), .A2(n717), .ZN(n718) );
  NAND2_X1 U778 ( .A1(n731), .A2(G469), .ZN(n723) );
  XNOR2_X1 U779 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n721) );
  XNOR2_X1 U780 ( .A(n719), .B(KEYINPUT57), .ZN(n720) );
  XNOR2_X1 U781 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U782 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U783 ( .A1(n737), .A2(n724), .ZN(G54) );
  XOR2_X1 U784 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n725) );
  XNOR2_X1 U785 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U786 ( .A(KEYINPUT60), .B(n730), .ZN(G60) );
  NAND2_X1 U787 ( .A1(n731), .A2(G478), .ZN(n733) );
  XNOR2_X1 U788 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U789 ( .A1(n737), .A2(n734), .ZN(G63) );
  XOR2_X1 U790 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n735) );
  XNOR2_X1 U791 ( .A(n738), .B(G110), .ZN(n740) );
  NOR2_X1 U792 ( .A1(n740), .A2(n739), .ZN(n747) );
  XNOR2_X1 U793 ( .A(n741), .B(KEYINPUT126), .ZN(n745) );
  NAND2_X1 U794 ( .A1(G953), .A2(G224), .ZN(n742) );
  XNOR2_X1 U795 ( .A(KEYINPUT61), .B(n742), .ZN(n743) );
  NAND2_X1 U796 ( .A1(n743), .A2(G898), .ZN(n744) );
  NAND2_X1 U797 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(G69) );
  XNOR2_X1 U799 ( .A(n749), .B(n748), .ZN(n751) );
  XOR2_X1 U800 ( .A(n751), .B(n750), .Z(n754) );
  XOR2_X1 U801 ( .A(n754), .B(n752), .Z(n753) );
  NAND2_X1 U802 ( .A1(n753), .A2(n459), .ZN(n758) );
  XNOR2_X1 U803 ( .A(G227), .B(n754), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(G953), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n758), .A2(n757), .ZN(G72) );
  XNOR2_X1 U807 ( .A(G134), .B(n759), .ZN(G36) );
  XOR2_X1 U808 ( .A(n760), .B(G131), .Z(G33) );
  XOR2_X1 U809 ( .A(n761), .B(G122), .Z(G24) );
  XOR2_X1 U810 ( .A(G137), .B(n762), .Z(G39) );
endmodule

