//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(G104), .ZN(new_n189));
  INV_X1    g003(.A(G131), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT69), .A2(G237), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT69), .A2(G237), .ZN(new_n193));
  OAI211_X1 g007(.A(G214), .B(new_n191), .C1(new_n192), .C2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT83), .B(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT69), .B(G237), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT83), .A2(G143), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(G214), .A3(new_n191), .A4(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n190), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT18), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n196), .A2(new_n199), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT18), .A2(G131), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT84), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT84), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n212), .A3(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(KEYINPUT73), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n202), .A2(new_n203), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n200), .A2(KEYINPUT17), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n221));
  OR3_X1    g035(.A1(new_n206), .A2(KEYINPUT16), .A3(G140), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n221), .A2(G146), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(G146), .B1(new_n221), .B2(new_n222), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT86), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n222), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n217), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n222), .A3(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT86), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n220), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n196), .A2(new_n199), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT85), .B1(new_n232), .B2(G131), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(G131), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT85), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n196), .A2(new_n199), .A3(new_n236), .A4(new_n190), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n233), .A2(new_n234), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  AOI221_X4 g052(.A(new_n189), .B1(new_n201), .B2(new_n219), .C1(new_n231), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n189), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n231), .A2(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n219), .A2(new_n201), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n187), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G475), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT20), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n241), .A2(new_n240), .A3(new_n242), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n209), .A2(new_n212), .A3(KEYINPUT19), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT19), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n214), .A2(new_n216), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n250), .A3(new_n217), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n228), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n235), .A2(new_n237), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n233), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n219), .A2(new_n201), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n189), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(G475), .A2(G902), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n246), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n258), .ZN(new_n260));
  AOI211_X1 g074(.A(KEYINPUT20), .B(new_n260), .C1(new_n247), .C2(new_n256), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n245), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT9), .B(G234), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(G217), .A3(new_n191), .ZN(new_n265));
  INV_X1    g079(.A(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(G143), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OR3_X1    g083(.A1(new_n267), .A2(new_n269), .A3(G134), .ZN(new_n270));
  OAI21_X1  g084(.A(G134), .B1(new_n269), .B2(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G122), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G116), .ZN(new_n274));
  INV_X1    g088(.A(G116), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G122), .ZN(new_n276));
  INV_X1    g090(.A(G107), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT14), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n276), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n273), .A2(G116), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n279), .B2(new_n274), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT88), .B1(new_n276), .B2(KEYINPUT14), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n282), .B(G107), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n272), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n274), .A2(new_n276), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G107), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n278), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT13), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n266), .B2(G143), .ZN(new_n292));
  INV_X1    g106(.A(G143), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT13), .A3(G128), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n268), .A3(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n295), .A2(KEYINPUT87), .A3(G134), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT87), .B1(new_n295), .B2(G134), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n270), .B(new_n290), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT89), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n287), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n287), .B2(new_n298), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n265), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n287), .A2(new_n298), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT89), .ZN(new_n305));
  INV_X1    g119(.A(new_n265), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n300), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n187), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(G234), .A2(G237), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(G952), .A3(new_n191), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT21), .B(G898), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT90), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(G902), .A3(G953), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n311), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n308), .A2(new_n187), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n312), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n262), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G469), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n217), .A2(G143), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n293), .A2(G146), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n217), .A2(KEYINPUT64), .A3(G143), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT64), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n293), .B2(G146), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n293), .A2(G146), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n333));
  OAI21_X1  g147(.A(G128), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n327), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n277), .A2(KEYINPUT78), .A3(G104), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n337));
  INV_X1    g151(.A(G104), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(G107), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n277), .A2(G104), .ZN(new_n340));
  OAI211_X1 g154(.A(G101), .B(new_n336), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT3), .B1(new_n338), .B2(G107), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n277), .A3(G104), .ZN(new_n344));
  INV_X1    g158(.A(G101), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n338), .A2(G107), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n342), .A2(new_n344), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT10), .B1(new_n335), .B2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n341), .A2(new_n347), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n325), .A2(new_n326), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n266), .B1(new_n325), .B2(KEYINPUT1), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G101), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT77), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n362), .A3(G101), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(KEYINPUT0), .A2(G128), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT0), .A2(G128), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n332), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n358), .A2(new_n369), .A3(G101), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n353), .A2(new_n365), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G134), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT65), .B1(new_n374), .B2(G137), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT11), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT11), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT65), .B(new_n377), .C1(new_n374), .C2(G137), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(G137), .ZN(new_n379));
  AND4_X1   g193(.A1(new_n190), .A2(new_n376), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n375), .A2(KEYINPUT11), .B1(new_n374), .B2(G137), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n190), .B1(new_n381), .B2(new_n378), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n357), .A2(new_n373), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT79), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n349), .A2(new_n356), .B1(new_n364), .B2(new_n372), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G110), .B(G140), .ZN(new_n390));
  INV_X1    g204(.A(G227), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G953), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n390), .B(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n350), .A2(new_n355), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n335), .A2(new_n348), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n383), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT12), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT12), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n389), .A2(new_n394), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n357), .A2(new_n373), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n398), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n394), .B1(new_n389), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n323), .B(new_n187), .C1(new_n404), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n387), .B1(new_n386), .B2(new_n383), .ZN(new_n409));
  AND4_X1   g223(.A1(new_n387), .A2(new_n357), .A3(new_n373), .A4(new_n383), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n394), .B(new_n406), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n385), .A2(new_n388), .B1(new_n402), .B2(new_n401), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n411), .B(G469), .C1(new_n412), .C2(new_n394), .ZN(new_n413));
  NAND2_X1  g227(.A1(G469), .A2(G902), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G214), .B1(G237), .B2(G902), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G210), .B1(G237), .B2(G902), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT2), .B(G113), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G119), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT68), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G119), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n425), .A3(G116), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n275), .A2(G119), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n421), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n426), .A2(KEYINPUT5), .A3(new_n427), .ZN(new_n429));
  OAI21_X1  g243(.A(G113), .B1(new_n426), .B2(KEYINPUT5), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n350), .B(new_n428), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n427), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT67), .A3(new_n420), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n420), .B1(new_n432), .B2(KEYINPUT67), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n370), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n431), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n439), .B(new_n431), .C1(new_n436), .C2(new_n437), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n438), .A2(new_n444), .A3(new_n440), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n368), .A2(new_n371), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G125), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n335), .A2(new_n206), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n191), .A2(G224), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT80), .Z(new_n451));
  XNOR2_X1  g265(.A(new_n449), .B(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n443), .A2(new_n445), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n348), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n431), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT81), .B(KEYINPUT8), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n439), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT82), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n456), .A2(new_n461), .A3(new_n458), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n447), .A2(new_n448), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(new_n447), .B2(new_n448), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n460), .A2(new_n442), .A3(new_n462), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n187), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n419), .B1(new_n453), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n467), .A2(new_n442), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n456), .A2(new_n461), .A3(new_n458), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n461), .B1(new_n456), .B2(new_n458), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n443), .A2(new_n445), .A3(new_n452), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n418), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n417), .B1(new_n470), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G221), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n264), .B2(new_n187), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n322), .A2(new_n415), .A3(new_n478), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n413), .A2(new_n414), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n480), .B1(new_n485), .B2(new_n408), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n486), .A2(KEYINPUT91), .A3(new_n322), .A4(new_n478), .ZN(new_n487));
  INV_X1    g301(.A(G472), .ZN(new_n488));
  INV_X1    g302(.A(new_n435), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n433), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n332), .A2(new_n367), .B1(new_n365), .B2(new_n353), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n380), .B2(new_n382), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n381), .A2(new_n190), .A3(new_n378), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT66), .B1(new_n374), .B2(G137), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n379), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n374), .A2(KEYINPUT66), .A3(G137), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n326), .A2(KEYINPUT64), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n325), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n354), .B1(new_n499), .B2(new_n328), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n493), .B(new_n497), .C1(new_n500), .C2(new_n327), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n490), .B1(new_n502), .B2(KEYINPUT71), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n492), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT28), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n502), .A2(new_n490), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n434), .A2(new_n435), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n492), .A3(new_n501), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n197), .A2(G210), .A3(new_n191), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT26), .B(G101), .Z(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n506), .A2(new_n511), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n518), .B2(KEYINPUT29), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n502), .A2(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n509), .A3(new_n505), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n507), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n508), .A2(new_n510), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT28), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n492), .A2(new_n501), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n492), .B2(new_n501), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n490), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n510), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n517), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n488), .B1(new_n519), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n529), .A2(new_n510), .A3(new_n516), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n517), .B1(new_n506), .B2(new_n511), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n529), .A2(new_n538), .A3(new_n510), .A4(new_n516), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G472), .A2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT32), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(new_n544), .A3(new_n541), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n534), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT22), .B(G137), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT74), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n218), .A2(new_n228), .ZN(new_n551));
  NOR2_X1   g365(.A1(G119), .A2(G128), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT68), .B(G119), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT23), .B(new_n553), .C1(new_n554), .C2(new_n266), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n554), .B2(G128), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n266), .B1(new_n423), .B2(new_n425), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT24), .B(G110), .Z(new_n561));
  OR3_X1    g375(.A1(new_n560), .A2(new_n561), .A3(new_n552), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n551), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n561), .B1(new_n560), .B2(new_n552), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n223), .B2(new_n224), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n556), .B1(new_n555), .B2(new_n558), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n550), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n559), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n218), .A2(new_n228), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n227), .A2(new_n228), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n555), .A2(new_n558), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(new_n564), .C1(new_n573), .C2(new_n556), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n574), .A3(new_n549), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n575), .A3(new_n187), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT25), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(G217), .A2(G902), .ZN(new_n580));
  INV_X1    g394(.A(G217), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(G234), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT72), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n576), .A2(new_n577), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n568), .A2(new_n575), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n187), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(KEYINPUT76), .Z(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n546), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n484), .A2(new_n487), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT92), .B(G101), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G3));
  INV_X1    g412(.A(new_n594), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n486), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n470), .A2(new_n477), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n318), .A3(new_n416), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n308), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n303), .A2(new_n307), .A3(KEYINPUT33), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(G478), .A3(new_n187), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n309), .A2(new_n310), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n262), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n488), .B1(new_n540), .B2(new_n187), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n542), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n601), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NAND3_X1  g432(.A1(new_n233), .A2(new_n235), .A3(new_n237), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n228), .A3(new_n251), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n240), .B1(new_n620), .B2(new_n242), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n258), .B1(new_n239), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT20), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n257), .A2(new_n246), .A3(new_n258), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n623), .A2(new_n624), .B1(G475), .B2(new_n244), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n319), .B1(new_n308), .B2(new_n187), .ZN(new_n626));
  AOI211_X1 g440(.A(G902), .B(new_n311), .C1(new_n303), .C2(new_n307), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n603), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n601), .A2(new_n615), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  AOI21_X1  g448(.A(KEYINPUT25), .B1(new_n576), .B2(new_n577), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n578), .A2(new_n635), .A3(new_n583), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n550), .A2(KEYINPUT36), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n563), .A2(new_n567), .A3(KEYINPUT93), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT93), .B1(new_n563), .B2(new_n567), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n638), .A2(new_n637), .A3(new_n639), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n591), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT94), .B1(new_n636), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT94), .ZN(new_n645));
  INV_X1    g459(.A(new_n642), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n592), .B1(new_n646), .B2(new_n640), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n587), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n484), .A2(new_n487), .A3(new_n615), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  XNOR2_X1  g466(.A(new_n314), .B(KEYINPUT95), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(G900), .B2(new_n317), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n625), .A2(new_n629), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT96), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n486), .A2(new_n478), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n644), .A2(new_n648), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n546), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  NAND2_X1  g476(.A1(new_n523), .A2(new_n517), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT97), .ZN(new_n664));
  INV_X1    g478(.A(new_n535), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n187), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G472), .ZN(new_n667));
  INV_X1    g481(.A(new_n545), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n544), .B1(new_n540), .B2(new_n541), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT98), .Z(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n654), .B(KEYINPUT39), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n486), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n602), .B(KEYINPUT38), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n625), .A2(new_n628), .A3(new_n417), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n677), .A2(new_n659), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n672), .A2(new_n675), .A3(new_n676), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  INV_X1    g495(.A(new_n654), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n610), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n660), .A2(new_n658), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  INV_X1    g499(.A(new_n534), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n668), .B2(new_n669), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n393), .B1(new_n385), .B2(new_n388), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n393), .A2(new_n688), .B1(new_n689), .B2(new_n403), .ZN(new_n690));
  OAI21_X1  g504(.A(G469), .B1(new_n690), .B2(G902), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n691), .A2(new_n481), .A3(new_n408), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n687), .A2(new_n599), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n611), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT41), .B(G113), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND4_X1  g511(.A1(new_n631), .A2(new_n687), .A3(new_n599), .A4(new_n692), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  NAND2_X1  g513(.A1(new_n687), .A2(new_n649), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n692), .A2(new_n322), .A3(new_n478), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n422), .ZN(G21));
  INV_X1    g517(.A(KEYINPUT99), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n536), .A2(new_n537), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n539), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n536), .B2(new_n537), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n541), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n613), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n594), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n691), .A2(new_n481), .A3(new_n408), .ZN(new_n711));
  INV_X1    g525(.A(new_n318), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n623), .A2(new_n624), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n628), .B1(new_n714), .B2(new_n245), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT100), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n715), .A2(new_n478), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n716), .B1(new_n715), .B2(new_n478), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n710), .B(new_n713), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT101), .B(G122), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G24));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n709), .B2(new_n659), .ZN(new_n723));
  INV_X1    g537(.A(new_n510), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n502), .A2(KEYINPUT30), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n492), .A2(new_n501), .A3(new_n526), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n724), .B1(new_n727), .B2(new_n490), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n538), .B1(new_n728), .B2(new_n516), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n516), .B1(new_n522), .B2(new_n524), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT99), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n539), .A3(new_n705), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n612), .B1(new_n732), .B2(new_n541), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(KEYINPUT102), .A3(new_n649), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n723), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n453), .A2(new_n469), .A3(new_n419), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n418), .B1(new_n475), .B2(new_n476), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n416), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n711), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n735), .A2(new_n683), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NOR2_X1   g555(.A1(new_n602), .A2(new_n417), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n688), .A2(new_n393), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n389), .A2(new_n394), .A3(new_n403), .ZN(new_n745));
  AOI211_X1 g559(.A(G469), .B(G902), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n414), .B(KEYINPUT103), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n413), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT104), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n408), .A2(new_n750), .A3(new_n413), .A4(new_n747), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n481), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n743), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n749), .A2(KEYINPUT105), .A3(new_n481), .A4(new_n751), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n595), .A3(new_n683), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT106), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n752), .A2(new_n753), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n761), .A2(new_n755), .A3(new_n742), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(KEYINPUT42), .A3(new_n595), .A4(new_n683), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n756), .A2(new_n757), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NAND4_X1  g582(.A1(new_n754), .A2(new_n657), .A3(new_n595), .A4(new_n755), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  XNOR2_X1  g584(.A(new_n625), .B(KEYINPUT108), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(KEYINPUT43), .A3(new_n609), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT109), .Z(new_n773));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n774));
  INV_X1    g588(.A(new_n609), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n775), .B2(new_n262), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n614), .B(new_n649), .C1(new_n777), .C2(new_n778), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n780), .B2(new_n781), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n411), .B1(new_n412), .B2(new_n394), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n323), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n786), .B2(new_n785), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT107), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n747), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n746), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n481), .A3(new_n673), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n743), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n783), .A2(new_n784), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n481), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n793), .A2(KEYINPUT47), .A3(new_n481), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n683), .A2(new_n546), .A3(new_n594), .A4(new_n742), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT111), .Z(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  NOR2_X1   g620(.A1(new_n672), .A2(new_n594), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n677), .A2(new_n417), .A3(new_n480), .A4(new_n775), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n691), .A2(new_n408), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT49), .Z(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(new_n771), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n653), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n777), .A2(new_n812), .A3(new_n710), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n677), .A2(new_n416), .A3(new_n711), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(KEYINPUT50), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n777), .A2(new_n812), .A3(new_n710), .A4(new_n814), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n743), .A2(new_n711), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n777), .A2(new_n812), .A3(new_n735), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n314), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n807), .A2(new_n822), .A3(new_n820), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n775), .A2(new_n625), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT119), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n813), .A2(new_n742), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n800), .B(new_n801), .C1(new_n481), .C2(new_n809), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n825), .B1(new_n815), .B2(new_n818), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n777), .A2(new_n595), .A3(new_n812), .A4(new_n820), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT48), .ZN(new_n838));
  OAI211_X1 g652(.A(G952), .B(new_n191), .C1(new_n823), .C2(new_n610), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n739), .B2(new_n813), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n838), .A2(new_n840), .A3(KEYINPUT122), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n835), .A2(new_n836), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n832), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n836), .B1(new_n829), .B2(new_n830), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n832), .B2(new_n847), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n846), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n827), .A2(KEYINPUT120), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT121), .A3(new_n848), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n845), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n658), .B(new_n660), .C1(new_n657), .C2(new_n683), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n715), .A2(new_n478), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT100), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n715), .A2(new_n478), .A3(new_n716), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n752), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n636), .A2(new_n643), .A3(new_n682), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n861), .A2(new_n670), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n740), .A2(new_n857), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n865), .A2(KEYINPUT52), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(KEYINPUT115), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n740), .A2(new_n857), .A3(new_n864), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT53), .B1(new_n758), .B2(new_n759), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n717), .A2(new_n718), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n713), .A2(new_n599), .A3(new_n733), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n698), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n693), .A2(new_n694), .B1(new_n700), .B2(new_n701), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n735), .A2(new_n683), .A3(new_n755), .A4(new_n754), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n629), .A2(new_n262), .A3(new_n682), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n660), .A2(new_n486), .A3(new_n742), .A4(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(new_n769), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n596), .A2(new_n616), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT112), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n630), .A2(KEYINPUT113), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n625), .B2(new_n629), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n603), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n601), .A3(new_n889), .A4(new_n615), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n650), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT112), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n596), .A2(new_n616), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n873), .A2(new_n882), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n872), .A2(KEYINPUT117), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT117), .B1(new_n872), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n546), .A2(new_n594), .A3(new_n711), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n714), .A2(new_n628), .A3(new_n245), .A4(new_n318), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n711), .A2(new_n738), .A3(new_n900), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n899), .A2(new_n611), .B1(new_n660), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(new_n698), .A3(new_n719), .A4(new_n881), .ZN(new_n903));
  INV_X1    g717(.A(new_n769), .ZN(new_n904));
  AND4_X1   g718(.A1(KEYINPUT102), .A2(new_n649), .A3(new_n613), .A4(new_n708), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT102), .B1(new_n733), .B2(new_n649), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n683), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n761), .A2(new_n755), .A3(new_n742), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n596), .A2(new_n892), .A3(new_n616), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n892), .B1(new_n596), .B2(new_n616), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n650), .A2(new_n890), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n760), .A2(new_n910), .A3(new_n766), .A4(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT114), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n867), .A2(KEYINPUT52), .A3(new_n869), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT52), .B1(new_n867), .B2(new_n869), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n882), .A2(new_n894), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(KEYINPUT114), .A3(new_n760), .A4(new_n766), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n898), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n917), .A2(new_n920), .A3(new_n922), .A4(KEYINPUT53), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(KEYINPUT116), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n917), .A2(new_n922), .A3(new_n872), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n924), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n933), .B2(new_n928), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n934), .B2(new_n926), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT118), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n927), .C1(new_n934), .C2(new_n926), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n856), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(G952), .A2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n811), .B1(new_n939), .B2(new_n940), .ZN(G75));
  NOR2_X1   g755(.A1(new_n191), .A2(G952), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n187), .B1(new_n898), .B2(new_n925), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT56), .B1(new_n944), .B2(G210), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n443), .A2(new_n445), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n452), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n943), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n945), .B2(new_n948), .ZN(G51));
  NAND2_X1  g764(.A1(new_n898), .A2(new_n925), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n927), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n747), .B(KEYINPUT57), .Z(new_n954));
  AOI21_X1  g768(.A(new_n690), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n789), .ZN(new_n956));
  AOI22_X1  g770(.A1(new_n955), .A2(KEYINPUT123), .B1(new_n956), .B2(new_n944), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n953), .A2(new_n954), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n690), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n942), .B1(new_n957), .B2(new_n960), .ZN(G54));
  NAND2_X1  g775(.A1(KEYINPUT58), .A2(G475), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT124), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n944), .A2(new_n257), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n257), .B1(new_n944), .B2(new_n963), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n966), .A2(new_n967), .A3(new_n942), .A4(new_n968), .ZN(G60));
  AND2_X1   g783(.A1(new_n605), .A2(new_n606), .ZN(new_n970));
  NAND2_X1  g784(.A1(G478), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT59), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n953), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n943), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n936), .A2(new_n938), .A3(new_n972), .ZN(new_n975));
  INV_X1    g789(.A(new_n970), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G63));
  XNOR2_X1  g791(.A(new_n580), .B(KEYINPUT60), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n898), .B2(new_n925), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n646), .B2(new_n640), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n980), .B(new_n943), .C1(new_n589), .C2(new_n979), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g796(.A(new_n191), .B1(new_n316), .B2(G224), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n914), .A2(new_n878), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n191), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n946), .B1(G898), .B2(new_n191), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n985), .B(new_n986), .Z(G69));
  AND2_X1   g801(.A1(new_n740), .A2(new_n857), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n680), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n610), .B1(new_n885), .B2(new_n887), .ZN(new_n991));
  NOR4_X1   g805(.A1(new_n674), .A2(new_n743), .A3(new_n546), .A4(new_n594), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n796), .A2(new_n993), .A3(new_n805), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n191), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n248), .A2(new_n250), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n727), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n191), .A2(G900), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n796), .A2(new_n805), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n988), .A2(new_n769), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n861), .A2(new_n595), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n767), .B(new_n1002), .C1(new_n794), .C2(new_n1003), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1000), .B1(new_n1005), .B2(new_n191), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n999), .B1(new_n1006), .B2(new_n998), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1000), .B1(new_n391), .B2(G953), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT126), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1009), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1011), .B(new_n999), .C1(new_n1006), .C2(new_n998), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n995), .B2(new_n984), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n728), .B(KEYINPUT127), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1016), .A2(new_n516), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1015), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1020));
  INV_X1    g834(.A(new_n984), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OR2_X1    g836(.A1(new_n1017), .A2(new_n516), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1018), .B(new_n943), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n934), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1019), .B1(new_n531), .B2(new_n535), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(G57));
endmodule


