//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1191,
    new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n465), .B1(new_n470), .B2(G137), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n463), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI211_X1 g053(.A(KEYINPUT69), .B(new_n463), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(G160));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n463), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(G136), .B2(new_n470), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT70), .Z(G162));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND2_X1  g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n468), .B2(new_n469), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n463), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n489), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n490), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n472), .B2(new_n473), .ZN(new_n497));
  INV_X1    g072(.A(G102), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(new_n463), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(new_n501), .A3(G2104), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n497), .A2(new_n502), .A3(KEYINPUT71), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n463), .C1(new_n472), .C2(new_n473), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n481), .A2(new_n506), .A3(G138), .A4(new_n463), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n495), .A2(new_n503), .B1(new_n505), .B2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(G543), .A3(new_n515), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(new_n509), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n518), .A2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(G51), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(G651), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n532), .A2(G63), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n527), .A2(new_n528), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n509), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT73), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT74), .B(G90), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n542), .A2(new_n520), .B1(new_n517), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n518), .A2(G81), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n521), .A2(G43), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n509), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  AOI22_X1  g131(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT75), .B1(new_n557), .B2(new_n509), .ZN(new_n558));
  OAI21_X1  g133(.A(G65), .B1(new_n529), .B2(new_n530), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(new_n562), .A3(G651), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n558), .A2(new_n563), .B1(new_n518), .B2(G91), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n514), .A2(G53), .A3(G543), .A4(new_n515), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n510), .A2(new_n513), .B1(KEYINPUT6), .B2(new_n509), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n567), .A2(new_n568), .A3(G53), .A4(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n564), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n573), .B(G651), .C1(new_n516), .C2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(G74), .A2(G651), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n531), .A2(KEYINPUT76), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n514), .A2(G49), .A3(G543), .A4(new_n515), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n514), .A2(G87), .A3(new_n515), .A4(new_n516), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OR2_X1    g156(.A1(KEYINPUT5), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(KEYINPUT5), .A2(G543), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(G73), .A2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT77), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n588), .B(G651), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n514), .A2(G48), .A3(G543), .A4(new_n515), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n514), .A2(G86), .A3(new_n515), .A4(new_n516), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n518), .A2(G85), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n521), .A2(G47), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n595), .B(new_n596), .C1(new_n509), .C2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n518), .A2(G92), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT10), .Z(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n520), .A2(new_n602), .B1(new_n603), .B2(new_n509), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT78), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n599), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n599), .B1(new_n607), .B2(G868), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G299), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NOR2_X1   g190(.A1(new_n551), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n607), .A2(new_n614), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT79), .Z(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n470), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n463), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(G123), .ZN(new_n624));
  OAI221_X1 g199(.A(new_n621), .B1(new_n622), .B2(new_n623), .C1(new_n624), .C2(new_n482), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n626), .A2(new_n631), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT80), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G1341), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G14), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n642), .A2(new_n646), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT17), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT81), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  INV_X1    g233(.A(new_n651), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n655), .C1(new_n659), .C2(new_n653), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n653), .A3(new_n654), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n670), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AOI211_X1 g250(.A(new_n672), .B(new_n675), .C1(new_n667), .C2(new_n671), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT83), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT84), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n678), .B(new_n684), .ZN(G229));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT32), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(G1981), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1971), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT33), .B(G1976), .ZN(new_n693));
  OR2_X1    g268(.A1(G16), .A2(G23), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n574), .A2(new_n576), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n578), .A2(new_n579), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n577), .A2(KEYINPUT89), .A3(new_n578), .A4(new_n579), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(new_n689), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n692), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n693), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n687), .A2(G1981), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n688), .A2(new_n702), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  MUX2_X1   g283(.A(G24), .B(G290), .S(G16), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT86), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n470), .A2(G131), .ZN(new_n716));
  INV_X1    g291(.A(G119), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n482), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n715), .A2(new_n718), .A3(KEYINPUT87), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT87), .B1(new_n715), .B2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n712), .B1(new_n722), .B2(new_n711), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n710), .B(new_n726), .C1(new_n727), .C2(KEYINPUT36), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n707), .A2(new_n708), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n727), .A2(KEYINPUT36), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT24), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n711), .B1(new_n734), .B2(G34), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n734), .B2(G34), .ZN(new_n738));
  AOI22_X1  g313(.A1(G160), .A2(G29), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n711), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n711), .ZN(new_n743));
  INV_X1    g318(.A(G2078), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n741), .B1(KEYINPUT99), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G5), .A2(G16), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT98), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G301), .B2(new_n689), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n746), .B(new_n751), .C1(KEYINPUT99), .C2(new_n745), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n711), .A2(G33), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n481), .A2(G127), .ZN(new_n754));
  INV_X1    g329(.A(G115), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(new_n467), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n463), .B1(new_n756), .B2(KEYINPUT94), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(KEYINPUT94), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n470), .A2(G139), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n753), .B1(new_n762), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2072), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n689), .A2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G168), .B2(new_n689), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n765), .B1(G1966), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G1966), .B2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n711), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G116), .B2(new_n463), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT92), .ZN(new_n775));
  INV_X1    g350(.A(new_n482), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n776), .A2(G128), .B1(G140), .B2(new_n470), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(new_n711), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT93), .B(G2067), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n779), .B(new_n780), .Z(new_n781));
  INV_X1    g356(.A(G28), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT30), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n782), .B2(KEYINPUT30), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n781), .B(new_n787), .C1(new_n711), .C2(new_n625), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n711), .A2(G32), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n776), .A2(G129), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT97), .ZN(new_n791));
  AND3_X1   g366(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT26), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n792), .B(new_n794), .C1(G141), .C2(new_n470), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(new_n711), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT27), .B(G1996), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G16), .A2(G19), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n551), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1341), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n769), .A2(new_n788), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n711), .A2(G35), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G162), .B2(new_n711), .ZN(new_n806));
  INV_X1    g381(.A(G2090), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n752), .A2(new_n804), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n607), .A2(new_n689), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G4), .B2(new_n689), .ZN(new_n813));
  INV_X1    g388(.A(G1348), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n689), .A2(G20), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT23), .Z(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G299), .B2(G16), .ZN(new_n818));
  INV_X1    g393(.A(G1956), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n763), .A2(new_n764), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT95), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n813), .B2(new_n814), .ZN(new_n823));
  NOR4_X1   g398(.A1(new_n811), .A2(new_n815), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n732), .A2(new_n733), .A3(new_n825), .ZN(G311));
  INV_X1    g401(.A(G311), .ZN(G150));
  NAND2_X1  g402(.A1(new_n607), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n830), .A2(new_n520), .B1(new_n517), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n516), .A2(G67), .ZN(new_n835));
  AND2_X1   g410(.A1(G80), .A2(G543), .ZN(new_n836));
  OAI21_X1  g411(.A(G651), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n550), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n829), .B(new_n839), .Z(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n841), .A2(new_n842), .A3(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n838), .A2(G860), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n491), .B2(new_n494), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n497), .A2(new_n502), .A3(KEYINPUT102), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n506), .B1(new_n470), .B2(G138), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n778), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n762), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n797), .ZN(new_n855));
  INV_X1    g430(.A(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n463), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n482), .A2(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G142), .B2(new_n470), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(new_n628), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n721), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G162), .B(new_n625), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(G160), .Z(new_n865));
  XOR2_X1   g440(.A(new_n862), .B(KEYINPUT103), .Z(new_n866));
  OAI211_X1 g441(.A(new_n863), .B(new_n865), .C1(new_n855), .C2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n866), .B(new_n855), .Z(new_n869));
  OAI211_X1 g444(.A(new_n867), .B(new_n868), .C1(new_n869), .C2(new_n865), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g446(.A(new_n606), .B(G299), .Z(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT41), .Z(new_n873));
  XOR2_X1   g448(.A(new_n839), .B(new_n617), .Z(new_n874));
  MUX2_X1   g449(.A(new_n872), .B(new_n873), .S(new_n874), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n700), .B(G305), .ZN(new_n876));
  XNOR2_X1  g451(.A(G166), .B(G290), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n875), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G868), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n838), .A2(new_n610), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(G331));
  NAND2_X1  g464(.A1(G331), .A2(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(G295));
  XNOR2_X1  g468(.A(new_n839), .B(G286), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G171), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n839), .B(G168), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G301), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n872), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n873), .A2(new_n895), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n898), .B2(new_n872), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n878), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n872), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT107), .ZN(new_n906));
  INV_X1    g481(.A(new_n878), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n901), .A4(new_n900), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n904), .A2(new_n908), .A3(new_n909), .A4(new_n868), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n901), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n911), .B2(new_n878), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(new_n908), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n910), .B(KEYINPUT44), .C1(new_n913), .C2(new_n909), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n908), .A2(new_n909), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n904), .A2(new_n868), .A3(new_n908), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n912), .A2(new_n915), .B1(new_n916), .B2(KEYINPUT43), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n918));
  OAI21_X1  g493(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(G397));
  XOR2_X1   g494(.A(KEYINPUT108), .B(G40), .Z(new_n920));
  NOR3_X1   g495(.A1(new_n478), .A2(new_n479), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1384), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n852), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n778), .B(G2067), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT110), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n928), .B2(new_n796), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n925), .A2(G1996), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT46), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n930), .A2(KEYINPUT46), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n928), .B1(G1996), .B2(new_n796), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n935), .A2(new_n925), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n797), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT109), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n722), .A2(new_n724), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n721), .A2(new_n725), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n926), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n925), .A2(G1986), .A3(G290), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT48), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n934), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n939), .A2(new_n941), .ZN(new_n947));
  INV_X1    g522(.A(G2067), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n778), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n925), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n505), .A2(new_n507), .ZN(new_n953));
  INV_X1    g528(.A(new_n503), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT71), .B1(new_n497), .B2(new_n502), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(KEYINPUT45), .A3(new_n922), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n497), .A2(new_n502), .A3(KEYINPUT102), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT102), .B1(new_n497), .B2(new_n502), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n960), .B2(new_n953), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n957), .B(new_n921), .C1(new_n961), .C2(KEYINPUT45), .ZN(new_n962));
  INV_X1    g537(.A(G1966), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  AND4_X1   g541(.A1(new_n965), .A2(new_n852), .A3(new_n966), .A4(new_n922), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n961), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n921), .A2(new_n740), .ZN(new_n971));
  OAI211_X1 g546(.A(G168), .B(new_n964), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n852), .A2(new_n966), .A3(new_n922), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n973), .A3(KEYINPUT112), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n961), .A2(new_n965), .A3(new_n966), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n475), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n481), .B2(G125), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT69), .B1(new_n978), .B2(new_n463), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n474), .A2(new_n475), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n477), .A3(G2105), .ZN(new_n981));
  INV_X1    g556(.A(new_n920), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n979), .A2(new_n981), .A3(new_n471), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n923), .B2(new_n924), .ZN(new_n984));
  AOI21_X1  g559(.A(G1966), .B1(new_n984), .B2(new_n957), .ZN(new_n985));
  OAI21_X1  g560(.A(G286), .B1(new_n976), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n972), .A2(new_n986), .A3(G8), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT51), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT62), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n974), .A2(new_n975), .ZN(new_n991));
  INV_X1    g566(.A(new_n971), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n991), .A2(new_n992), .B1(new_n963), .B2(new_n962), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n993), .B2(G168), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n988), .A2(new_n989), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n924), .B1(G164), .B2(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n922), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n921), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n998), .A2(new_n999), .A3(new_n921), .A4(KEYINPUT111), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n744), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n983), .B1(new_n974), .B2(new_n975), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1006), .A2(G2078), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI22_X1  g585(.A1(new_n1008), .A2(G1961), .B1(new_n962), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(G301), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n590), .A2(new_n1015), .A3(new_n593), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n590), .B2(new_n593), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT49), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n990), .B1(new_n921), .B2(new_n961), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1014), .B(new_n1021), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n698), .A2(G1976), .A3(new_n699), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1020), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1029), .B(new_n1030), .C1(new_n1020), .C2(new_n1024), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n921), .A2(new_n961), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n1024), .A3(G8), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT114), .B1(new_n1033), .B2(KEYINPUT52), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1971), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1002), .A2(new_n1037), .A3(new_n1003), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n495), .A2(new_n503), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1384), .B1(new_n1039), .B2(new_n953), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n983), .B1(new_n1040), .B2(new_n966), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n923), .A2(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n807), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G303), .A2(G8), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1008), .A2(new_n807), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n990), .B1(new_n1054), .B2(new_n1038), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1051), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1013), .A2(new_n1036), .A3(new_n1053), .A4(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n952), .B1(new_n997), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1038), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1059), .A2(G8), .A3(new_n1051), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1051), .B1(new_n1044), .B2(G8), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1023), .B(new_n1027), .C1(new_n1034), .C2(new_n1031), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n988), .A2(new_n989), .A3(new_n996), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(KEYINPUT125), .A4(new_n1013), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n995), .B1(new_n994), .B2(new_n986), .ZN(new_n1066));
  AOI211_X1 g641(.A(KEYINPUT51), .B(new_n990), .C1(new_n993), .C2(G168), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT62), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1058), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n750), .B1(new_n970), .B2(new_n983), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n923), .A2(new_n924), .ZN(new_n1071));
  INV_X1    g646(.A(new_n476), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n470), .A2(G137), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n464), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n471), .A2(KEYINPUT122), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1009), .A2(G40), .ZN(new_n1078));
  AND4_X1   g653(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1071), .A2(new_n1079), .A3(new_n999), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT123), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1071), .A2(new_n1079), .A3(new_n1082), .A4(new_n999), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G2078), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1070), .B(new_n1084), .C1(KEYINPUT53), .C2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT124), .B1(new_n1086), .B2(G171), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(KEYINPUT53), .ZN(new_n1088));
  OAI21_X1  g663(.A(G171), .B1(new_n1088), .B2(new_n1011), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1008), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1090), .A2(new_n750), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1007), .A2(new_n1091), .A3(new_n1092), .A4(G301), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1087), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n566), .A2(new_n569), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n567), .A2(G91), .A3(new_n516), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n562), .B1(new_n561), .B2(G651), .ZN(new_n1099));
  AOI211_X1 g674(.A(KEYINPUT75), .B(new_n509), .C1(new_n559), .C2(new_n560), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT119), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n570), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n564), .A2(new_n1105), .A3(new_n570), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1104), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1956), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  AND4_X1   g685(.A1(new_n921), .A2(new_n998), .A3(new_n999), .A4(new_n1110), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1107), .A2(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1104), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1097), .A2(new_n1101), .A3(KEYINPUT119), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1105), .B1(new_n564), .B2(new_n570), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n956), .A2(new_n966), .A3(new_n922), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n921), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n966), .B1(new_n852), .B2(new_n922), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n819), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1102), .A2(new_n1106), .A3(new_n1104), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n998), .A2(new_n999), .A3(new_n921), .A4(new_n1110), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1116), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1112), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n923), .A2(new_n983), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT58), .B(G1341), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1000), .A2(G1996), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n551), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT59), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1131), .A3(new_n551), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1124), .A2(new_n1125), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1112), .A2(KEYINPUT120), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n1139));
  OAI221_X1 g714(.A(new_n1139), .B1(new_n1109), .B2(new_n1111), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1126), .A2(new_n948), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1008), .B2(G1348), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT60), .B(new_n1142), .C1(new_n1008), .C2(G1348), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n607), .A3(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1133), .A2(new_n1141), .A3(new_n1145), .A4(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1138), .B(new_n1140), .C1(new_n606), .C2(new_n1144), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1123), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1036), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1086), .A2(G171), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1007), .A2(new_n1012), .A3(G301), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(KEYINPUT54), .A3(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1096), .A2(new_n1153), .A3(new_n1156), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(G288), .A2(G1976), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT116), .Z(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1020), .B1(new_n1163), .B2(new_n1016), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1036), .B(KEYINPUT117), .C1(new_n1051), .C2(new_n1055), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n993), .A2(new_n990), .A3(G286), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1056), .A2(KEYINPUT63), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1055), .A2(new_n1051), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1169), .B1(new_n1170), .B2(new_n1062), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1166), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1036), .A2(new_n1053), .A3(new_n1056), .A4(new_n1167), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1165), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1069), .A2(new_n1160), .A3(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(G290), .B(G1986), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n943), .B1(new_n926), .B2(new_n1178), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1177), .A2(KEYINPUT126), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT126), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n951), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(KEYINPUT127), .B(new_n951), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g761(.A1(G229), .A2(G401), .A3(new_n461), .A4(G227), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1188), .A2(new_n870), .ZN(new_n1189));
  NOR2_X1   g763(.A1(new_n917), .A2(new_n1189), .ZN(G308));
  AND2_X1   g764(.A1(new_n915), .A2(new_n912), .ZN(new_n1191));
  AND2_X1   g765(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n870), .B(new_n1188), .C1(new_n1191), .C2(new_n1192), .ZN(G225));
endmodule


