//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n465), .A2(new_n468), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n463), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n468), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n468), .A2(new_n463), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n463), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G124), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n468), .A2(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n463), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n488), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT71), .B1(new_n488), .B2(G2105), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n468), .A2(KEYINPUT4), .A3(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n463), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n492), .A2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G50), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n501), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT72), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n509), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n508), .A2(new_n516), .ZN(G166));
  OAI21_X1  g092(.A(G89), .B1(new_n505), .B2(new_n506), .ZN(new_n518));
  NAND2_X1  g093(.A1(G63), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(new_n512), .B1(G51), .B2(new_n500), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT73), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n524), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n523), .A2(KEYINPUT7), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT7), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(new_n500), .A2(G52), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OAI221_X1 g108(.A(new_n531), .B1(new_n532), .B2(new_n507), .C1(new_n533), .C2(new_n509), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  AOI22_X1  g110(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n509), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT6), .B(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n512), .A2(new_n538), .A3(G81), .ZN(new_n539));
  OAI211_X1 g114(.A(G43), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(KEYINPUT74), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT74), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n537), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n510), .B2(new_n511), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n504), .A2(new_n503), .ZN(new_n557));
  OAI211_X1 g132(.A(KEYINPUT76), .B(new_n554), .C1(new_n557), .C2(new_n552), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(G651), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT77), .A4(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n500), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n500), .A2(new_n567), .A3(G53), .ZN(new_n568));
  INV_X1    g143(.A(new_n507), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n569), .A2(KEYINPUT75), .A3(G91), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n507), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n566), .A2(new_n568), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n563), .A2(new_n574), .ZN(G299));
  NAND2_X1  g150(.A1(new_n500), .A2(G51), .ZN(new_n576));
  INV_X1    g151(.A(new_n519), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n538), .B2(G89), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n578), .B2(new_n557), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n523), .A2(new_n525), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n523), .A2(KEYINPUT7), .A3(new_n525), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n521), .A2(new_n586), .A3(new_n528), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G286));
  INV_X1    g164(.A(G166), .ZN(G303));
  NAND2_X1  g165(.A1(new_n569), .A2(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n500), .A2(G49), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  AOI22_X1  g169(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n509), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n500), .A2(G48), .ZN(new_n597));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n507), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n509), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n569), .A2(G85), .B1(G47), .B2(new_n500), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT79), .B(G66), .Z(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n557), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n500), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n507), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n512), .A2(new_n538), .A3(KEYINPUT10), .A4(G92), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n619), .A2(KEYINPUT80), .B1(G299), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(KEYINPUT80), .B2(new_n619), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(KEYINPUT80), .B2(new_n619), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n616), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n624), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  MUX2_X1   g203(.A(new_n544), .B(new_n628), .S(G868), .Z(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g205(.A1(new_n461), .A2(new_n462), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n470), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT82), .Z(new_n637));
  AOI22_X1  g212(.A1(new_n479), .A2(G123), .B1(new_n480), .B2(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n639), .A2(KEYINPUT83), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(KEYINPUT83), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n468), .B2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n638), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  OAI211_X1 g219(.A(new_n637), .B(new_n644), .C1(new_n635), .C2(new_n634), .ZN(G156));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  OAI21_X1  g224(.A(KEYINPUT14), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT85), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(KEYINPUT17), .ZN(new_n670));
  INV_X1    g245(.A(new_n664), .ZN(new_n671));
  INV_X1    g246(.A(new_n665), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n667), .A3(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(new_n666), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n669), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n680), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT87), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  OR2_X1    g271(.A1(G288), .A2(KEYINPUT89), .ZN(new_n697));
  NAND2_X1  g272(.A1(G288), .A2(KEYINPUT89), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  MUX2_X1   g274(.A(G23), .B(new_n699), .S(G16), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT33), .B(G1976), .Z(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G6), .A2(G16), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n600), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT32), .B(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n700), .B2(new_n701), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n708), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  INV_X1    g286(.A(G1971), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n702), .A2(new_n707), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n479), .A2(G119), .ZN(new_n720));
  OAI221_X1 g295(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n480), .A2(G131), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT88), .Z(new_n724));
  OAI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(new_n718), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n708), .A2(G24), .ZN(new_n730));
  INV_X1    g305(.A(G290), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n708), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1986), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n728), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n716), .A2(new_n717), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT36), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n479), .A2(G128), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT92), .Z(new_n738));
  OR2_X1    g313(.A1(new_n468), .A2(G116), .ZN(new_n739));
  INV_X1    g314(.A(G104), .ZN(new_n740));
  INV_X1    g315(.A(G2105), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT93), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT93), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n742), .A2(new_n743), .A3(new_n469), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n739), .A2(new_n744), .B1(new_n480), .B2(G140), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n738), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n718), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2067), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n708), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n708), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT98), .B(G1966), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n708), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n616), .B2(new_n708), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT91), .B(G1348), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n758), .B(new_n759), .Z(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT24), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n761), .B2(KEYINPUT24), .ZN(new_n763));
  AOI22_X1  g338(.A1(G160), .A2(G29), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G2084), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT31), .B(G11), .Z(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n718), .B1(new_n768), .B2(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT99), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n769), .A2(KEYINPUT99), .B1(new_n768), .B2(G28), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n643), .B2(new_n718), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n718), .A2(G32), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n479), .A2(G129), .B1(new_n480), .B2(G141), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT97), .B(KEYINPUT26), .Z(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n470), .A2(G105), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT27), .B(G1996), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n773), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  NOR2_X1   g359(.A1(G171), .A2(new_n708), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G5), .B2(new_n708), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n766), .B(new_n783), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n752), .A2(new_n756), .A3(new_n760), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G29), .A2(G35), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G162), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT29), .B(G2090), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n708), .A2(G19), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n545), .B2(new_n708), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1341), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n718), .A2(G27), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n718), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT101), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n788), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT25), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n480), .A2(G139), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n631), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n803), .B(new_n804), .C1(new_n468), .C2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G33), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT95), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2072), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n708), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  INV_X1    g386(.A(G299), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n708), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1956), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n786), .A2(new_n784), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n815), .B1(new_n781), .B2(new_n782), .C1(new_n764), .C2(G2084), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT100), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n809), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n736), .A2(new_n801), .A3(new_n818), .ZN(G311));
  INV_X1    g394(.A(G311), .ZN(G150));
  NAND2_X1  g395(.A1(new_n616), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT103), .ZN(new_n822));
  OAI211_X1 g397(.A(G55), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n507), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(G67), .B1(new_n504), .B2(new_n503), .ZN(new_n826));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n509), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(new_n537), .C1(new_n542), .C2(new_n543), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G81), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n540), .B1(new_n507), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(new_n541), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n829), .B1(new_n836), .B2(new_n537), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n822), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g417(.A(G860), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  INV_X1    g419(.A(new_n829), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(G145));
  XOR2_X1   g423(.A(new_n723), .B(KEYINPUT105), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n633), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n479), .A2(G130), .B1(new_n480), .B2(G142), .ZN(new_n851));
  OAI221_X1 g426(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n850), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT106), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(KEYINPUT106), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n746), .B(new_n780), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n806), .ZN(new_n859));
  XNOR2_X1  g434(.A(G164), .B(KEYINPUT104), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n856), .A2(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n854), .A2(KEYINPUT106), .ZN(new_n865));
  INV_X1    g440(.A(new_n863), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n861), .A4(new_n855), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G162), .B(G160), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n643), .ZN(new_n870));
  AOI21_X1  g445(.A(G37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n856), .A2(new_n857), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n862), .A2(new_n863), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n850), .B(new_n853), .Z(new_n875));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT107), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g456(.A(new_n838), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n628), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n616), .B1(new_n563), .B2(new_n574), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n563), .A2(new_n616), .A3(new_n574), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n885), .B2(new_n884), .ZN(new_n888));
  INV_X1    g463(.A(new_n616), .ZN(new_n889));
  NAND2_X1  g464(.A1(G299), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n563), .A2(new_n616), .A3(new_n574), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n886), .B1(new_n883), .B2(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n894), .A2(KEYINPUT42), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(KEYINPUT42), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G290), .B(G166), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n697), .A2(new_n698), .A3(G305), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G305), .B1(new_n697), .B2(new_n698), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n699), .A2(new_n600), .ZN(new_n903));
  XNOR2_X1  g478(.A(G303), .B(G290), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n897), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n895), .A2(new_n906), .A3(new_n896), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(G868), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n910), .A2(new_n911), .B1(new_n620), .B2(new_n845), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n908), .A2(KEYINPUT108), .A3(G868), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G295));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(G331));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n579), .A2(new_n584), .A3(KEYINPUT78), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n586), .B1(new_n521), .B2(new_n528), .ZN(new_n918));
  OAI21_X1  g493(.A(G171), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n544), .A2(new_n845), .ZN(new_n920));
  NAND2_X1  g495(.A1(G301), .A2(new_n529), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n830), .A4(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n533), .A2(new_n509), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n569), .A2(G90), .B1(G52), .B2(new_n500), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n926), .A2(new_n927), .B1(new_n521), .B2(new_n528), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n588), .B2(G171), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n838), .A2(new_n929), .A3(KEYINPUT109), .ZN(new_n930));
  AOI21_X1  g505(.A(G301), .B1(new_n585), .B2(new_n587), .ZN(new_n931));
  OAI22_X1  g506(.A1(new_n837), .A2(new_n831), .B1(new_n931), .B2(new_n928), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n924), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n893), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n885), .A2(new_n884), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n932), .A3(new_n922), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n906), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n924), .A2(new_n930), .A3(new_n935), .A4(new_n932), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n922), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n888), .A3(new_n892), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n940), .A3(new_n906), .ZN(new_n941));
  INV_X1    g516(.A(G37), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n916), .B1(new_n944), .B2(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n907), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(KEYINPUT110), .A3(new_n942), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n906), .B1(new_n938), .B2(new_n940), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n950), .B2(G37), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n941), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n946), .B2(new_n907), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n941), .B1(new_n955), .B2(KEYINPUT110), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n950), .A2(new_n949), .A3(G37), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT43), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n937), .A2(new_n943), .A3(KEYINPUT43), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n954), .B1(new_n961), .B2(new_n916), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n952), .B2(KEYINPUT43), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n963), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n953), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT112), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n953), .C1(new_n962), .C2(new_n964), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(G397));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n970));
  NAND3_X1  g545(.A1(G160), .A2(new_n970), .A3(G40), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n492), .B2(new_n495), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT115), .B1(new_n477), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1976), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n977), .B(G8), .C1(new_n978), .C2(new_n699), .ZN(new_n979));
  INV_X1    g554(.A(G288), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G1976), .ZN(new_n981));
  OR3_X1    g556(.A1(new_n979), .A2(KEYINPUT52), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(KEYINPUT52), .ZN(new_n983));
  INV_X1    g558(.A(new_n977), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1981), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n600), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT119), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(G1981), .B2(G305), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n986), .B1(new_n990), .B2(KEYINPUT49), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n992));
  AOI211_X1 g567(.A(new_n992), .B(new_n989), .C1(G1981), .C2(G305), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n982), .B(new_n983), .C1(new_n991), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(new_n971), .A3(new_n976), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n997));
  OR3_X1    g572(.A1(new_n996), .A2(G2090), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G164), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT113), .B(G1384), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n973), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1002), .A2(new_n1004), .A3(new_n976), .A4(new_n971), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT118), .B(G1971), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n985), .B1(new_n998), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G303), .A2(G8), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT55), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n994), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  OR4_X1    g589(.A1(new_n1014), .A2(new_n996), .A3(G2084), .A4(new_n997), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n971), .A2(new_n976), .ZN(new_n1016));
  INV_X1    g591(.A(new_n997), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n995), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1018), .B2(G2084), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1003), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n974), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1016), .B(new_n1021), .C1(KEYINPUT45), .C2(new_n974), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1015), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(G8), .A3(new_n588), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT63), .B1(new_n1013), .B2(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n997), .A2(KEYINPUT120), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1016), .A2(new_n1029), .A3(new_n995), .A4(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1007), .B1(new_n1032), .B2(G2090), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1011), .B1(new_n1033), .B2(G8), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n994), .A2(new_n1028), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1026), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n989), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n991), .A2(new_n993), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n980), .A2(new_n978), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n994), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n986), .A2(new_n1042), .B1(new_n1043), .B2(new_n1028), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1027), .A2(new_n1038), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT62), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1015), .A2(new_n1019), .A3(new_n1024), .A4(G168), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(G8), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1025), .A2(G8), .A3(new_n529), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1047), .B2(G8), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1046), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1047), .A2(G8), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT51), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1055), .A2(KEYINPUT62), .A3(new_n1050), .A4(new_n1049), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1005), .A2(G2078), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1058), .A2(new_n1059), .B1(new_n784), .B2(new_n1018), .ZN(new_n1060));
  OR3_X1    g635(.A1(new_n1022), .A2(new_n1059), .A3(G2078), .ZN(new_n1061));
  AOI21_X1  g636(.A(G301), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(new_n1035), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT122), .B(G1956), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1032), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n971), .A2(new_n976), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n973), .B2(new_n1003), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1002), .A3(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(G299), .B(KEYINPUT57), .Z(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G2067), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n984), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n759), .B1(new_n996), .B2(new_n997), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1074), .A2(new_n1075), .A3(KEYINPUT123), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT123), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1077));
  OR3_X1    g652(.A1(new_n1076), .A2(new_n1077), .A3(new_n889), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1070), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1072), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(KEYINPUT61), .A3(new_n1071), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1076), .A2(new_n1077), .A3(KEYINPUT60), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT60), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n889), .A2(KEYINPUT126), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n889), .A2(KEYINPUT126), .ZN(new_n1090));
  OR3_X1    g665(.A1(new_n1087), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1996), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1067), .A2(KEYINPUT124), .A3(new_n1093), .A4(new_n1002), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1005), .B2(G1996), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT58), .B(G1341), .Z(new_n1098));
  NAND2_X1  g673(.A1(new_n977), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT125), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1099), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1101), .B(new_n1102), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n545), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT59), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n545), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1081), .B1(new_n1092), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1020), .B1(new_n999), .B2(new_n1001), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n477), .A2(new_n975), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1059), .A2(G2078), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1002), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1060), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(G171), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1110), .B1(new_n1117), .B2(new_n1062), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1055), .A2(new_n1050), .A3(new_n1049), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(G171), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1060), .A2(G301), .A3(new_n1061), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(KEYINPUT54), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1118), .A2(new_n1119), .A3(new_n1035), .A4(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1045), .B(new_n1063), .C1(new_n1109), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1016), .A2(new_n1111), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n746), .B(new_n1073), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n780), .A2(G1996), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1125), .A2(G1996), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT117), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n780), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1125), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n723), .B(new_n727), .Z(new_n1134));
  AOI211_X1 g709(.A(new_n1128), .B(new_n1132), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G290), .A2(G1986), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT116), .ZN(new_n1137));
  AND2_X1   g712(.A1(G290), .A2(G1986), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1133), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1124), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1126), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1133), .B1(new_n1142), .B2(new_n780), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1131), .A2(KEYINPUT46), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT46), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1130), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT47), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT48), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1135), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n724), .A2(new_n727), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1132), .A2(new_n1128), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n746), .A2(G2067), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1133), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1148), .A2(new_n1151), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1141), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g732(.A(G319), .ZN(new_n1159));
  NOR2_X1   g733(.A1(G227), .A2(new_n1159), .ZN(new_n1160));
  XOR2_X1   g734(.A(new_n1160), .B(KEYINPUT127), .Z(new_n1161));
  NOR3_X1   g735(.A1(new_n662), .A2(G229), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g736(.A1(new_n880), .A2(new_n1162), .A3(new_n961), .ZN(G225));
  INV_X1    g737(.A(G225), .ZN(G308));
endmodule


