//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(G2106), .B2(new_n453), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n464), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(KEYINPUT3), .A3(new_n471), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n474), .A2(G137), .A3(new_n475), .A4(new_n463), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  AND3_X1   g053(.A1(new_n474), .A2(new_n475), .A3(new_n463), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n474), .A2(G2105), .A3(new_n463), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  MUX2_X1   g057(.A(G100), .B(G112), .S(G2105), .Z(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2104), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND2_X1  g061(.A1(new_n463), .A2(new_n465), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(new_n475), .A3(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n474), .A2(G138), .A3(new_n475), .A4(new_n463), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n474), .A2(G126), .A3(G2105), .A4(new_n463), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G102), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n494), .B1(new_n497), .B2(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n475), .A2(G102), .ZN(new_n499));
  AOI211_X1 g074(.A(KEYINPUT69), .B(new_n464), .C1(new_n499), .C2(new_n495), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n493), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n492), .A2(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(G50), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT70), .A3(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(new_n516), .B1(KEYINPUT6), .B2(new_n505), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT71), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n512), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n506), .B1(new_n519), .B2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT72), .Z(new_n524));
  XOR2_X1   g099(.A(KEYINPUT74), .B(G89), .Z(new_n525));
  NAND3_X1  g100(.A1(new_n517), .A2(new_n503), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n514), .A2(new_n516), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  OAI211_X1 g111(.A(G51), .B(G543), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n526), .A2(KEYINPUT75), .A3(new_n528), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n524), .A2(new_n531), .A3(new_n537), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n510), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n505), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(new_n544), .B2(new_n543), .ZN(new_n546));
  OAI211_X1 g121(.A(G52), .B(G543), .C1(new_n535), .C2(new_n536), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n532), .A2(new_n534), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n510), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G90), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n548), .B1(new_n547), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n546), .B1(new_n552), .B2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n510), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n550), .A2(G81), .B1(G651), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g134(.A(G43), .B(G543), .C1(new_n535), .C2(new_n536), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT78), .Z(G188));
  OAI21_X1  g143(.A(G543), .B1(new_n535), .B2(new_n536), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n549), .A2(KEYINPUT73), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n517), .A2(new_n533), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(new_n576), .A3(G53), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g153(.A(KEYINPUT79), .B(G65), .Z(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(new_n503), .B1(G78), .B2(G543), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n505), .B1(new_n580), .B2(new_n581), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n582), .A2(new_n583), .B1(G91), .B2(new_n550), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n578), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(new_n521), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n520), .B1(new_n512), .B2(new_n517), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n586), .A2(new_n587), .B1(new_n505), .B2(new_n504), .ZN(G303));
  NAND2_X1  g163(.A1(new_n575), .A2(G49), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n503), .A2(G74), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n550), .A2(G87), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G288));
  OAI211_X1 g167(.A(KEYINPUT81), .B(G61), .C1(new_n508), .C2(new_n509), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(KEYINPUT81), .B1(new_n503), .B2(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n503), .A2(G86), .ZN(new_n598));
  AND2_X1   g173(.A1(G48), .A2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n517), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n575), .A2(G47), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n510), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n550), .A2(G85), .B1(G651), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(G290));
  NAND3_X1  g182(.A1(new_n517), .A2(G92), .A3(new_n503), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .A4(new_n503), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g187(.A(G54), .B(G543), .C1(new_n535), .C2(new_n536), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n503), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(new_n505), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g193(.A(new_n617), .B1(G171), .B2(G868), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NOR2_X1   g195(.A1(G286), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G299), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n620), .ZN(G297));
  XNOR2_X1  g198(.A(G297), .B(KEYINPUT82), .ZN(G280));
  AND3_X1   g199(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  NOR2_X1   g202(.A1(new_n561), .A2(G868), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n616), .A2(G559), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g206(.A1(new_n472), .A2(new_n463), .A3(new_n465), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT13), .B(G2100), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n479), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n481), .A2(G123), .ZN(new_n638));
  AND2_X1   g213(.A1(G111), .A2(G2105), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(G99), .B2(new_n475), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n637), .B(new_n638), .C1(new_n464), .C2(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n642), .A3(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2427), .ZN(new_n648));
  INV_X1    g223(.A(G2430), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(KEYINPUT17), .ZN(new_n666));
  INV_X1    g241(.A(new_n662), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(new_n661), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n661), .B1(new_n666), .B2(new_n662), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(KEYINPUT84), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(new_n667), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT85), .B1(new_n669), .B2(new_n671), .ZN(new_n675));
  OAI221_X1 g250(.A(new_n665), .B1(new_n666), .B2(new_n668), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2096), .ZN(new_n677));
  INV_X1    g252(.A(G2100), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(G2096), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n676), .A2(G2096), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(G2100), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n688), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(new_n694), .B(new_n693), .S(new_n686), .Z(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  XOR2_X1   g275(.A(G1981), .B(G1986), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n698), .B(new_n702), .ZN(G229));
  NAND2_X1  g278(.A1(new_n562), .A2(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G16), .B2(G19), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G1341), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n705), .B(KEYINPUT91), .ZN(new_n709));
  INV_X1    g284(.A(G1341), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  NOR2_X1   g287(.A1(G5), .A2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT95), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(G301), .B2(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n708), .A2(new_n711), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G4), .A2(G16), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n625), .B2(G16), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT90), .B(G1348), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G32), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n479), .A2(G141), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n481), .A2(G129), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT26), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  AOI22_X1  g304(.A1(G105), .A2(new_n472), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n724), .A2(new_n725), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n723), .B1(new_n732), .B2(new_n722), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT27), .B(G1996), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  NOR2_X1   g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n722), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n477), .B2(new_n722), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT31), .B(G11), .Z(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n722), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n641), .B2(new_n722), .ZN(new_n746));
  NOR4_X1   g321(.A1(new_n735), .A2(new_n741), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n722), .A2(G33), .ZN(new_n748));
  NAND2_X1  g323(.A1(G115), .A2(G2104), .ZN(new_n749));
  INV_X1    g324(.A(G127), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n487), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G2105), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT25), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n479), .B2(G139), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n748), .B1(new_n757), .B2(new_n722), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G2072), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n722), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  NAND2_X1  g336(.A1(G116), .A2(G2105), .ZN(new_n762));
  INV_X1    g337(.A(G104), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G2105), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G2104), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT92), .ZN(new_n766));
  INV_X1    g341(.A(G128), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n474), .A2(G2105), .A3(new_n463), .ZN(new_n768));
  INV_X1    g343(.A(G140), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n474), .A2(new_n475), .A3(new_n463), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n766), .B1(new_n767), .B2(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n761), .B1(new_n772), .B2(new_n722), .ZN(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AND4_X1   g350(.A1(new_n721), .A2(new_n747), .A3(new_n759), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G29), .A2(G35), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G162), .B2(G29), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT29), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2090), .ZN(new_n780));
  NOR2_X1   g355(.A1(G27), .A2(G29), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G164), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT96), .B(G2078), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G168), .A2(new_n715), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n715), .B2(G21), .ZN(new_n786));
  INV_X1    g361(.A(G1966), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n717), .A2(new_n776), .A3(new_n780), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n715), .A2(G20), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT23), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n622), .B2(new_n715), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1956), .Z(new_n795));
  OAI211_X1 g370(.A(new_n791), .B(new_n795), .C1(new_n712), .C2(new_n716), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n789), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G290), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G16), .ZN(new_n799));
  OR2_X1    g374(.A1(G16), .A2(G24), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  OAI21_X1  g380(.A(G1986), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n799), .A2(new_n800), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT88), .ZN(new_n808));
  INV_X1    g383(.A(G1986), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n808), .A2(new_n809), .A3(new_n803), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n715), .A2(G23), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n589), .A2(new_n591), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n715), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT33), .B(G1976), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT89), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  MUX2_X1   g392(.A(G6), .B(G305), .S(G16), .Z(new_n818));
  XOR2_X1   g393(.A(KEYINPUT32), .B(G1981), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(G16), .A2(G22), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G166), .B2(G16), .ZN(new_n822));
  INV_X1    g397(.A(G1971), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n817), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT34), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n817), .A2(new_n827), .A3(new_n820), .A4(new_n824), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n479), .A2(G131), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n481), .A2(G119), .ZN(new_n830));
  AND2_X1   g405(.A1(G107), .A2(G2105), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G95), .B2(new_n475), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n464), .C2(new_n832), .ZN(new_n833));
  MUX2_X1   g408(.A(G25), .B(new_n833), .S(G29), .Z(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT35), .B(G1991), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT87), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n834), .B(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n811), .A2(new_n826), .A3(new_n828), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n828), .A2(new_n838), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n841), .A2(new_n842), .A3(new_n826), .A4(new_n811), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n797), .A2(new_n844), .ZN(G311));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n797), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n846), .B1(new_n797), .B2(new_n844), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(G150));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n510), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G651), .ZN(new_n853));
  OAI211_X1 g428(.A(G55), .B(G543), .C1(new_n535), .C2(new_n536), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT98), .B(G93), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n550), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(KEYINPUT99), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT99), .B1(new_n854), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NOR2_X1   g437(.A1(new_n616), .A2(new_n626), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT38), .Z(new_n864));
  NAND3_X1  g439(.A1(new_n559), .A2(KEYINPUT100), .A3(new_n560), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n866), .B(new_n853), .C1(new_n858), .C2(new_n859), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n854), .A2(new_n856), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n870), .A2(new_n857), .B1(G651), .B2(new_n852), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n561), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n865), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n867), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n864), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(G860), .B1(new_n876), .B2(new_n877), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n878), .A2(KEYINPUT101), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT101), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n862), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT102), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n884), .B(new_n862), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G145));
  XNOR2_X1  g461(.A(G160), .B(new_n485), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(new_n641), .Z(new_n888));
  MUX2_X1   g463(.A(G106), .B(G118), .S(G2105), .Z(new_n889));
  AOI22_X1  g464(.A1(new_n481), .A2(G130), .B1(G2104), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n479), .A2(G142), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n833), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n634), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n501), .B1(new_n492), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n897));
  INV_X1    g472(.A(new_n490), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT103), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n731), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n894), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n771), .B(KEYINPUT104), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n757), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n894), .A2(new_n902), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n905), .B1(new_n903), .B2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n888), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n894), .B(new_n902), .ZN(new_n912));
  INV_X1    g487(.A(new_n905), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n888), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n907), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n910), .A2(new_n911), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g493(.A(new_n875), .B(new_n629), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n578), .A2(new_n625), .A3(new_n584), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n625), .B1(new_n578), .B2(new_n584), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(G299), .A2(new_n616), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n578), .A2(new_n625), .A3(new_n584), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(KEYINPUT105), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n924), .A2(new_n929), .A3(new_n925), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT41), .B1(new_n921), .B2(new_n922), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n919), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n934));
  NAND2_X1  g509(.A1(G288), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(G288), .A2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n798), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n813), .A2(KEYINPUT106), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(G290), .A3(new_n935), .ZN(new_n940));
  XNOR2_X1  g515(.A(G166), .B(G305), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n942), .B1(new_n938), .B2(new_n940), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n940), .ZN(new_n952));
  AOI21_X1  g527(.A(G290), .B1(new_n939), .B2(new_n935), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n941), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n954), .B2(new_n943), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n933), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n928), .A2(new_n948), .A3(new_n956), .A4(new_n932), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G868), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n871), .A2(new_n620), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(KEYINPUT108), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n620), .B1(new_n958), .B2(new_n959), .ZN(new_n965));
  INV_X1    g540(.A(new_n962), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n963), .A2(new_n967), .ZN(G295));
  NAND3_X1  g543(.A1(new_n961), .A2(KEYINPUT109), .A3(new_n962), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n965), .B2(new_n966), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(G331));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  OAI211_X1 g548(.A(G168), .B(new_n546), .C1(new_n553), .C2(new_n552), .ZN(new_n974));
  NAND2_X1  g549(.A1(G301), .A2(G286), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n875), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n860), .A2(new_n873), .A3(new_n865), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(new_n867), .A3(new_n974), .A4(new_n975), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n927), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n931), .A2(new_n930), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n921), .A2(new_n922), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(KEYINPUT110), .A3(new_n929), .ZN(new_n986));
  INV_X1    g561(.A(new_n979), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n978), .A2(new_n867), .B1(new_n974), .B2(new_n975), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n984), .B(new_n986), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n927), .A2(new_n977), .A3(KEYINPUT111), .A4(new_n979), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n982), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n946), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n977), .A2(new_n985), .A3(new_n979), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n977), .A2(new_n979), .B1(new_n930), .B2(new_n931), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n954), .A2(new_n943), .ZN(new_n996));
  AOI21_X1  g571(.A(G37), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n973), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n994), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n977), .A2(new_n979), .A3(new_n985), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n996), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n946), .B1(new_n993), .B2(new_n994), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n973), .A2(new_n1001), .A3(new_n911), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT44), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n992), .B2(new_n997), .ZN(new_n1006));
  AND4_X1   g581(.A1(KEYINPUT43), .A2(new_n1001), .A3(new_n911), .A4(new_n1002), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1004), .A2(new_n1008), .ZN(G397));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n897), .A2(new_n895), .A3(new_n898), .ZN(new_n1011));
  INV_X1    g586(.A(new_n501), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n492), .A2(new_n895), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n468), .A2(G2105), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n472), .A2(G101), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1016), .A2(G40), .A3(new_n476), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n473), .A2(new_n1020), .A3(G40), .A4(new_n476), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n1024));
  NAND3_X1  g599(.A1(new_n1015), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT115), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1015), .A2(new_n1023), .A3(new_n1027), .A4(new_n1024), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n771), .B(G2067), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(KEYINPUT116), .A3(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1026), .A2(G1996), .A3(new_n731), .A4(new_n1028), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1025), .A2(G1996), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n732), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G290), .A2(G1986), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT114), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G290), .A2(G1986), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1025), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n833), .B(new_n837), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1029), .A2(new_n1045), .ZN(new_n1046));
  NOR4_X1   g621(.A1(new_n1036), .A2(new_n1040), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT45), .B1(new_n901), .B2(new_n1010), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1010), .B1(new_n492), .B2(new_n501), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1019), .B(new_n1021), .C1(new_n1049), .C2(new_n1024), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n787), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(new_n1010), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1049), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT117), .B1(new_n1049), .B2(KEYINPUT50), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1053), .B(new_n1023), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1051), .B(G168), .C1(G2084), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT51), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1051), .B1(G2084), .B2(new_n1056), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(G286), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1059), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(G166), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT50), .B(new_n1010), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1022), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT118), .B(G2090), .Z(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT45), .B(new_n1010), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1049), .A2(new_n1024), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1023), .A3(new_n1075), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1072), .A2(new_n1073), .B1(new_n1076), .B2(new_n823), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1069), .B1(new_n1077), .B2(new_n1065), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT119), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1073), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1056), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1075), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1971), .B1(new_n1086), .B2(new_n1074), .ZN(new_n1087));
  OAI211_X1 g662(.A(G8), .B(new_n1082), .C1(new_n1084), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n589), .A2(G1976), .A3(new_n591), .ZN(new_n1090));
  OAI211_X1 g665(.A(G8), .B(new_n1090), .C1(new_n1015), .C2(new_n1022), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n813), .B2(G1976), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1089), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1384), .B1(new_n896), .B2(new_n900), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1065), .B1(new_n1023), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1976), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(G288), .B2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1096), .A2(KEYINPUT120), .A3(new_n1090), .A4(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n597), .A2(new_n600), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n597), .B2(new_n600), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT121), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(new_n1104), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1105), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1110), .A2(new_n1096), .B1(KEYINPUT52), .B2(new_n1091), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1078), .A2(new_n1088), .A3(new_n1100), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT125), .B(KEYINPUT53), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1076), .B2(G2078), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1056), .A2(new_n712), .ZN(new_n1117));
  INV_X1    g692(.A(G2078), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT53), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1018), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1024), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1074), .B(new_n1120), .C1(new_n1095), .C2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1116), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1114), .B1(new_n1123), .B2(G171), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT45), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1050), .B1(new_n1015), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1119), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1056), .A2(new_n712), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1116), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1124), .B1(G171), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1123), .A2(G171), .ZN(new_n1131));
  AOI21_X1  g706(.A(G301), .B1(new_n1128), .B2(new_n1116), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1114), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1063), .A2(new_n1113), .A3(new_n1130), .A4(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT56), .B(G2072), .Z(new_n1135));
  OAI22_X1  g710(.A1(new_n1072), .A2(G1956), .B1(new_n1076), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G299), .B(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1138), .A2(KEYINPUT123), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(KEYINPUT123), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1076), .A2(new_n1135), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1138), .B(new_n1142), .C1(G1956), .C2(new_n1072), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  INV_X1    g720(.A(G1348), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1056), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1023), .A2(new_n1095), .A3(new_n774), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n625), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n616), .A3(new_n1148), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1145), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n1153));
  INV_X1    g728(.A(G1996), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1074), .A2(new_n1023), .A3(new_n1154), .A4(new_n1075), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT58), .B(G1341), .Z(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n1158), .B2(new_n562), .ZN(new_n1159));
  AOI211_X1 g734(.A(KEYINPUT59), .B(new_n561), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n625), .A2(new_n1145), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1159), .A2(new_n1160), .B1(new_n1149), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1152), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  XNOR2_X1  g739(.A(G299), .B(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1136), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1143), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g744(.A(KEYINPUT124), .B(KEYINPUT61), .C1(new_n1143), .C2(new_n1166), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1144), .B(new_n1163), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1143), .A2(new_n625), .A3(new_n1149), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1141), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1134), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n1175));
  NOR2_X1   g750(.A1(G286), .A2(new_n1065), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1049), .A2(KEYINPUT50), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT117), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1049), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1182), .A2(new_n740), .A3(new_n1023), .A4(new_n1053), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1177), .B1(new_n1183), .B2(new_n1051), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1175), .B1(new_n1112), .B2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1182), .A2(new_n1023), .A3(new_n1053), .A4(new_n1073), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1125), .B(G1384), .C1(new_n896), .C2(new_n900), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n823), .B1(new_n1188), .B2(new_n1085), .ZN(new_n1189));
  AOI221_X4 g764(.A(new_n1065), .B1(new_n1080), .B2(new_n1081), .C1(new_n1187), .C2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1189), .B1(new_n1056), .B2(new_n1083), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1068), .B1(new_n1191), .B2(G8), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1100), .A2(new_n1111), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1061), .A2(KEYINPUT63), .A3(new_n1176), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1193), .A2(new_n1196), .A3(KEYINPUT122), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1065), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1088), .B1(new_n1068), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1184), .A2(new_n1100), .A3(new_n1111), .A4(KEYINPUT63), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1186), .A2(new_n1197), .A3(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1062), .A2(new_n1058), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1060), .B1(new_n1057), .B2(G8), .ZN(new_n1205));
  OAI21_X1  g780(.A(KEYINPUT62), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1132), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1112), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1059), .B(new_n1209), .C1(new_n1058), .C2(new_n1062), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1194), .A2(new_n1088), .ZN(new_n1212));
  AOI211_X1 g787(.A(G1976), .B(G288), .C1(new_n1110), .C2(new_n1096), .ZN(new_n1213));
  OR2_X1    g788(.A1(new_n1213), .A2(new_n1102), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1212), .B1(new_n1096), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1203), .A2(new_n1211), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1047), .B1(new_n1174), .B2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1038), .B(KEYINPUT46), .ZN(new_n1218));
  OAI211_X1 g793(.A(new_n1026), .B(new_n1028), .C1(new_n731), .C2(new_n1031), .ZN(new_n1219));
  OR2_X1    g794(.A1(new_n1219), .A2(KEYINPUT126), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(KEYINPUT126), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1218), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT47), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n1042), .A2(new_n1025), .ZN(new_n1224));
  XNOR2_X1  g799(.A(new_n1224), .B(KEYINPUT48), .ZN(new_n1225));
  NOR4_X1   g800(.A1(new_n1036), .A2(new_n1225), .A3(new_n1046), .A4(new_n1040), .ZN(new_n1226));
  NOR2_X1   g801(.A1(new_n833), .A2(new_n836), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1040), .ZN(new_n1228));
  NAND4_X1  g803(.A1(new_n1034), .A2(new_n1227), .A3(new_n1228), .A4(new_n1035), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n772), .A2(new_n774), .ZN(new_n1230));
  AOI21_X1  g805(.A(new_n1029), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g806(.A1(new_n1223), .A2(new_n1226), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1217), .A2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g808(.A1(G229), .A2(G401), .ZN(new_n1235));
  NAND3_X1  g809(.A1(new_n679), .A2(G319), .A3(new_n682), .ZN(new_n1236));
  OAI21_X1  g810(.A(new_n1235), .B1(new_n1236), .B2(KEYINPUT127), .ZN(new_n1237));
  AND2_X1   g811(.A1(new_n1236), .A2(KEYINPUT127), .ZN(new_n1238));
  NOR2_X1   g812(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n917), .A2(new_n1239), .ZN(new_n1240));
  NOR3_X1   g814(.A1(new_n1240), .A2(new_n1006), .A3(new_n1007), .ZN(G308));
  OR3_X1    g815(.A1(new_n1240), .A2(new_n1006), .A3(new_n1007), .ZN(G225));
endmodule


