//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n205), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n205), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n216), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n215), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT9), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT72), .ZN(new_n246));
  NOR3_X1   g0046(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n220), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  OAI22_X1  g0050(.A1(new_n247), .A2(new_n220), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT8), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G58), .ZN(new_n254));
  INV_X1    g0054(.A(G58), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(KEYINPUT8), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(KEYINPUT8), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(G58), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT66), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n220), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(new_n220), .A3(G33), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n251), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n219), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT68), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n275), .A2(new_n272), .A3(G13), .A4(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n220), .A2(G1), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n207), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n270), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(G50), .B2(new_n277), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n246), .B1(new_n271), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n267), .A2(new_n270), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(KEYINPUT72), .A3(new_n281), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n245), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G222), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(G223), .A3(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n289), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  AND2_X1   g0102(.A1(G1), .A2(G13), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n295), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  INV_X1    g0105(.A(G45), .ZN(new_n306));
  AOI21_X1  g0106(.A(G1), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n301), .A2(G226), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n298), .A2(G190), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n271), .A2(new_n246), .A3(new_n282), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT72), .B1(new_n284), .B2(new_n281), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(KEYINPUT9), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n286), .A2(KEYINPUT73), .A3(new_n309), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n298), .A2(new_n308), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G200), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n286), .A2(new_n317), .A3(new_n309), .A4(new_n312), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n313), .A3(new_n314), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT74), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n271), .A2(new_n282), .B1(new_n324), .B2(new_n316), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G179), .B2(new_n316), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n210), .A2(G1698), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(G232), .B2(G1698), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n328), .A2(new_n289), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n297), .B1(new_n289), .B2(G107), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n307), .A2(new_n296), .A3(G274), .ZN(new_n332));
  INV_X1    g0132(.A(G244), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n300), .ZN(new_n334));
  OR3_X1    g0134(.A1(new_n331), .A2(KEYINPUT69), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT69), .B1(new_n331), .B2(new_n334), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(new_n324), .A3(new_n336), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n277), .A2(new_n270), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n278), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(G77), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n274), .A2(new_n276), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n293), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G20), .A2(G33), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n349), .A2(KEYINPUT70), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(KEYINPUT70), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n354), .A2(new_n262), .B1(new_n220), .B2(new_n293), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n346), .B(new_n348), .C1(new_n270), .C2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n342), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n337), .A2(KEYINPUT71), .A3(new_n338), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n341), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n357), .B1(new_n337), .B2(G190), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(new_n337), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n322), .A2(new_n323), .A3(new_n326), .A4(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n320), .A2(new_n321), .A3(new_n326), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT74), .B1(new_n367), .B2(new_n364), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n263), .A2(G77), .A3(new_n265), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n349), .A2(G50), .B1(G20), .B2(new_n209), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n270), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(KEYINPUT11), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n343), .A2(new_n209), .A3(new_n278), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OR3_X1    g0174(.A1(new_n277), .A2(KEYINPUT12), .A3(G68), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT12), .B1(new_n277), .B2(G68), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n375), .A2(new_n376), .B1(KEYINPUT11), .B2(new_n371), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT77), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT77), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n229), .A2(G1698), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(G226), .B2(G1698), .ZN(new_n385));
  AND2_X1   g0185(.A1(KEYINPUT3), .A2(G33), .ZN(new_n386));
  NOR2_X1   g0186(.A1(KEYINPUT3), .A2(G33), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n383), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n297), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n296), .A2(G238), .A3(new_n299), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n332), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(new_n332), .B2(new_n391), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT13), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(new_n390), .C1(new_n393), .C2(new_n394), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n396), .A2(G179), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(KEYINPUT76), .A3(new_n398), .ZN(new_n400));
  OR3_X1    g0200(.A1(new_n395), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(G169), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(KEYINPUT78), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n399), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n404), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n400), .A2(new_n401), .A3(G169), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n382), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G190), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n395), .B2(KEYINPUT13), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n379), .A2(new_n381), .B1(new_n398), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n400), .A2(new_n401), .A3(G200), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n287), .A2(new_n220), .A3(new_n288), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n388), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n209), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n255), .A2(new_n209), .ZN(new_n421));
  NOR2_X1   g0221(.A1(G58), .A2(G68), .ZN(new_n422));
  OAI21_X1  g0222(.A(G20), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n349), .A2(G159), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n415), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT7), .B1(new_n388), .B2(new_n220), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n386), .A2(new_n387), .A3(new_n417), .A4(G20), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n425), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT16), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n431), .A3(new_n269), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n261), .A2(new_n277), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n257), .A2(new_n260), .A3(new_n345), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n343), .B1(KEYINPUT79), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n257), .A2(new_n436), .A3(new_n260), .A4(new_n345), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n433), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(G223), .A2(G1698), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n208), .A2(G1698), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n441), .C1(new_n386), .C2(new_n387), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G87), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n297), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n296), .A2(G232), .A3(new_n299), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n332), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n447), .A3(new_n338), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n296), .B1(new_n442), .B2(new_n443), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n332), .A2(new_n446), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n324), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n439), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT18), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n362), .B1(new_n445), .B2(new_n447), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT80), .B(G190), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n449), .A2(new_n450), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n432), .A2(new_n438), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT17), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n452), .B1(new_n432), .B2(new_n438), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT18), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n432), .A2(new_n438), .A3(new_n459), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT17), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n455), .A2(new_n461), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n408), .A2(new_n414), .A3(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n366), .A2(new_n368), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT4), .A2(G244), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n290), .B(new_n472), .C1(new_n386), .C2(new_n387), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n333), .B1(new_n287), .B2(new_n288), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(KEYINPUT4), .ZN(new_n476));
  OAI21_X1  g0276(.A(G250), .B1(new_n386), .B2(new_n387), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n290), .B1(new_n477), .B2(KEYINPUT4), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n297), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n306), .A2(G1), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(G33), .A2(G41), .ZN(new_n484));
  OAI21_X1  g0284(.A(G274), .B1(new_n484), .B2(new_n219), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT81), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n304), .A2(new_n487), .A3(new_n488), .A4(new_n480), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n488), .A2(new_n480), .B1(new_n303), .B2(new_n295), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n486), .A2(new_n489), .B1(new_n490), .B2(G257), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n479), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G200), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n272), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n277), .A2(G97), .A3(new_n270), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G97), .B2(new_n277), .ZN(new_n496));
  OAI21_X1  g0296(.A(G107), .B1(new_n427), .B2(new_n428), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  AND2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n202), .ZN(new_n500));
  INV_X1    g0300(.A(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n349), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n496), .B1(new_n269), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n479), .A2(new_n491), .A3(G190), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n493), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(G20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n349), .A2(G77), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n501), .B1(new_n418), .B2(new_n419), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n269), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n277), .A2(G97), .ZN(new_n514));
  INV_X1    g0314(.A(new_n494), .ZN(new_n515));
  AOI211_X1 g0315(.A(new_n269), .B(new_n515), .C1(new_n274), .C2(new_n276), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n479), .A2(new_n491), .A3(G179), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n324), .B1(new_n479), .B2(new_n491), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n471), .B1(new_n508), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n507), .A2(new_n513), .A3(new_n517), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT82), .B1(new_n523), .B2(new_n493), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n475), .A2(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n289), .A2(G238), .A3(new_n290), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n297), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n272), .A2(G45), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G250), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n297), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n296), .A2(KEYINPUT83), .A3(G250), .A4(new_n531), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(new_n304), .B2(new_n480), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n289), .A2(new_n220), .A3(G68), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n220), .B1(new_n383), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(G87), .B2(new_n203), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n220), .A2(G33), .A3(G97), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n543), .A2(KEYINPUT84), .A3(new_n539), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT84), .B1(new_n543), .B2(new_n539), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n269), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n347), .A2(new_n354), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n529), .A2(G190), .A3(new_n535), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n516), .A2(G87), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n537), .A2(new_n549), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n536), .A2(new_n324), .ZN(new_n553));
  INV_X1    g0353(.A(new_n354), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n516), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n547), .A2(new_n548), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n529), .A2(new_n338), .A3(new_n535), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n522), .A2(new_n524), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n220), .B(G87), .C1(new_n386), .C2(new_n387), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n289), .A2(new_n563), .A3(new_n220), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OR3_X1    g0365(.A1(new_n220), .A2(KEYINPUT23), .A3(G107), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT86), .B1(new_n527), .B2(G20), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT23), .B1(new_n220), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n527), .A2(KEYINPUT86), .A3(G20), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n565), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n565), .B2(new_n571), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n269), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n347), .A2(KEYINPUT25), .A3(new_n501), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT25), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n277), .B2(G107), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n576), .A2(new_n578), .B1(new_n516), .B2(G107), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(G1698), .C1(new_n386), .C2(new_n387), .ZN(new_n581));
  OAI211_X1 g0381(.A(G250), .B(new_n290), .C1(new_n386), .C2(new_n387), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G294), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n296), .B1(new_n584), .B2(KEYINPUT87), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT87), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n581), .A2(new_n582), .A3(new_n586), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n486), .A2(new_n489), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n490), .A2(G264), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n324), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n585), .A2(new_n587), .B1(G264), .B2(new_n490), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n338), .A3(new_n589), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n580), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(G264), .B(G1698), .C1(new_n386), .C2(new_n387), .ZN(new_n596));
  OAI211_X1 g0396(.A(G257), .B(new_n290), .C1(new_n386), .C2(new_n387), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n287), .A2(G303), .A3(new_n288), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n297), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n490), .A2(G270), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n589), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  INV_X1    g0403(.A(G116), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n347), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n277), .A2(G116), .A3(new_n270), .A4(new_n494), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n268), .A2(new_n219), .B1(G20), .B2(new_n604), .ZN(new_n607));
  INV_X1    g0407(.A(G97), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n474), .B(new_n220), .C1(G33), .C2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT20), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n607), .A2(KEYINPUT20), .A3(new_n609), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n605), .B(new_n606), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n486), .A2(new_n489), .B1(new_n490), .B2(G270), .ZN(new_n614));
  INV_X1    g0414(.A(new_n457), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n600), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n603), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT85), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT85), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n603), .A2(new_n613), .A3(new_n619), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n602), .A2(new_n612), .A3(G169), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n612), .A2(G179), .A3(new_n600), .A4(new_n614), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n602), .A2(new_n612), .A3(KEYINPUT21), .A4(G169), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n591), .A2(G200), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n593), .A2(G190), .A3(new_n589), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n628), .A2(new_n575), .A3(new_n579), .A4(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n621), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n470), .A2(new_n560), .A3(new_n595), .A4(new_n631), .ZN(G372));
  OAI21_X1  g0432(.A(KEYINPUT89), .B1(new_n519), .B2(new_n520), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n492), .A2(G169), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT89), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n479), .A2(new_n491), .A3(G179), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n637), .A3(new_n518), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT90), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  INV_X1    g0440(.A(new_n559), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n633), .A2(new_n637), .A3(new_n642), .A4(new_n518), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n558), .A2(KEYINPUT88), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n553), .A2(new_n556), .A3(new_n646), .A4(new_n557), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n521), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n558), .A3(new_n552), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(KEYINPUT26), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT91), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT91), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n644), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n522), .A2(new_n524), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n627), .A2(new_n595), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(new_n641), .A3(new_n657), .A4(new_n630), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n653), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n470), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n326), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n463), .B1(new_n439), .B2(new_n453), .ZN(new_n663));
  AOI211_X1 g0463(.A(KEYINPUT18), .B(new_n452), .C1(new_n432), .C2(new_n438), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n455), .A2(KEYINPUT92), .A3(new_n464), .ZN(new_n666));
  INV_X1    g0466(.A(new_n360), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n408), .B1(new_n667), .B2(new_n413), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n465), .B(KEYINPUT17), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n665), .B(new_n666), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n661), .B1(new_n671), .B2(new_n322), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n660), .A2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n272), .A2(new_n220), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n612), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n621), .A2(new_n627), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n627), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n580), .A2(new_n592), .A3(new_n594), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n580), .A2(new_n679), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n630), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n595), .A2(new_n679), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n627), .A2(new_n679), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n223), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n218), .ZN(new_n697));
  INV_X1    g0497(.A(G87), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n202), .A2(new_n698), .A3(new_n604), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT93), .Z(new_n700));
  NOR3_X1   g0500(.A1(new_n700), .A2(new_n272), .A3(new_n696), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT94), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n702), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  XNOR2_X1  g0505(.A(KEYINPUT96), .B(KEYINPUT30), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n589), .A2(new_n600), .A3(G179), .A4(new_n601), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT95), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n529), .A2(new_n535), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n614), .A2(new_n710), .A3(G179), .A4(new_n600), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n593), .A4(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n706), .B1(new_n712), .B2(new_n492), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n709), .A2(new_n593), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n479), .A2(new_n491), .A3(KEYINPUT30), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n708), .A3(new_n711), .A4(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n591), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n536), .A2(new_n492), .A3(new_n338), .A4(new_n602), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n713), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT31), .B1(new_n720), .B2(new_n679), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT97), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n706), .ZN(new_n724));
  INV_X1    g0524(.A(new_n712), .ZN(new_n725));
  INV_X1    g0525(.A(new_n492), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n715), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n712), .A2(new_n728), .B1(new_n717), .B2(new_n718), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n679), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT97), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n679), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n631), .A2(new_n560), .A3(new_n595), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n723), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n648), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT98), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n641), .A4(new_n643), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n658), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT98), .B1(new_n650), .B2(new_n640), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(KEYINPUT29), .B(new_n736), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT29), .ZN(new_n748));
  INV_X1    g0548(.A(new_n659), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n749), .B2(new_n679), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n740), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n705), .B1(new_n751), .B2(G1), .ZN(G364));
  INV_X1    g0552(.A(new_n683), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n220), .A2(G13), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n754), .A2(G45), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT99), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT99), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(G1), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n696), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n682), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n219), .B1(G20), .B2(new_n324), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n695), .A2(new_n289), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n240), .A2(G45), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT100), .Z(new_n770));
  AOI211_X1 g0570(.A(new_n768), .B(new_n770), .C1(new_n306), .C2(new_n218), .ZN(new_n771));
  NAND3_X1  g0571(.A1(G355), .A2(new_n289), .A3(new_n223), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G116), .B2(new_n223), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n766), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n759), .ZN(new_n775));
  NAND2_X1  g0575(.A1(G20), .A2(G179), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT101), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n615), .A3(new_n362), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n777), .A2(new_n409), .A3(new_n362), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G58), .A2(new_n779), .B1(new_n781), .B2(G77), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n777), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n457), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n783), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n782), .B1(new_n207), .B2(new_n785), .C1(new_n209), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(G20), .A3(new_n409), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT102), .B(KEYINPUT32), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n220), .B1(new_n789), .B2(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n388), .B1(new_n796), .B2(G97), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n220), .A2(G179), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n698), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n798), .A2(new_n409), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(G107), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n794), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT103), .B(G326), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n784), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n802), .A2(G283), .ZN(new_n807));
  INV_X1    g0607(.A(new_n790), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n289), .B1(new_n808), .B2(G329), .ZN(new_n809));
  INV_X1    g0609(.A(new_n799), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(G303), .B1(new_n796), .B2(G294), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n806), .A2(new_n807), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G322), .A2(new_n779), .B1(new_n781), .B2(G311), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT33), .B(G317), .Z(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n787), .B2(new_n814), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n788), .A2(new_n804), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n775), .B1(new_n816), .B2(new_n765), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n774), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT104), .ZN(new_n819));
  INV_X1    g0619(.A(new_n764), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n682), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n761), .B1(new_n819), .B2(new_n821), .ZN(G396));
  NAND3_X1  g0622(.A1(new_n659), .A2(new_n365), .A3(new_n736), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n508), .A2(new_n521), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT82), .ZN(new_n825));
  INV_X1    g0625(.A(new_n524), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n826), .A3(new_n641), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n630), .B1(new_n684), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n652), .B2(KEYINPUT91), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n679), .B1(new_n831), .B2(new_n655), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n360), .A2(new_n363), .B1(new_n357), .B2(new_n679), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n357), .A2(new_n679), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n359), .A2(new_n342), .A3(new_n357), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n341), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n823), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n838), .A2(new_n739), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n759), .B1(new_n838), .B2(new_n739), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n765), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n763), .ZN(new_n843));
  INV_X1    g0643(.A(G303), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n785), .A2(new_n844), .B1(new_n604), .B2(new_n780), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n801), .A2(new_n698), .ZN(new_n846));
  INV_X1    g0646(.A(G311), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n388), .B1(new_n790), .B2(new_n847), .C1(new_n608), .C2(new_n795), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n846), .B(new_n848), .C1(G107), .C2(new_n810), .ZN(new_n849));
  INV_X1    g0649(.A(G283), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n787), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n845), .B(new_n851), .C1(G294), .C2(new_n779), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G143), .A2(new_n779), .B1(new_n781), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n853), .B1(new_n854), .B2(new_n785), .C1(new_n250), .C2(new_n787), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT34), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n289), .B1(new_n790), .B2(new_n857), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n207), .A2(new_n799), .B1(new_n801), .B2(new_n209), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n858), .B(new_n859), .C1(G58), .C2(new_n796), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n852), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n759), .B1(G77), .B2(new_n843), .C1(new_n861), .C2(new_n842), .ZN(new_n862));
  INV_X1    g0662(.A(new_n837), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(new_n762), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT105), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n841), .A2(new_n865), .ZN(G384));
  OR2_X1    g0666(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n867), .A2(G116), .A3(new_n221), .A4(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  OAI211_X1 g0670(.A(new_n218), .B(G77), .C1(new_n255), .C2(new_n209), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n207), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n272), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n470), .A2(new_n747), .A3(new_n750), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n672), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n460), .A2(new_n462), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT107), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n434), .A2(KEYINPUT79), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n344), .A3(new_n437), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n261), .A2(new_n277), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n429), .A2(new_n430), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n270), .B1(new_n884), .B2(new_n415), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n885), .B2(new_n431), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n879), .B1(new_n886), .B2(new_n677), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  INV_X1    g0688(.A(new_n677), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n439), .A2(KEYINPUT107), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n878), .A2(new_n887), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n454), .A2(new_n465), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n886), .A2(new_n677), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n468), .A2(new_n893), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n666), .A2(new_n665), .A3(new_n669), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n887), .A2(new_n890), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n878), .A2(new_n887), .A3(new_n890), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n891), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT108), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n899), .A2(new_n898), .B1(new_n902), .B2(new_n891), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n907), .A2(KEYINPUT108), .A3(KEYINPUT38), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n877), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n895), .B2(new_n896), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n897), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n877), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n405), .A2(new_n407), .ZN(new_n915));
  INV_X1    g0715(.A(new_n382), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n679), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n909), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n360), .A2(new_n679), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n823), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n379), .A2(new_n381), .A3(new_n679), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT106), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n917), .A2(new_n925), .A3(new_n413), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n923), .B(KEYINPUT106), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n408), .B2(new_n414), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n922), .A2(new_n912), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n666), .A2(new_n665), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n677), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n919), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n876), .B(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(G330), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n737), .A2(new_n732), .A3(new_n734), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n937), .A2(new_n837), .A3(new_n926), .A4(new_n928), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT40), .ZN(new_n939));
  INV_X1    g0739(.A(new_n897), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n910), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n737), .A2(new_n732), .A3(new_n734), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n926), .A2(new_n928), .A3(new_n837), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n906), .B2(new_n908), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(new_n946), .B2(KEYINPUT40), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n470), .A2(new_n937), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n936), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n935), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n272), .B2(new_n754), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n935), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n874), .B1(new_n953), .B2(new_n954), .ZN(G367));
  OAI221_X1 g0755(.A(new_n766), .B1(new_n223), .B2(new_n354), .C1(new_n235), .C2(new_n768), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n956), .A2(new_n759), .ZN(new_n957));
  INV_X1    g0757(.A(G317), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n388), .B1(new_n790), .B2(new_n958), .C1(new_n801), .C2(new_n608), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT112), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n784), .A2(G311), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n810), .A2(G116), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT46), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n962), .A2(new_n963), .B1(G107), .B2(new_n796), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n961), .B(new_n964), .C1(new_n844), .C2(new_n778), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n962), .A2(new_n963), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT111), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G294), .A2(new_n786), .B1(new_n781), .B2(G283), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n960), .C2(new_n959), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n786), .A2(G159), .B1(new_n784), .B2(G143), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n250), .B2(new_n778), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n799), .A2(new_n255), .B1(new_n854), .B2(new_n790), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT113), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n801), .A2(new_n293), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n795), .A2(new_n209), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n975), .A2(new_n976), .A3(new_n388), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n974), .B(new_n977), .C1(new_n207), .C2(new_n780), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n970), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n736), .B1(new_n549), .B2(new_n551), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n648), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n559), .B2(new_n981), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n957), .B1(new_n980), .B2(new_n842), .C1(new_n987), .C2(new_n820), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n656), .B1(new_n506), .B2(new_n736), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n638), .A2(new_n736), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n693), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n991), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n691), .A2(new_n692), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n997), .B(KEYINPUT44), .C1(new_n998), .C2(new_n687), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT44), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n693), .B2(new_n991), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n689), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n996), .A2(new_n1002), .A3(new_n690), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n691), .B(new_n692), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT110), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n683), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n683), .B(new_n1008), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n751), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n751), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n696), .B(KEYINPUT41), .Z(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n758), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n998), .A2(new_n991), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT42), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n521), .B1(new_n997), .B2(new_n595), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n736), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(KEYINPUT42), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT43), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n986), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1027), .A2(new_n1028), .B1(new_n690), .B2(new_n997), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1028), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n690), .A2(new_n997), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n1026), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n988), .B1(new_n1016), .B2(new_n1033), .ZN(G387));
  NAND2_X1  g0834(.A1(new_n688), .A2(new_n764), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n232), .A2(new_n306), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n351), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  AOI211_X1 g0838(.A(G45), .B(new_n700), .C1(G68), .C2(G77), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n768), .B(new_n1036), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n700), .A2(new_n223), .A3(new_n289), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(G107), .B2(new_n223), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT114), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n766), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n759), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n799), .A2(new_n293), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n289), .B1(new_n790), .B2(new_n250), .C1(new_n801), .C2(new_n608), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n554), .C2(new_n796), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n786), .A2(new_n261), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n784), .A2(G159), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G50), .A2(new_n779), .B1(new_n781), .B2(G68), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n289), .B1(new_n808), .B2(new_n805), .ZN(new_n1053));
  INV_X1    g0853(.A(G294), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n799), .A2(new_n1054), .B1(new_n795), .B2(new_n850), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n786), .A2(G311), .B1(new_n784), .B2(G322), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n844), .B2(new_n780), .C1(new_n958), .C2(new_n778), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1053), .B1(new_n604), .B2(new_n801), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1052), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1045), .B1(new_n1064), .B2(new_n765), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1011), .A2(new_n758), .B1(new_n1035), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1012), .A2(new_n696), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n751), .A2(new_n1011), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(G393));
  NAND3_X1  g0869(.A1(new_n1004), .A2(new_n758), .A3(new_n1005), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n243), .A2(new_n767), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n765), .B(new_n764), .C1(G97), .C2(new_n695), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n775), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n785), .A2(new_n250), .B1(new_n791), .B2(new_n778), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n780), .A2(new_n351), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n388), .B(new_n846), .C1(G143), .C2(new_n808), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n209), .B2(new_n799), .C1(new_n293), .C2(new_n795), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G50), .C2(new_n786), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n289), .B1(new_n808), .B2(G322), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n501), .B2(new_n801), .C1(new_n850), .C2(new_n799), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT115), .Z(new_n1082));
  NOR2_X1   g0882(.A1(new_n787), .A2(new_n844), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n780), .A2(new_n1054), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n795), .A2(new_n604), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n785), .A2(new_n958), .B1(new_n847), .B2(new_n778), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1075), .A2(new_n1079), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1073), .B1(new_n1089), .B2(new_n842), .C1(new_n991), .C2(new_n820), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1070), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n696), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1091), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(G390));
  NAND2_X1  g0897(.A1(new_n937), .A2(G330), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1099), .A2(KEYINPUT117), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n837), .B1(new_n1099), .B2(KEYINPUT117), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n929), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n736), .B(new_n837), .C1(new_n744), .C2(new_n746), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n921), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n944), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n740), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n738), .A2(G330), .A3(new_n837), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n929), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1098), .A2(new_n944), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT116), .B1(new_n1112), .B2(new_n922), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1110), .B1(new_n1108), .B2(new_n929), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT116), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n920), .B1(new_n832), .B2(new_n365), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n470), .A2(new_n1099), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n875), .A2(new_n672), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n364), .B(new_n679), .C1(new_n831), .C2(new_n655), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n930), .B1(new_n1123), .B2(new_n920), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n918), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1124), .A2(new_n1125), .B1(new_n909), .B2(new_n914), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1104), .A2(new_n930), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n904), .A2(new_n905), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT108), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n897), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1127), .A2(new_n1125), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1110), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(new_n1125), .A3(new_n1130), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n740), .A2(new_n1105), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n929), .B1(new_n823), .B2(new_n921), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n918), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n913), .B1(new_n1130), .B2(new_n877), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1133), .B(new_n1134), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1122), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1118), .A2(new_n1138), .A3(new_n1132), .A4(new_n1121), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n696), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n909), .A2(new_n914), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n762), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n759), .B1(new_n261), .B2(new_n843), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n801), .A2(new_n207), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n388), .B(new_n1146), .C1(G125), .C2(new_n808), .ZN(new_n1147));
  INV_X1    g0947(.A(G128), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1147), .B1(new_n791), .B2(new_n795), .C1(new_n785), .C2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT54), .B(G143), .Z(new_n1150));
  AOI22_X1  g0950(.A1(G132), .A2(new_n779), .B1(new_n781), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n799), .A2(new_n250), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n854), .C2(new_n787), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n289), .B(new_n800), .C1(G294), .C2(new_n808), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n802), .A2(G68), .B1(new_n796), .B2(G77), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n850), .C2(new_n785), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G107), .A2(new_n786), .B1(new_n781), .B2(G97), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n604), .B2(new_n778), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1149), .A2(new_n1154), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1145), .B1(new_n1160), .B2(new_n765), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1144), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n758), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1139), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1142), .A2(new_n1165), .ZN(G378));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n677), .B1(new_n310), .B2(new_n311), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n367), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n320), .A2(new_n321), .A3(new_n326), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1169), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n947), .B2(new_n936), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n939), .B1(new_n1130), .B2(new_n945), .ZN(new_n1180));
  OAI211_X1 g0980(.A(G330), .B(new_n1177), .C1(new_n1180), .C2(new_n942), .ZN(new_n1181));
  AND4_X1   g0981(.A1(new_n1167), .A2(new_n1179), .A3(new_n934), .A4(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1179), .A2(new_n1181), .B1(new_n934), .B2(new_n1167), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n762), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n759), .B1(G50), .B2(new_n843), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G97), .A2(new_n786), .B1(new_n781), .B2(new_n554), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n388), .B(new_n305), .C1(new_n790), .C2(new_n850), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n801), .A2(new_n255), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1046), .A2(new_n1188), .A3(new_n1189), .A4(new_n976), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1187), .B(new_n1190), .C1(new_n604), .C2(new_n785), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n778), .A2(new_n501), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT119), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  XOR2_X1   g0995(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G50), .B1(new_n248), .B2(new_n305), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n289), .B2(G41), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT118), .Z(new_n1200));
  AND2_X1   g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1148), .A2(new_n778), .B1(new_n780), .B2(new_n854), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n810), .A2(new_n1150), .B1(new_n796), .B2(G150), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n787), .B2(new_n857), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(G125), .C2(new_n784), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n802), .A2(G159), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G33), .B(G41), .C1(new_n808), .C2(G124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1201), .B1(new_n1196), .B2(new_n1195), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1186), .B1(new_n1212), .B2(new_n765), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1184), .A2(new_n758), .B1(new_n1185), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT122), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1120), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n875), .A2(new_n1119), .A3(KEYINPUT122), .A4(new_n672), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1138), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1143), .B1(new_n1135), .B2(new_n918), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1111), .B1(new_n1220), .B2(new_n1133), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1112), .A2(KEYINPUT116), .A3(new_n922), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1115), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1120), .B1(new_n1225), .B2(new_n1107), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1218), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n919), .A2(new_n931), .A3(new_n933), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1228), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n696), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1141), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1184), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1214), .B1(new_n1232), .B2(new_n1235), .ZN(G375));
  OAI21_X1  g1036(.A(new_n759), .B1(G68), .B2(new_n843), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n289), .B(new_n975), .C1(G303), .C2(new_n808), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n810), .A2(G97), .B1(new_n796), .B2(new_n554), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n604), .C2(new_n787), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G294), .A2(new_n784), .B1(new_n781), .B2(G107), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n850), .B2(new_n778), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n786), .A2(new_n1150), .B1(new_n781), .B2(G150), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n854), .B2(new_n778), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n799), .A2(new_n791), .B1(new_n795), .B2(new_n207), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n289), .B1(new_n790), .B2(new_n1148), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1245), .A2(new_n1189), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n785), .B2(new_n857), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n1240), .A2(new_n1242), .B1(new_n1244), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1237), .B1(new_n1249), .B2(new_n765), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n930), .B2(new_n763), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1223), .A2(new_n1224), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1163), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT123), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT123), .B(new_n1251), .C1(new_n1252), .C2(new_n1163), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1252), .A2(new_n1120), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1122), .A2(new_n1258), .A3(new_n1015), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(G381));
  NOR3_X1   g1061(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1016), .A2(new_n1033), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n988), .A3(new_n1096), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1263), .A2(G375), .A3(G378), .A4(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT124), .ZN(G407));
  AOI21_X1  g1067(.A(new_n1093), .B1(new_n1122), .B2(new_n1139), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1164), .B1(new_n1268), .B2(new_n1141), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n678), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G375), .C2(new_n1270), .ZN(G409));
  XNOR2_X1  g1071(.A(G393), .B(G396), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G390), .A2(G387), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(G390), .B2(G387), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1273), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1265), .A2(new_n1276), .A3(new_n1274), .A4(new_n1272), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G378), .B(new_n1214), .C1(new_n1232), .C2(new_n1235), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1234), .A2(new_n1184), .A3(new_n1015), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n758), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1185), .A2(new_n1213), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1269), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G213), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(G343), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT60), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1258), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1252), .A2(KEYINPUT60), .A3(new_n1120), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(new_n696), .A3(new_n1122), .A4(new_n1294), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1257), .A2(new_n1295), .A3(G384), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G384), .B1(new_n1257), .B2(new_n1295), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1288), .A2(new_n1291), .A3(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1281), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1290), .B1(new_n1282), .B2(new_n1287), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1298), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT125), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1257), .A2(new_n1295), .ZN(new_n1306));
  INV_X1    g1106(.A(G384), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1257), .A2(new_n1295), .A3(G384), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1290), .A2(G2897), .ZN(new_n1310));
  XOR2_X1   g1110(.A(new_n1310), .B(KEYINPUT126), .Z(new_n1311));
  NAND3_X1  g1111(.A1(new_n1308), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1311), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1312), .B(new_n1314), .C1(new_n1302), .C2(new_n1304), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1301), .B(new_n1303), .C1(new_n1305), .C2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1312), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1279), .B1(new_n1317), .B2(new_n1302), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  AND4_X1   g1119(.A1(new_n1319), .A2(new_n1288), .A3(new_n1291), .A4(new_n1298), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1302), .B2(new_n1298), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1318), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1316), .B1(new_n1322), .B2(new_n1324), .ZN(G405));
  NAND2_X1  g1125(.A1(G375), .A2(new_n1269), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1282), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1298), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1327), .A2(new_n1298), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1323), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1330), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1324), .A3(new_n1328), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(G402));
endmodule


