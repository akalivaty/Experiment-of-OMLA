//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  OR3_X1    g001(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT26), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(KEYINPUT26), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT68), .B(G190gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n211), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT23), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n228), .B(new_n231), .C1(new_n209), .C2(new_n206), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n226), .A2(KEYINPUT25), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n236), .A2(new_n221), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n211), .A2(KEYINPUT64), .A3(new_n223), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT64), .B1(new_n211), .B2(new_n223), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n232), .B1(new_n240), .B2(KEYINPUT65), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n237), .B(new_n242), .C1(new_n238), .C2(new_n239), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(KEYINPUT69), .B(new_n234), .C1(new_n244), .C2(KEYINPUT25), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT25), .B1(new_n241), .B2(new_n243), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  AOI211_X1 g047(.A(new_n248), .B(new_n232), .C1(new_n222), .C2(new_n225), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n218), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n202), .B1(new_n251), .B2(KEYINPUT29), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT79), .ZN(new_n253));
  INV_X1    g052(.A(new_n218), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n247), .B2(new_n249), .ZN(new_n255));
  INV_X1    g054(.A(new_n202), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n253), .B(new_n202), .C1(new_n251), .C2(KEYINPUT29), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G197gat), .B(G204gat), .Z(new_n261));
  AOI21_X1  g060(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT78), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT77), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n264), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n267), .B2(new_n263), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n274), .A3(new_n202), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n245), .A2(new_n250), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n254), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n277), .B2(new_n202), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(new_n271), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(new_n273), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n270), .B1(new_n258), .B2(new_n259), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT80), .B1(new_n286), .B2(new_n279), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n281), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n280), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n284), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT30), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(G127gat), .A2(G134gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(G127gat), .A2(G134gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  AOI211_X1 g097(.A(KEYINPUT1), .B(new_n297), .C1(KEYINPUT74), .C2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(KEYINPUT74), .B2(new_n298), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n298), .B2(KEYINPUT73), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(KEYINPUT73), .B2(new_n298), .ZN(new_n302));
  XOR2_X1   g101(.A(KEYINPUT72), .B(G127gat), .Z(new_n303));
  AOI21_X1  g102(.A(new_n296), .B1(new_n303), .B2(G134gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G155gat), .ZN(new_n307));
  INV_X1    g106(.A(G162gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT2), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n309), .A2(KEYINPUT84), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(KEYINPUT84), .ZN(new_n311));
  XOR2_X1   g110(.A(G155gat), .B(G162gat), .Z(new_n312));
  NOR3_X1   g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT82), .B(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G141gat), .ZN(new_n315));
  INV_X1    g114(.A(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G148gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(KEYINPUT83), .A3(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n313), .B(new_n318), .C1(KEYINPUT83), .C2(new_n315), .ZN(new_n319));
  XNOR2_X1  g118(.A(G141gat), .B(G148gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n309), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n312), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n306), .B1(new_n325), .B2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n319), .B2(new_n324), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n325), .ZN(new_n330));
  INV_X1    g129(.A(new_n306), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT4), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n325), .A2(new_n306), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT85), .B(KEYINPUT4), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n329), .A2(new_n334), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n336), .B1(new_n325), .B2(new_n306), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n339), .B(new_n343), .C1(new_n332), .C2(new_n333), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n326), .A2(new_n328), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n347), .B2(new_n335), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT5), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n342), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G57gat), .B(G85gat), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT87), .ZN(new_n352));
  XOR2_X1   g151(.A(G1gat), .B(G29gat), .Z(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n342), .B(new_n356), .C1(new_n346), .C2(new_n349), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n350), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n292), .A2(new_n294), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT29), .B1(new_n266), .B2(new_n269), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n325), .B1(new_n365), .B2(KEYINPUT3), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n274), .B1(new_n325), .B2(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n271), .ZN(new_n368));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n265), .B(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n263), .A2(new_n264), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n274), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n327), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n325), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n370), .B1(new_n378), .B2(new_n368), .ZN(new_n379));
  OR3_X1    g178(.A1(new_n372), .A2(new_n379), .A3(G22gat), .ZN(new_n380));
  OAI21_X1  g179(.A(G22gat), .B1(new_n372), .B2(new_n379), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT88), .ZN(new_n382));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT31), .B(G50gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  AND4_X1   g184(.A1(new_n380), .A2(new_n382), .A3(new_n381), .A4(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n382), .A2(new_n385), .B1(new_n380), .B2(new_n381), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n277), .A2(new_n331), .ZN(new_n389));
  INV_X1    g188(.A(G227gat), .ZN(new_n390));
  INV_X1    g189(.A(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n251), .A2(new_n306), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(G71gat), .B(G99gat), .Z(new_n395));
  XNOR2_X1  g194(.A(G15gat), .B(G43gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT33), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(KEYINPUT32), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT75), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n394), .A2(new_n401), .A3(KEYINPUT32), .A4(new_n398), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT34), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n393), .ZN(new_n405));
  INV_X1    g204(.A(new_n392), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI211_X1 g206(.A(KEYINPUT34), .B(new_n392), .C1(new_n389), .C2(new_n393), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(new_n394), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n410), .B(new_n397), .C1(new_n411), .C2(KEYINPUT33), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n403), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n403), .A2(new_n412), .ZN(new_n414));
  INV_X1    g213(.A(new_n409), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n388), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT35), .B1(new_n364), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n413), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n386), .A2(new_n387), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n293), .B1(new_n288), .B2(new_n290), .ZN(new_n422));
  INV_X1    g221(.A(new_n294), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT35), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n421), .A2(new_n424), .A3(new_n425), .A4(new_n363), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n418), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n286), .A2(new_n279), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n361), .B(new_n362), .C1(new_n428), .C2(new_n285), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n285), .B1(new_n428), .B2(KEYINPUT37), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n258), .A2(new_n270), .A3(new_n259), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT37), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n278), .B2(new_n271), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT38), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n429), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n281), .A2(KEYINPUT37), .A3(new_n287), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT38), .B1(new_n437), .B2(new_n430), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  OR3_X1    g239(.A1(new_n347), .A2(new_n340), .A3(new_n335), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT39), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT89), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n334), .A2(new_n338), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n340), .B1(new_n444), .B2(new_n345), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n446), .A3(KEYINPUT39), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n356), .B1(new_n445), .B2(KEYINPUT39), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n440), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n445), .A2(KEYINPUT39), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT40), .A4(new_n356), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n450), .A2(new_n453), .A3(new_n358), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n422), .B2(new_n423), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n455), .A3(new_n388), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n364), .A2(new_n420), .ZN(new_n457));
  NAND2_X1  g256(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n419), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n416), .B(new_n413), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n456), .A2(new_n457), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n427), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G71gat), .A2(G78gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT9), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT95), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT95), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  INV_X1    g272(.A(G57gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G64gat), .ZN(new_n475));
  INV_X1    g274(.A(G64gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G57gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n471), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G71gat), .B(G78gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT96), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n474), .A3(G64gat), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT96), .B1(new_n476), .B2(G57gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n476), .A2(G57gat), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(new_n480), .A3(new_n473), .A4(new_n471), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G231gat), .A2(G233gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G127gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT16), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(G1gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n497), .B(new_n498), .C1(G1gat), .C2(new_n495), .ZN(new_n499));
  NOR2_X1   g298(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n500), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT21), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n489), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n494), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G183gat), .B(G211gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT98), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(new_n307), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n508), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n506), .B(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT41), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n515), .B(KEYINPUT99), .Z(new_n516));
  XNOR2_X1  g315(.A(G134gat), .B(G162gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  INV_X1    g320(.A(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT14), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT92), .B1(new_n520), .B2(KEYINPUT15), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n526), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n530), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n527), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n521), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n532), .A2(KEYINPUT91), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n528), .A4(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n531), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT7), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(G85gat), .A3(G92gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  INV_X1    g347(.A(G92gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n546), .A2(new_n550), .A3(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n541), .A2(new_n556), .B1(new_n514), .B2(new_n513), .ZN(new_n557));
  INV_X1    g356(.A(new_n539), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n532), .A2(KEYINPUT91), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n520), .A2(KEYINPUT15), .A3(new_n528), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n529), .A2(new_n530), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n534), .A2(new_n561), .B1(new_n562), .B2(new_n521), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT93), .B1(new_n541), .B2(KEYINPUT17), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n541), .A2(KEYINPUT17), .B1(new_n555), .B2(new_n554), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n557), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT100), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AOI211_X1 g373(.A(new_n572), .B(new_n557), .C1(new_n568), .C2(new_n569), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n519), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n573), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n556), .B1(new_n563), .B2(new_n565), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n578), .B1(new_n567), .B2(new_n566), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n572), .B1(new_n579), .B2(new_n557), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n580), .A3(new_n518), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n512), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n489), .A2(new_n556), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n482), .A2(new_n488), .A3(new_n554), .A4(new_n555), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(KEYINPUT101), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n489), .A2(new_n587), .A3(new_n556), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT102), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT10), .B1(new_n586), .B2(new_n588), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n585), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n592), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n599), .A2(new_n601), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n591), .B(KEYINPUT104), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n605), .A2(new_n606), .B1(new_n592), .B2(new_n589), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n596), .B(KEYINPUT103), .Z(new_n608));
  AOI21_X1  g407(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n583), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n541), .A2(KEYINPUT17), .B1(new_n502), .B2(new_n501), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n541), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G229gat), .A2(G233gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n503), .A2(new_n541), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n620), .A2(KEYINPUT18), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n503), .B(new_n541), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n621), .B(KEYINPUT13), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n622), .B1(new_n568), .B2(new_n617), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT18), .B1(new_n629), .B2(new_n621), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n616), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT18), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n616), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n634), .A2(new_n624), .A3(new_n627), .A4(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n610), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n467), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n363), .B(KEYINPUT105), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g442(.A1(new_n292), .A2(new_n294), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  AND3_X1   g444(.A1(new_n639), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G8gat), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n639), .B2(new_n644), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT42), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n639), .A2(new_n644), .A3(new_n645), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT106), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n655), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(G1325gat));
  INV_X1    g456(.A(new_n639), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n658), .A2(G15gat), .A3(new_n419), .ZN(new_n659));
  OAI21_X1  g458(.A(G15gat), .B1(new_n658), .B2(new_n465), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(G1326gat));
  NAND2_X1  g460(.A1(new_n639), .A2(new_n420), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  INV_X1    g463(.A(new_n512), .ZN(new_n665));
  INV_X1    g464(.A(new_n609), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n665), .A2(new_n637), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n467), .A2(new_n582), .A3(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(G29gat), .A3(new_n640), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT45), .Z(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n364), .A2(new_n420), .B1(new_n459), .B2(new_n464), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n456), .A2(new_n672), .B1(new_n418), .B2(new_n426), .ZN(new_n673));
  INV_X1    g472(.A(new_n582), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n467), .A2(KEYINPUT44), .A3(new_n582), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n667), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n640), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n670), .A2(new_n679), .ZN(G1328gat));
  OAI21_X1  g479(.A(G36gat), .B1(new_n678), .B2(new_n424), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n668), .A2(G36gat), .A3(new_n424), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT46), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1329gat));
  NOR2_X1   g483(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n419), .A2(G43gat), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n467), .A2(new_n582), .A3(new_n667), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT107), .ZN(new_n691));
  INV_X1    g490(.A(new_n465), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n676), .A3(new_n692), .A4(new_n667), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  AOI211_X1 g493(.A(new_n685), .B(new_n688), .C1(new_n691), .C2(new_n694), .ZN(new_n695));
  AND4_X1   g494(.A1(new_n686), .A2(new_n691), .A3(new_n694), .A4(new_n687), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(G1330gat));
  INV_X1    g496(.A(G50gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n668), .B2(new_n388), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n388), .A2(new_n698), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n678), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT48), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n704), .B(new_n699), .C1(new_n678), .C2(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1331gat));
  NAND2_X1  g505(.A1(new_n631), .A2(new_n636), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n609), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n583), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT109), .B1(new_n673), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n467), .A2(new_n711), .A3(new_n583), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n640), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(new_n474), .ZN(G1332gat));
  NOR2_X1   g514(.A1(new_n713), .A2(new_n424), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n713), .B2(new_n465), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n419), .B(KEYINPUT110), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(G71gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n710), .A2(new_n712), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1334gat));
  NOR2_X1   g526(.A1(new_n713), .A2(new_n388), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(G78gat), .Z(G1335gat));
  AND2_X1   g528(.A1(new_n708), .A2(new_n512), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n677), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731), .B2(new_n640), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n665), .A2(new_n707), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n467), .A2(new_n582), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n736), .A2(new_n548), .A3(new_n666), .A4(new_n641), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n737), .ZN(G1336gat));
  NOR2_X1   g537(.A1(new_n424), .A2(new_n609), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n549), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n675), .A2(new_n676), .A3(new_n644), .A4(new_n730), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G92gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n734), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n734), .A2(new_n747), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n750), .A2(new_n741), .B1(G92gat), .B2(new_n744), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n746), .B1(new_n751), .B2(new_n743), .ZN(G1337gat));
  OAI21_X1  g551(.A(G99gat), .B1(new_n731), .B2(new_n465), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n419), .A2(G99gat), .A3(new_n609), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1338gat));
  NOR3_X1   g555(.A1(new_n388), .A2(G106gat), .A3(new_n609), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT53), .B1(new_n736), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n675), .A2(new_n676), .A3(new_n420), .A4(new_n730), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G106gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n759), .A2(new_n760), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n757), .B1(new_n748), .B2(new_n749), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n759), .A2(G106gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  INV_X1    g569(.A(new_n606), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n770), .B(new_n771), .C1(new_n599), .C2(new_n601), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(new_n597), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n599), .A2(new_n601), .A3(new_n771), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT54), .B(new_n602), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n589), .A2(new_n600), .ZN(new_n777));
  INV_X1    g576(.A(new_n601), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n778), .A3(new_n606), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT114), .ZN(new_n780));
  OAI211_X1 g579(.A(KEYINPUT55), .B(new_n773), .C1(new_n776), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n603), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(KEYINPUT114), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n774), .A2(new_n775), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n784), .A2(new_n785), .A3(KEYINPUT54), .A4(new_n602), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT55), .B1(new_n786), .B2(new_n773), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(KEYINPUT115), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(KEYINPUT115), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n707), .B(new_n783), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n615), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n629), .A2(new_n621), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n625), .A2(new_n626), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n666), .A2(new_n636), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n674), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n582), .A2(new_n636), .A3(new_n794), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n798), .B(new_n783), .C1(new_n789), .C2(new_n788), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n665), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n610), .A2(new_n707), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n641), .A2(new_n424), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n417), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G113gat), .B1(new_n805), .B2(new_n637), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(KEYINPUT116), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n637), .A2(G113gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(G1340gat));
  OAI21_X1  g608(.A(G120gat), .B1(new_n805), .B2(new_n609), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n609), .A2(G120gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT117), .Z(G1341gat));
  NOR2_X1   g613(.A1(new_n805), .A2(new_n512), .ZN(new_n815));
  INV_X1    g614(.A(new_n303), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT118), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n815), .B(new_n817), .Z(G1342gat));
  NOR3_X1   g617(.A1(new_n805), .A2(G134gat), .A3(new_n674), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  OAI21_X1  g621(.A(G134gat), .B1(new_n805), .B2(new_n674), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(G1343gat));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n802), .A2(new_n825), .A3(new_n420), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n692), .A2(new_n803), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT119), .B1(new_n782), .B2(new_n787), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n773), .B1(new_n776), .B2(new_n780), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n603), .A4(new_n781), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n707), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n582), .B1(new_n834), .B2(new_n795), .ZN(new_n835));
  INV_X1    g634(.A(new_n799), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n512), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n801), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n388), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n826), .B(new_n827), .C1(new_n825), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G141gat), .B1(new_n840), .B2(new_n637), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n802), .A2(new_n420), .A3(new_n827), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n316), .A3(new_n707), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT58), .ZN(G1344gat));
  NOR2_X1   g644(.A1(new_n314), .A2(KEYINPUT59), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n840), .B2(new_n609), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848));
  INV_X1    g647(.A(new_n795), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n782), .A2(new_n787), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n637), .B1(new_n850), .B2(new_n832), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n828), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n799), .B1(new_n852), .B2(new_n582), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n801), .B1(new_n853), .B2(new_n512), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT120), .B(new_n825), .C1(new_n854), .C2(new_n388), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n857));
  OAI211_X1 g656(.A(KEYINPUT57), .B(new_n420), .C1(new_n800), .C2(new_n801), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n666), .A3(new_n827), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G148gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n848), .B1(new_n861), .B2(KEYINPUT59), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT121), .B(new_n863), .C1(new_n860), .C2(G148gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n847), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n314), .A3(new_n666), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1345gat));
  OAI21_X1  g666(.A(G155gat), .B1(new_n840), .B2(new_n512), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n842), .A2(new_n307), .A3(new_n665), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  NAND3_X1  g669(.A1(new_n842), .A2(new_n308), .A3(new_n582), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT122), .Z(new_n872));
  OAI21_X1  g671(.A(G162gat), .B1(new_n840), .B2(new_n674), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1347gat));
  NAND3_X1  g673(.A1(new_n644), .A2(new_n640), .A3(KEYINPUT123), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT123), .B1(new_n644), .B2(new_n640), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n722), .A2(new_n420), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n802), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n802), .A2(new_n878), .A3(KEYINPUT124), .A4(new_n879), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n707), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n802), .A2(new_n421), .A3(new_n640), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n424), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n637), .A2(G169gat), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n884), .A2(G169gat), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT125), .ZN(G1348gat));
  AND2_X1   g688(.A1(new_n882), .A2(new_n883), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n666), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n739), .A2(new_n230), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n891), .A2(new_n230), .B1(new_n885), .B2(new_n892), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n882), .A2(new_n665), .A3(new_n883), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G183gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n886), .A2(new_n214), .A3(new_n665), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n886), .A2(new_n213), .A3(new_n582), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n890), .A2(new_n582), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(G190gat), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT61), .B(new_n235), .C1(new_n890), .C2(new_n582), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(G1351gat));
  INV_X1    g703(.A(G197gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n876), .A2(new_n692), .A3(new_n877), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n859), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(new_n707), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n802), .A2(new_n420), .A3(new_n465), .A4(new_n640), .ZN(new_n909));
  NOR4_X1   g708(.A1(new_n909), .A2(G197gat), .A3(new_n424), .A4(new_n637), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n908), .A2(KEYINPUT126), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT126), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1352gat));
  NOR4_X1   g712(.A1(new_n909), .A2(G204gat), .A3(new_n424), .A4(new_n609), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT62), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n859), .A2(new_n906), .A3(new_n666), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G204gat), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1353gat));
  NOR2_X1   g717(.A1(new_n909), .A2(new_n424), .ZN(new_n919));
  INV_X1    g718(.A(G211gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n665), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n907), .A2(new_n665), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n922), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT63), .B1(new_n922), .B2(G211gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1354gat));
  AOI21_X1  g724(.A(G218gat), .B1(new_n919), .B2(new_n582), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n582), .A2(G218gat), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT127), .Z(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n907), .B2(new_n928), .ZN(G1355gat));
endmodule


