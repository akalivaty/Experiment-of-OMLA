//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G214), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT67), .B(G131), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n194), .B(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n197), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT76), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT16), .B1(new_n204), .B2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n206), .A2(KEYINPUT74), .A3(G140), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(KEYINPUT74), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n209), .B2(KEYINPUT16), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n203), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n204), .A2(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT74), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n215), .B(KEYINPUT16), .C1(KEYINPUT74), .C2(new_n213), .ZN(new_n216));
  INV_X1    g030(.A(new_n205), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT76), .A3(G146), .ZN(new_n219));
  INV_X1    g033(.A(new_n208), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT19), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n209), .B2(new_n221), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n211), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n212), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n202), .B1(new_n225), .B2(KEYINPUT88), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT88), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n212), .A2(new_n219), .A3(new_n227), .A4(new_n224), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT18), .A2(G131), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n200), .B(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n220), .A2(G146), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(new_n209), .B2(G146), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n187), .B(new_n191), .C1(new_n229), .C2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n234), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n196), .A2(KEYINPUT17), .A3(new_n198), .ZN(new_n237));
  INV_X1    g051(.A(new_n202), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(KEYINPUT17), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n218), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n210), .A2(new_n211), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n190), .B(new_n236), .C1(new_n239), .C2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n234), .B1(new_n226), .B2(new_n228), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT89), .B1(new_n244), .B2(new_n190), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n235), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(G475), .A2(G902), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT20), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT20), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(new_n250), .A3(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n236), .B1(new_n239), .B2(new_n242), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(new_n190), .Z(new_n254));
  INV_X1    g068(.A(G902), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G475), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT9), .B(G234), .ZN(new_n258));
  INV_X1    g072(.A(G217), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n258), .A2(new_n259), .A3(G953), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT92), .ZN(new_n262));
  INV_X1    g076(.A(G122), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT90), .B1(new_n263), .B2(G116), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT90), .ZN(new_n265));
  INV_X1    g079(.A(G116), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G122), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT91), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n263), .A2(G116), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n268), .B2(new_n270), .ZN(new_n273));
  INV_X1    g087(.A(G107), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(new_n270), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT91), .ZN(new_n277));
  AOI21_X1  g091(.A(G107), .B1(new_n277), .B2(new_n271), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n262), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n274), .B1(new_n272), .B2(new_n273), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(G107), .A3(new_n271), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT92), .ZN(new_n282));
  INV_X1    g096(.A(G128), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT13), .B1(new_n283), .B2(G143), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G128), .B(G143), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n279), .A2(new_n282), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT95), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT93), .B(G134), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n287), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n268), .A2(KEYINPUT14), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT14), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n264), .A2(new_n267), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n270), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT94), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n296), .A2(new_n297), .A3(G107), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n296), .B2(G107), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n280), .B(new_n292), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n289), .A2(new_n290), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n290), .B1(new_n289), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n261), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n289), .A2(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT95), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n289), .A2(new_n290), .A3(new_n300), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n260), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT73), .B(G902), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n314), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n303), .A2(new_n307), .A3(new_n308), .A4(new_n316), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n193), .B(new_n308), .C1(G234), .C2(G237), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT21), .B(G898), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G952), .ZN(new_n321));
  AOI211_X1 g135(.A(G953), .B(new_n321), .C1(G234), .C2(G237), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT97), .Z(new_n325));
  AND3_X1   g139(.A1(new_n315), .A2(new_n317), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n252), .A2(new_n257), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G221), .ZN(new_n329));
  INV_X1    g143(.A(new_n258), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n255), .ZN(new_n331));
  XOR2_X1   g145(.A(G110), .B(G140), .Z(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT78), .ZN(new_n333));
  INV_X1    g147(.A(G227), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n285), .A2(G137), .ZN(new_n337));
  INV_X1    g151(.A(G137), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G134), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT11), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT66), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(new_n339), .ZN(new_n345));
  AND2_X1   g159(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n346));
  NOR2_X1   g160(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n339), .B(new_n343), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n342), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G131), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n197), .B(new_n342), .C1(new_n345), .C2(new_n349), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n274), .B2(G104), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n274), .A2(G104), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n189), .A2(KEYINPUT84), .A3(G107), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G101), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n189), .A2(G107), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT80), .B1(new_n274), .B2(G104), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n189), .A3(G107), .ZN(new_n367));
  OAI22_X1  g181(.A1(new_n189), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT83), .B(G101), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n359), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT64), .B1(new_n195), .B2(G146), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT64), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n211), .A3(G143), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n195), .A2(G146), .ZN(new_n376));
  AND4_X1   g190(.A1(G128), .A2(new_n373), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n211), .A2(G143), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT1), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G128), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n377), .A2(new_n378), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n373), .A2(new_n375), .A3(G128), .A4(new_n376), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n380), .A2(new_n376), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n283), .B1(new_n380), .B2(KEYINPUT1), .ZN(new_n387));
  OAI22_X1  g201(.A1(new_n385), .A2(KEYINPUT1), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n368), .A2(new_n365), .A3(new_n367), .ZN(new_n389));
  OR2_X1    g203(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n356), .B1(new_n390), .B2(new_n361), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n370), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n388), .B1(new_n393), .B2(new_n359), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n353), .B1(new_n384), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n353), .B(KEYINPUT12), .C1(new_n384), .C2(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n353), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT10), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n372), .B2(new_n383), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n393), .A2(KEYINPUT10), .A3(new_n388), .A4(new_n359), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n392), .B2(new_n370), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n368), .A2(new_n367), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n364), .A4(new_n365), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT81), .B1(new_n389), .B2(new_n391), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G101), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n406), .B1(new_n411), .B2(KEYINPUT82), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n413));
  INV_X1    g227(.A(G101), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(new_n369), .B2(KEYINPUT81), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n415), .B2(new_n409), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n409), .A2(new_n410), .A3(new_n405), .A4(G101), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT0), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT0), .B(G128), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n385), .A2(new_n419), .B1(new_n386), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n400), .B(new_n404), .C1(new_n417), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n399), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n402), .A2(new_n403), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n415), .A2(new_n413), .A3(new_n409), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n406), .ZN(new_n429));
  INV_X1    g243(.A(new_n423), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n336), .B1(new_n431), .B2(new_n400), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n404), .B1(new_n417), .B2(new_n423), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n353), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n336), .A2(new_n425), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G469), .B1(new_n435), .B2(G902), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  INV_X1    g251(.A(new_n336), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n434), .B2(new_n424), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n399), .A2(new_n424), .A3(new_n438), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n437), .B(new_n308), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n331), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G214), .B1(G237), .B2(G902), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n444));
  INV_X1    g258(.A(G119), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G116), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n266), .A2(G119), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT2), .B(G113), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n448), .A2(KEYINPUT69), .ZN(new_n451));
  XNOR2_X1  g265(.A(G116), .B(G119), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n450), .B1(new_n455), .B2(new_n449), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n457), .B(new_n418), .C1(new_n412), .C2(new_n416), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT5), .B1(new_n451), .B2(new_n454), .ZN(new_n459));
  OAI21_X1  g273(.A(G113), .B1(new_n446), .B2(KEYINPUT5), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n450), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n372), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n450), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n448), .A2(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n452), .A2(new_n453), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n466), .B1(new_n470), .B2(new_n460), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT85), .B1(new_n471), .B2(new_n372), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n458), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n444), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n457), .A2(new_n418), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n478), .A2(new_n429), .B1(new_n472), .B2(new_n465), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT86), .B1(new_n479), .B2(new_n475), .ZN(new_n480));
  AND4_X1   g294(.A1(KEYINPUT86), .A2(new_n458), .A3(new_n475), .A4(new_n473), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n479), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n388), .A2(G125), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n421), .A2(G125), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G224), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(G953), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT87), .Z(new_n490));
  XNOR2_X1  g304(.A(new_n487), .B(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n482), .A2(new_n484), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n474), .B2(new_n476), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n479), .A2(KEYINPUT86), .A3(new_n475), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(new_n488), .B2(G953), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n487), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n448), .A2(new_n467), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n466), .B1(new_n499), .B2(new_n460), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n463), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n475), .B(KEYINPUT8), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n501), .B(new_n502), .C1(new_n471), .C2(new_n463), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n487), .A2(new_n497), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n496), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G210), .B1(G237), .B2(G902), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n492), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n492), .B2(new_n506), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n442), .B(new_n443), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n512), .B(new_n513), .Z(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT23), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n445), .B2(G128), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n445), .A2(G128), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n283), .A2(KEYINPUT23), .A3(G119), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(G110), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT75), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n283), .A2(G119), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT24), .B(G110), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n521), .A2(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT75), .B1(new_n520), .B2(G110), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n232), .ZN(new_n529));
  AND4_X1   g343(.A1(new_n212), .A2(new_n528), .A3(new_n219), .A4(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n524), .A2(new_n525), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n520), .A2(G110), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n240), .B2(new_n241), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n515), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n534), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n528), .A2(new_n212), .A3(new_n219), .A4(new_n529), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n514), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n308), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n535), .A2(new_n538), .A3(KEYINPUT25), .A4(new_n308), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n259), .B1(new_n308), .B2(G234), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(G902), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n535), .A2(new_n538), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT77), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n421), .B1(new_n351), .B2(new_n352), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n339), .A2(KEYINPUT68), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n339), .A2(KEYINPUT68), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n337), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G131), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n352), .A2(new_n556), .A3(new_n388), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n551), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n339), .B1(new_n346), .B2(new_n347), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT66), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n341), .B1(new_n560), .B2(new_n348), .ZN(new_n561));
  INV_X1    g375(.A(G131), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n341), .B(new_n198), .C1(new_n560), .C2(new_n348), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n422), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n352), .A2(new_n556), .A3(new_n388), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(KEYINPUT30), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n558), .A2(new_n457), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n192), .A2(new_n193), .A3(G210), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n569), .B(KEYINPUT27), .Z(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT26), .B(G101), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n561), .A2(new_n197), .B1(new_n555), .B2(G131), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n353), .A2(new_n422), .B1(new_n573), .B2(new_n388), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n574), .B2(new_n456), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT31), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT70), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n580));
  NAND3_X1  g394(.A1(new_n568), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT28), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n456), .B1(new_n565), .B2(new_n566), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n583), .B2(KEYINPUT71), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n457), .B1(new_n552), .B2(new_n557), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT71), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n565), .A2(new_n456), .A3(new_n566), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n584), .A2(new_n588), .B1(new_n582), .B2(new_n587), .ZN(new_n589));
  INV_X1    g403(.A(new_n572), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n579), .B(new_n581), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(G472), .A2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT32), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT32), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n595), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n584), .A2(new_n588), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n582), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n590), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT29), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n568), .A2(new_n587), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n572), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n308), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n552), .A2(new_n557), .A3(new_n457), .ZN(new_n606));
  OAI211_X1 g420(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n606), .C2(new_n583), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT72), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n599), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n582), .B1(new_n585), .B2(new_n587), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n572), .A2(new_n601), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n605), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G472), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n550), .B1(new_n597), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n328), .A2(new_n511), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(new_n371), .ZN(G3));
  NOR2_X1   g432(.A1(new_n605), .A2(new_n310), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n622), .B(new_n623), .C1(new_n303), .C2(new_n307), .ZN(new_n624));
  AND4_X1   g438(.A1(KEYINPUT99), .A2(new_n303), .A3(new_n307), .A4(KEYINPUT33), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n619), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n309), .A2(new_n310), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n246), .A2(new_n250), .A3(new_n247), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n250), .B1(new_n246), .B2(new_n247), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n257), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(new_n631), .A3(new_n325), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n579), .A2(new_n581), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n590), .B1(new_n598), .B2(new_n599), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n633), .B(new_n308), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n633), .B1(new_n591), .B2(new_n308), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n593), .B(new_n549), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n632), .A2(new_n510), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT34), .B(G104), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  NAND2_X1  g456(.A1(new_n315), .A2(new_n317), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n643), .B(new_n257), .C1(new_n629), .C2(new_n630), .ZN(new_n644));
  INV_X1    g458(.A(new_n325), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT100), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n252), .A2(new_n257), .A3(new_n643), .A4(new_n325), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI211_X1 g464(.A(new_n510), .B(new_n639), .C1(new_n647), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT101), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n651), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n536), .A2(new_n537), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n546), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n545), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n593), .B(new_n659), .C1(new_n637), .C2(new_n638), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n327), .A2(new_n510), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT102), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  AND3_X1   g478(.A1(new_n591), .A2(new_n595), .A3(new_n592), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n595), .B1(new_n591), .B2(new_n592), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n615), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n667), .A2(new_n442), .A3(new_n659), .ZN(new_n668));
  INV_X1    g482(.A(new_n443), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n492), .A2(new_n506), .ZN(new_n670));
  INV_X1    g484(.A(new_n507), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n492), .A2(new_n506), .A3(new_n507), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n322), .B1(new_n318), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n644), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n668), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  OAI21_X1  g493(.A(new_n572), .B1(new_n606), .B2(new_n583), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n576), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT103), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n255), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n681), .A2(KEYINPUT103), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n597), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n669), .A3(new_n659), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n672), .A2(new_n673), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT38), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n631), .A2(new_n643), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n688), .A2(new_n689), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n659), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n692), .A2(new_n443), .A3(new_n694), .A4(new_n686), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n690), .B(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT104), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n676), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n442), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT40), .Z(new_n701));
  NAND3_X1  g515(.A1(new_n693), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  INV_X1    g519(.A(new_n676), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n628), .A2(new_n631), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n628), .A2(new_n631), .A3(KEYINPUT106), .A4(new_n706), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n674), .A3(new_n668), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT107), .B(G146), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G48));
  NOR2_X1   g527(.A1(new_n439), .A2(new_n440), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n714), .B2(new_n605), .ZN(new_n715));
  INV_X1    g529(.A(new_n331), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n715), .A2(new_n716), .A3(new_n441), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n674), .A2(new_n667), .A3(new_n549), .A4(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n632), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT41), .B(G113), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  AOI21_X1  g535(.A(new_n718), .B1(new_n647), .B2(new_n650), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n266), .ZN(G18));
  AOI22_X1  g537(.A1(new_n249), .A2(new_n251), .B1(G475), .B2(new_n256), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n667), .A3(new_n326), .A4(new_n659), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n674), .A2(new_n717), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n445), .ZN(G21));
  NAND4_X1  g542(.A1(new_n690), .A2(new_n631), .A3(new_n443), .A4(new_n643), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n591), .A2(new_n308), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n581), .B(new_n579), .C1(new_n611), .C2(new_n590), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n730), .A2(G472), .B1(new_n592), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n717), .A2(new_n549), .A3(new_n325), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n263), .ZN(G24));
  OAI21_X1  g549(.A(new_n443), .B1(new_n508), .B2(new_n509), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n730), .A2(G472), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n731), .A2(new_n592), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n659), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n715), .A2(new_n716), .A3(new_n441), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n709), .A2(new_n741), .A3(new_n710), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT108), .B(G125), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G27));
  NAND2_X1  g558(.A1(new_n667), .A2(new_n549), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n672), .A2(new_n442), .A3(new_n443), .A4(new_n673), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n709), .A3(new_n710), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n597), .A2(KEYINPUT109), .B1(G472), .B2(new_n614), .ZN(new_n751));
  OR3_X1    g565(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT109), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n550), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n746), .A2(new_n749), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n709), .A3(new_n710), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND2_X1  g571(.A1(new_n747), .A2(new_n677), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  XNOR2_X1  g573(.A(new_n724), .B(KEYINPUT110), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n303), .A2(new_n307), .ZN(new_n761));
  INV_X1    g575(.A(new_n622), .ZN(new_n762));
  INV_X1    g576(.A(new_n623), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n303), .A2(new_n307), .A3(KEYINPUT99), .A4(KEYINPUT33), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n766), .A2(new_n619), .B1(new_n310), .B2(new_n309), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n768), .B1(new_n767), .B2(new_n631), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n770), .A2(KEYINPUT111), .A3(new_n771), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n637), .A2(new_n638), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n694), .B1(new_n776), .B2(new_n593), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n435), .A2(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n435), .A2(KEYINPUT45), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(G469), .A2(G902), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n785), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n441), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n716), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n508), .A2(new_n509), .A3(new_n669), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n792), .A2(new_n699), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n780), .A2(new_n781), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  NOR2_X1   g610(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n790), .A2(KEYINPUT47), .A3(new_n716), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n709), .A2(new_n710), .ZN(new_n800));
  INV_X1    g614(.A(new_n793), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(new_n667), .A3(new_n549), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NAND4_X1  g619(.A1(new_n628), .A2(new_n549), .A3(new_n443), .A4(new_n716), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n715), .A2(new_n441), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n686), .B(new_n806), .C1(KEYINPUT49), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(KEYINPUT49), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT112), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n808), .A2(new_n697), .A3(new_n760), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n801), .A2(new_n740), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n549), .A2(new_n812), .A3(new_n322), .A4(new_n687), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n724), .A3(new_n767), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n323), .B1(new_n770), .B2(new_n771), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n812), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n659), .A3(new_n732), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n732), .A2(new_n549), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n691), .A2(new_n443), .A3(new_n740), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT50), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n807), .A2(new_n716), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n797), .A2(new_n798), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n817), .A2(new_n822), .A3(new_n793), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n816), .A3(new_n819), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n825), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n724), .A2(new_n767), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n321), .B(G953), .C1(new_n813), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n817), .A2(new_n822), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n836), .B1(new_n837), .B2(new_n726), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n818), .A2(new_n753), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT48), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n840), .A2(new_n841), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n839), .B2(new_n842), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n838), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n831), .A2(new_n834), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n745), .A2(new_n327), .A3(new_n510), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n640), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n639), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n511), .A2(new_n835), .A3(new_n851), .A4(new_n325), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n617), .A3(KEYINPUT113), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n648), .A2(new_n510), .A3(new_n639), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT114), .B1(new_n661), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n660), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n328), .A2(new_n511), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n511), .A2(new_n851), .A3(new_n646), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n850), .A2(new_n853), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n725), .A2(new_n726), .B1(new_n729), .B2(new_n733), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n722), .A2(new_n862), .A3(new_n719), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n746), .A2(new_n739), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n709), .A2(new_n710), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n793), .A2(new_n667), .A3(new_n549), .A4(new_n442), .ZN(new_n866));
  INV_X1    g680(.A(new_n677), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n643), .A2(new_n676), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n724), .A2(new_n667), .A3(new_n659), .A4(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n866), .A2(new_n867), .B1(new_n869), .B2(new_n746), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n861), .A2(new_n756), .A3(new_n863), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n659), .A2(new_n676), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n511), .A2(new_n692), .A3(new_n686), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n711), .A2(new_n742), .A3(new_n678), .A4(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT52), .ZN(new_n876));
  XNOR2_X1  g690(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n872), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n850), .A2(new_n853), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n855), .A2(new_n860), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n871), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n756), .A2(new_n863), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n875), .B(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT54), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n881), .A2(KEYINPUT116), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n861), .A2(new_n889), .A3(new_n871), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n756), .A2(new_n863), .A3(KEYINPUT53), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n888), .A2(new_n885), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n877), .B1(new_n872), .B2(new_n876), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n847), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT119), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n811), .B1(new_n897), .B2(new_n899), .ZN(G75));
  NAND2_X1  g714(.A1(new_n892), .A2(new_n893), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n605), .A3(new_n671), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n483), .B1(new_n496), .B2(new_n477), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(new_n491), .Z(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  XOR2_X1   g719(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n906));
  AND3_X1   g720(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n193), .A2(G952), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(G51));
  XOR2_X1   g725(.A(new_n785), .B(KEYINPUT57), .Z(new_n912));
  INV_X1    g726(.A(new_n895), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n894), .B1(new_n892), .B2(new_n893), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n439), .B2(new_n440), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n901), .A2(new_n605), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(new_n784), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n910), .B1(new_n916), .B2(new_n918), .ZN(G54));
  NAND4_X1  g733(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .A4(new_n605), .ZN(new_n920));
  INV_X1    g734(.A(new_n246), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n920), .A2(KEYINPUT121), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n910), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT121), .B1(new_n920), .B2(new_n921), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(G60));
  XNOR2_X1  g740(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n887), .B2(new_n895), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n930), .B2(new_n766), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n764), .B2(new_n765), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n913), .B2(new_n914), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(new_n932), .C1(new_n913), .C2(new_n914), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n931), .B1(new_n934), .B2(new_n936), .ZN(G63));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n892), .B2(new_n893), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n657), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n535), .A2(new_n538), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n923), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n938), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n941), .A2(new_n945), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n923), .A4(new_n942), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(G953), .B1(new_n319), .B2(new_n488), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n861), .A2(new_n863), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n954), .B2(G953), .ZN(new_n955));
  INV_X1    g769(.A(G898), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n903), .B1(new_n956), .B2(G953), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT125), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n955), .B(new_n958), .ZN(G69));
  INV_X1    g773(.A(new_n729), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n792), .A2(new_n699), .A3(new_n960), .A4(new_n753), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n758), .B(new_n961), .C1(new_n799), .C2(new_n803), .ZN(new_n962));
  INV_X1    g776(.A(new_n756), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n711), .A2(new_n678), .A3(new_n742), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n795), .A2(new_n966), .A3(new_n193), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n558), .A2(new_n567), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(new_n223), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(G900), .B2(G953), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n644), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n747), .B(new_n699), .C1(new_n835), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n804), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n781), .A2(new_n794), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n780), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n978), .A3(new_n964), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n704), .A2(KEYINPUT62), .A3(new_n964), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(G953), .B1(new_n976), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n969), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n971), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI221_X1 g800(.A(G953), .B1(new_n334), .B2(new_n675), .C1(new_n969), .C2(KEYINPUT126), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n971), .B(new_n987), .C1(new_n984), .C2(new_n985), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G72));
  XOR2_X1   g805(.A(new_n602), .B(KEYINPUT127), .Z(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n590), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n976), .A2(new_n983), .A3(new_n954), .ZN(new_n994));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  AOI21_X1  g810(.A(new_n993), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n954), .A2(new_n795), .A3(new_n966), .ZN(new_n998));
  AOI211_X1 g812(.A(new_n590), .B(new_n992), .C1(new_n998), .C2(new_n996), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n878), .A2(new_n886), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n603), .A2(new_n576), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n996), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n923), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n997), .A2(new_n999), .A3(new_n1003), .ZN(G57));
endmodule


