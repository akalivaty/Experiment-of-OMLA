

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U550 ( .A1(n545), .A2(n544), .ZN(G164) );
  XNOR2_X1 U551 ( .A(n518), .B(KEYINPUT69), .ZN(n582) );
  INV_X1 U552 ( .A(KEYINPUT17), .ZN(n536) );
  NOR2_X1 U553 ( .A1(n697), .A2(KEYINPUT33), .ZN(n698) );
  AND2_X1 U554 ( .A1(n740), .A2(n739), .ZN(n741) );
  BUF_X1 U555 ( .A(n702), .Z(n703) );
  BUF_X1 U556 ( .A(n706), .Z(n707) );
  NOR2_X2 U557 ( .A1(G651), .A2(n582), .ZN(n519) );
  NAND2_X2 U558 ( .A1(n609), .A2(n608), .ZN(n984) );
  XNOR2_X2 U559 ( .A(n554), .B(KEYINPUT23), .ZN(n555) );
  NOR2_X4 U560 ( .A1(n556), .A2(n555), .ZN(G160) );
  NAND2_X1 U561 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U562 ( .A(n612), .B(KEYINPUT26), .ZN(n615) );
  INV_X2 U563 ( .A(n539), .ZN(n547) );
  XNOR2_X2 U564 ( .A(G2104), .B(KEYINPUT66), .ZN(n539) );
  NOR2_X1 U565 ( .A1(n551), .A2(n517), .ZN(n552) );
  INV_X1 U566 ( .A(G651), .ZN(n528) );
  XNOR2_X1 U567 ( .A(KEYINPUT5), .B(KEYINPUT79), .ZN(n531) );
  BUF_X1 U568 ( .A(n549), .Z(n891) );
  NOR2_X1 U569 ( .A1(n516), .A2(n726), .ZN(n515) );
  NAND2_X1 U570 ( .A1(n999), .A2(n723), .ZN(n516) );
  XOR2_X1 U571 ( .A(KEYINPUT68), .B(n550), .Z(n517) );
  INV_X1 U572 ( .A(KEYINPUT101), .ZN(n660) );
  XNOR2_X1 U573 ( .A(n660), .B(KEYINPUT30), .ZN(n661) );
  INV_X1 U574 ( .A(KEYINPUT29), .ZN(n645) );
  BUF_X1 U575 ( .A(n647), .Z(n683) );
  INV_X1 U576 ( .A(KEYINPUT103), .ZN(n677) );
  XNOR2_X1 U577 ( .A(KEYINPUT78), .B(KEYINPUT4), .ZN(n526) );
  XNOR2_X1 U578 ( .A(n527), .B(n526), .ZN(n530) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n549) );
  INV_X1 U580 ( .A(KEYINPUT77), .ZN(n625) );
  XNOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n626), .B(n625), .ZN(n987) );
  XNOR2_X1 U583 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U584 ( .A(KEYINPUT80), .B(KEYINPUT6), .ZN(n525) );
  XOR2_X2 U585 ( .A(KEYINPUT65), .B(n519), .Z(n804) );
  NAND2_X1 U586 ( .A1(n804), .A2(G51), .ZN(n523) );
  NOR2_X1 U587 ( .A1(G543), .A2(n528), .ZN(n520) );
  XOR2_X1 U588 ( .A(KEYINPUT70), .B(n520), .Z(n521) );
  XNOR2_X2 U589 ( .A(KEYINPUT1), .B(n521), .ZN(n805) );
  NAND2_X1 U590 ( .A1(G63), .A2(n805), .ZN(n522) );
  NAND2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n534) );
  NOR2_X2 U593 ( .A1(G651), .A2(G543), .ZN(n808) );
  NAND2_X1 U594 ( .A1(G89), .A2(n808), .ZN(n527) );
  NOR2_X2 U595 ( .A1(n582), .A2(n528), .ZN(n809) );
  NAND2_X1 U596 ( .A1(G76), .A2(n809), .ZN(n529) );
  NAND2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n532) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT7), .B(n535), .Z(G168) );
  XOR2_X1 U600 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X2 U601 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XNOR2_X2 U602 ( .A(n537), .B(n536), .ZN(n888) );
  NAND2_X1 U603 ( .A1(n888), .A2(G138), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT90), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n891), .A2(G114), .ZN(n543) );
  NOR2_X2 U606 ( .A1(n547), .A2(G2105), .ZN(n702) );
  NAND2_X1 U607 ( .A1(G102), .A2(n702), .ZN(n541) );
  AND2_X1 U608 ( .A1(G2105), .A2(n547), .ZN(n706) );
  NAND2_X1 U609 ( .A1(G126), .A2(n706), .ZN(n540) );
  AND2_X1 U610 ( .A1(n541), .A2(n540), .ZN(n542) );
  AND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n888), .A2(G137), .ZN(n553) );
  AND2_X1 U613 ( .A1(G2105), .A2(G125), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT67), .ZN(n551) );
  NAND2_X1 U616 ( .A1(G113), .A2(n549), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G101), .A2(n702), .ZN(n554) );
  NAND2_X1 U619 ( .A1(G91), .A2(n808), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT72), .B(n557), .Z(n562) );
  NAND2_X1 U621 ( .A1(n804), .A2(G53), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G65), .A2(n805), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT73), .B(n560), .Z(n561) );
  NOR2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n809), .A2(G78), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(G299) );
  NAND2_X1 U628 ( .A1(n804), .A2(G52), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G64), .A2(n805), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G90), .A2(n808), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G77), .A2(n809), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(G171) );
  NAND2_X1 U636 ( .A1(G88), .A2(n808), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G75), .A2(n809), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n804), .A2(G50), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G62), .A2(n805), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(G166) );
  INV_X1 U643 ( .A(G166), .ZN(G303) );
  NAND2_X1 U644 ( .A1(G49), .A2(n804), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U647 ( .A(KEYINPUT85), .B(n580), .Z(n581) );
  NOR2_X1 U648 ( .A1(n805), .A2(n581), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n582), .A2(G87), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(G288) );
  NAND2_X1 U651 ( .A1(G86), .A2(n808), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G61), .A2(n805), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n809), .A2(G73), .ZN(n587) );
  XOR2_X1 U655 ( .A(KEYINPUT2), .B(n587), .Z(n588) );
  NOR2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n804), .A2(G48), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(G305) );
  NAND2_X1 U659 ( .A1(G85), .A2(n808), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G60), .A2(n805), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G47), .A2(n804), .ZN(n594) );
  XNOR2_X1 U663 ( .A(KEYINPUT71), .B(n594), .ZN(n595) );
  NOR2_X1 U664 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n809), .A2(G72), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(G290) );
  NAND2_X1 U667 ( .A1(G56), .A2(n805), .ZN(n599) );
  XOR2_X1 U668 ( .A(KEYINPUT14), .B(n599), .Z(n605) );
  NAND2_X1 U669 ( .A1(n808), .A2(G81), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT12), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G68), .A2(n809), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT13), .B(n603), .Z(n604) );
  NOR2_X2 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U675 ( .A(KEYINPUT74), .B(n606), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n804), .A2(G43), .ZN(n607) );
  XOR2_X1 U677 ( .A(KEYINPUT75), .B(n607), .Z(n608) );
  NAND2_X1 U678 ( .A1(G160), .A2(G40), .ZN(n699) );
  INV_X1 U679 ( .A(n699), .ZN(n611) );
  NOR2_X2 U680 ( .A1(G164), .A2(G1384), .ZN(n701) );
  NAND2_X1 U681 ( .A1(n611), .A2(n701), .ZN(n655) );
  INV_X2 U682 ( .A(n655), .ZN(n647) );
  NAND2_X1 U683 ( .A1(n683), .A2(G1996), .ZN(n612) );
  BUF_X1 U684 ( .A(n655), .Z(n613) );
  NAND2_X1 U685 ( .A1(n613), .A2(G1341), .ZN(n614) );
  NOR2_X2 U686 ( .A1(n984), .A2(n616), .ZN(n632) );
  NAND2_X1 U687 ( .A1(G54), .A2(n804), .ZN(n623) );
  NAND2_X1 U688 ( .A1(n809), .A2(G79), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G66), .A2(n805), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n808), .A2(G92), .ZN(n619) );
  XOR2_X1 U692 ( .A(KEYINPUT76), .B(n619), .Z(n620) );
  NOR2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT15), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n632), .A2(n987), .ZN(n631) );
  XNOR2_X2 U697 ( .A(n647), .B(KEYINPUT98), .ZN(n649) );
  NAND2_X1 U698 ( .A1(G2067), .A2(n649), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G1348), .A2(n613), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n629), .B(KEYINPUT100), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n634) );
  OR2_X1 U703 ( .A1(n632), .A2(n987), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n639) );
  NAND2_X1 U705 ( .A1(G2072), .A2(n649), .ZN(n635) );
  XNOR2_X2 U706 ( .A(n635), .B(KEYINPUT27), .ZN(n637) );
  INV_X1 U707 ( .A(G1956), .ZN(n1008) );
  NOR2_X1 U708 ( .A1(n649), .A2(n1008), .ZN(n636) );
  NOR2_X2 U709 ( .A1(n637), .A2(n636), .ZN(n640) );
  INV_X1 U710 ( .A(G299), .ZN(n996) );
  NAND2_X1 U711 ( .A1(n640), .A2(n996), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n644) );
  NOR2_X1 U713 ( .A1(n640), .A2(n996), .ZN(n642) );
  INV_X1 U714 ( .A(KEYINPUT28), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(n645), .ZN(n654) );
  NOR2_X1 U718 ( .A1(n647), .A2(G1961), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n648), .B(KEYINPUT97), .ZN(n651) );
  XNOR2_X1 U720 ( .A(G2078), .B(KEYINPUT25), .ZN(n962) );
  NAND2_X1 U721 ( .A1(n649), .A2(n962), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT99), .B(n652), .Z(n664) );
  NAND2_X1 U724 ( .A1(n664), .A2(G171), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n654), .A2(n653), .ZN(n670) );
  INV_X1 U726 ( .A(KEYINPUT96), .ZN(n657) );
  NAND2_X1 U727 ( .A1(G8), .A2(n655), .ZN(n736) );
  NOR2_X1 U728 ( .A1(G1966), .A2(n736), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(n687) );
  NAND2_X1 U730 ( .A1(G2084), .A2(G8), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n658), .A2(n736), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n687), .A2(n659), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X1 U734 ( .A1(G168), .A2(n663), .ZN(n666) );
  NOR2_X1 U735 ( .A1(G171), .A2(n664), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U737 ( .A(KEYINPUT31), .B(n667), .ZN(n668) );
  INV_X1 U738 ( .A(n668), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n681) );
  NAND2_X1 U740 ( .A1(n681), .A2(G286), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(KEYINPUT102), .ZN(n676) );
  NOR2_X1 U742 ( .A1(G1971), .A2(n736), .ZN(n673) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n613), .ZN(n672) );
  NOR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n674), .A2(G303), .ZN(n675) );
  NAND2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n679), .A2(G8), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n680), .B(KEYINPUT32), .ZN(n731) );
  BUF_X1 U750 ( .A(n681), .Z(n682) );
  INV_X1 U751 ( .A(n682), .ZN(n686) );
  NAND2_X1 U752 ( .A1(G8), .A2(n683), .ZN(n684) );
  NOR2_X1 U753 ( .A1(G2084), .A2(n684), .ZN(n685) );
  NOR2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n730) );
  NAND2_X1 U756 ( .A1(G288), .A2(G1976), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n689), .B(KEYINPUT104), .ZN(n986) );
  AND2_X1 U758 ( .A1(n730), .A2(n986), .ZN(n690) );
  AND2_X1 U759 ( .A1(n731), .A2(n690), .ZN(n694) );
  INV_X1 U760 ( .A(n986), .ZN(n692) );
  NOR2_X1 U761 ( .A1(G1976), .A2(G288), .ZN(n724) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n724), .A2(n691), .ZN(n997) );
  NOR2_X1 U764 ( .A1(n692), .A2(n997), .ZN(n693) );
  NOR2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U766 ( .A1(n695), .A2(n736), .ZN(n696) );
  XNOR2_X1 U767 ( .A(n696), .B(KEYINPUT64), .ZN(n697) );
  INV_X1 U768 ( .A(n698), .ZN(n727) );
  XOR2_X1 U769 ( .A(G1981), .B(G305), .Z(n999) );
  BUF_X1 U770 ( .A(n699), .Z(n700) );
  NOR2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n772) );
  NAND2_X1 U772 ( .A1(G107), .A2(n891), .ZN(n705) );
  NAND2_X1 U773 ( .A1(G95), .A2(n703), .ZN(n704) );
  NAND2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n711) );
  NAND2_X1 U775 ( .A1(G131), .A2(n888), .ZN(n709) );
  NAND2_X1 U776 ( .A1(G119), .A2(n707), .ZN(n708) );
  NAND2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n710) );
  OR2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n901) );
  NAND2_X1 U779 ( .A1(G1991), .A2(n901), .ZN(n721) );
  NAND2_X1 U780 ( .A1(G117), .A2(n891), .ZN(n713) );
  NAND2_X1 U781 ( .A1(G129), .A2(n707), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U783 ( .A(KEYINPUT94), .B(n714), .ZN(n717) );
  NAND2_X1 U784 ( .A1(n703), .A2(G105), .ZN(n715) );
  XOR2_X1 U785 ( .A(KEYINPUT38), .B(n715), .Z(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U787 ( .A1(n888), .A2(G141), .ZN(n718) );
  NAND2_X1 U788 ( .A1(n719), .A2(n718), .ZN(n898) );
  NAND2_X1 U789 ( .A1(G1996), .A2(n898), .ZN(n720) );
  NAND2_X1 U790 ( .A1(n721), .A2(n720), .ZN(n932) );
  NAND2_X1 U791 ( .A1(n772), .A2(n932), .ZN(n722) );
  XNOR2_X1 U792 ( .A(n722), .B(KEYINPUT95), .ZN(n742) );
  INV_X1 U793 ( .A(n742), .ZN(n723) );
  NAND2_X1 U794 ( .A1(n724), .A2(KEYINPUT33), .ZN(n725) );
  NOR2_X1 U795 ( .A1(n725), .A2(n736), .ZN(n726) );
  NAND2_X1 U796 ( .A1(n727), .A2(n515), .ZN(n744) );
  NOR2_X1 U797 ( .A1(G1981), .A2(G305), .ZN(n728) );
  XOR2_X1 U798 ( .A(n728), .B(KEYINPUT24), .Z(n729) );
  OR2_X1 U799 ( .A1(n736), .A2(n729), .ZN(n740) );
  NAND2_X1 U800 ( .A1(n731), .A2(n730), .ZN(n735) );
  NOR2_X1 U801 ( .A1(G2090), .A2(G303), .ZN(n732) );
  XOR2_X1 U802 ( .A(KEYINPUT105), .B(n732), .Z(n733) );
  NAND2_X1 U803 ( .A1(G8), .A2(n733), .ZN(n734) );
  NAND2_X1 U804 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U805 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U806 ( .A(n738), .B(KEYINPUT106), .ZN(n739) );
  OR2_X2 U807 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U808 ( .A1(n744), .A2(n743), .ZN(n757) );
  XOR2_X1 U809 ( .A(G2067), .B(KEYINPUT37), .Z(n745) );
  XOR2_X1 U810 ( .A(KEYINPUT92), .B(n745), .Z(n770) );
  NAND2_X1 U811 ( .A1(G116), .A2(n891), .ZN(n747) );
  NAND2_X1 U812 ( .A1(G128), .A2(n707), .ZN(n746) );
  NAND2_X1 U813 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U814 ( .A(n748), .B(KEYINPUT35), .ZN(n753) );
  NAND2_X1 U815 ( .A1(G140), .A2(n888), .ZN(n750) );
  NAND2_X1 U816 ( .A1(G104), .A2(n703), .ZN(n749) );
  NAND2_X1 U817 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U818 ( .A(KEYINPUT34), .B(n751), .Z(n752) );
  NAND2_X1 U819 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U820 ( .A(n754), .B(KEYINPUT36), .Z(n908) );
  OR2_X1 U821 ( .A1(n770), .A2(n908), .ZN(n755) );
  XOR2_X1 U822 ( .A(KEYINPUT93), .B(n755), .Z(n768) );
  INV_X1 U823 ( .A(n768), .ZN(n951) );
  NAND2_X1 U824 ( .A1(n772), .A2(n951), .ZN(n756) );
  NAND2_X1 U825 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U826 ( .A(n758), .B(KEYINPUT107), .ZN(n761) );
  XOR2_X1 U827 ( .A(KEYINPUT91), .B(G1986), .Z(n759) );
  XNOR2_X1 U828 ( .A(G290), .B(n759), .ZN(n991) );
  NAND2_X1 U829 ( .A1(n991), .A2(n772), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n761), .A2(n760), .ZN(n775) );
  NOR2_X1 U831 ( .A1(G1996), .A2(n898), .ZN(n945) );
  NOR2_X1 U832 ( .A1(G1991), .A2(n901), .ZN(n762) );
  XOR2_X1 U833 ( .A(KEYINPUT109), .B(n762), .Z(n948) );
  NOR2_X1 U834 ( .A1(G1986), .A2(G290), .ZN(n763) );
  XNOR2_X1 U835 ( .A(KEYINPUT108), .B(n763), .ZN(n764) );
  NOR2_X1 U836 ( .A1(n948), .A2(n764), .ZN(n765) );
  NOR2_X1 U837 ( .A1(n765), .A2(n932), .ZN(n766) );
  NOR2_X1 U838 ( .A1(n945), .A2(n766), .ZN(n767) );
  XNOR2_X1 U839 ( .A(n767), .B(KEYINPUT39), .ZN(n769) );
  NAND2_X1 U840 ( .A1(n769), .A2(n768), .ZN(n771) );
  NAND2_X1 U841 ( .A1(n770), .A2(n908), .ZN(n933) );
  NAND2_X1 U842 ( .A1(n771), .A2(n933), .ZN(n773) );
  NAND2_X1 U843 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U844 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U845 ( .A(n776), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U847 ( .A(G132), .ZN(G219) );
  INV_X1 U848 ( .A(G82), .ZN(G220) );
  INV_X1 U849 ( .A(G57), .ZN(G237) );
  INV_X1 U850 ( .A(G120), .ZN(G236) );
  INV_X1 U851 ( .A(G69), .ZN(G235) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n777) );
  XNOR2_X1 U853 ( .A(n777), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U854 ( .A(G223), .ZN(n843) );
  NAND2_X1 U855 ( .A1(n843), .A2(G567), .ZN(n778) );
  XOR2_X1 U856 ( .A(KEYINPUT11), .B(n778), .Z(G234) );
  INV_X1 U857 ( .A(G860), .ZN(n803) );
  OR2_X1 U858 ( .A1(n984), .A2(n803), .ZN(G153) );
  INV_X1 U859 ( .A(G171), .ZN(G301) );
  NAND2_X1 U860 ( .A1(G868), .A2(G301), .ZN(n780) );
  INV_X1 U861 ( .A(n987), .ZN(n785) );
  INV_X1 U862 ( .A(G868), .ZN(n825) );
  NAND2_X1 U863 ( .A1(n785), .A2(n825), .ZN(n779) );
  NAND2_X1 U864 ( .A1(n780), .A2(n779), .ZN(G284) );
  NOR2_X1 U865 ( .A1(G286), .A2(n825), .ZN(n782) );
  NOR2_X1 U866 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U867 ( .A1(n782), .A2(n781), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n803), .A2(G559), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n783), .A2(n987), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U871 ( .A1(n785), .A2(n825), .ZN(n786) );
  XOR2_X1 U872 ( .A(KEYINPUT82), .B(n786), .Z(n787) );
  NOR2_X1 U873 ( .A1(G559), .A2(n787), .ZN(n788) );
  XOR2_X1 U874 ( .A(KEYINPUT83), .B(n788), .Z(n791) );
  NOR2_X1 U875 ( .A1(G868), .A2(n984), .ZN(n789) );
  XOR2_X1 U876 ( .A(KEYINPUT81), .B(n789), .Z(n790) );
  NOR2_X1 U877 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U878 ( .A1(G111), .A2(n891), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G99), .A2(n703), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U881 ( .A(KEYINPUT84), .B(n794), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G123), .A2(n707), .ZN(n795) );
  XNOR2_X1 U883 ( .A(n795), .B(KEYINPUT18), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n888), .A2(G135), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n943) );
  XNOR2_X1 U887 ( .A(G2096), .B(n943), .ZN(n801) );
  INV_X1 U888 ( .A(G2100), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(G156) );
  NAND2_X1 U890 ( .A1(G559), .A2(n987), .ZN(n802) );
  XOR2_X1 U891 ( .A(n984), .B(n802), .Z(n822) );
  NAND2_X1 U892 ( .A1(n803), .A2(n822), .ZN(n814) );
  NAND2_X1 U893 ( .A1(n804), .A2(G55), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G67), .A2(n805), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n813) );
  NAND2_X1 U896 ( .A1(G93), .A2(n808), .ZN(n811) );
  NAND2_X1 U897 ( .A1(G80), .A2(n809), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U899 ( .A1(n813), .A2(n812), .ZN(n824) );
  XOR2_X1 U900 ( .A(n814), .B(n824), .Z(G145) );
  XNOR2_X1 U901 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n816) );
  XNOR2_X1 U902 ( .A(G290), .B(KEYINPUT86), .ZN(n815) );
  XNOR2_X1 U903 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U904 ( .A(n824), .B(n817), .ZN(n819) );
  XNOR2_X1 U905 ( .A(G305), .B(G166), .ZN(n818) );
  XNOR2_X1 U906 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U907 ( .A(n820), .B(G288), .ZN(n821) );
  XNOR2_X1 U908 ( .A(n821), .B(G299), .ZN(n911) );
  XOR2_X1 U909 ( .A(n911), .B(n822), .Z(n823) );
  NOR2_X1 U910 ( .A1(n825), .A2(n823), .ZN(n827) );
  AND2_X1 U911 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U912 ( .A1(n827), .A2(n826), .ZN(G295) );
  NAND2_X1 U913 ( .A1(G2078), .A2(G2084), .ZN(n828) );
  XOR2_X1 U914 ( .A(KEYINPUT20), .B(n828), .Z(n829) );
  NAND2_X1 U915 ( .A1(G2090), .A2(n829), .ZN(n830) );
  XNOR2_X1 U916 ( .A(KEYINPUT21), .B(n830), .ZN(n831) );
  NAND2_X1 U917 ( .A1(n831), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U918 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U919 ( .A1(G235), .A2(G236), .ZN(n832) );
  NAND2_X1 U920 ( .A1(G108), .A2(n832), .ZN(n833) );
  NOR2_X1 U921 ( .A1(n833), .A2(G237), .ZN(n834) );
  XNOR2_X1 U922 ( .A(n834), .B(KEYINPUT89), .ZN(n849) );
  AND2_X1 U923 ( .A1(G567), .A2(n849), .ZN(n840) );
  NOR2_X1 U924 ( .A1(G220), .A2(G219), .ZN(n835) );
  XOR2_X1 U925 ( .A(KEYINPUT22), .B(n835), .Z(n836) );
  NOR2_X1 U926 ( .A1(G218), .A2(n836), .ZN(n837) );
  NAND2_X1 U927 ( .A1(G96), .A2(n837), .ZN(n850) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n850), .ZN(n838) );
  XOR2_X1 U929 ( .A(KEYINPUT88), .B(n838), .Z(n839) );
  NOR2_X1 U930 ( .A1(n840), .A2(n839), .ZN(G319) );
  INV_X1 U931 ( .A(G319), .ZN(n842) );
  NAND2_X1 U932 ( .A1(G661), .A2(G483), .ZN(n841) );
  NOR2_X1 U933 ( .A1(n842), .A2(n841), .ZN(n848) );
  NAND2_X1 U934 ( .A1(n848), .A2(G36), .ZN(G176) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n843), .ZN(G217) );
  NAND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n844) );
  XOR2_X1 U937 ( .A(KEYINPUT110), .B(n844), .Z(n845) );
  NAND2_X1 U938 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n846) );
  XOR2_X1 U940 ( .A(KEYINPUT111), .B(n846), .Z(n847) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(G188) );
  XNOR2_X1 U942 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  NOR2_X1 U945 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n851), .B(KEYINPUT112), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2090), .Z(n853) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U951 ( .A(n854), .B(G2096), .Z(n856) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U954 ( .A(KEYINPUT43), .B(G2678), .Z(n858) );
  XNOR2_X1 U955 ( .A(KEYINPUT113), .B(G2100), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n860), .B(n859), .Z(G227) );
  XOR2_X1 U958 ( .A(KEYINPUT115), .B(G1956), .Z(n862) );
  XNOR2_X1 U959 ( .A(G1981), .B(G1961), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(n863), .B(KEYINPUT41), .Z(n865) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U964 ( .A(G1966), .B(G1971), .Z(n867) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1976), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U968 ( .A(KEYINPUT114), .B(G2474), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U970 ( .A1(G136), .A2(n888), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G112), .A2(n891), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G124), .A2(n707), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n703), .A2(G100), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G142), .A2(n888), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G106), .A2(n703), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n881), .B(KEYINPUT45), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G130), .A2(n707), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n891), .A2(G118), .ZN(n884) );
  XOR2_X1 U985 ( .A(KEYINPUT116), .B(n884), .Z(n885) );
  NOR2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n943), .B(n887), .ZN(n900) );
  NAND2_X1 U988 ( .A1(G139), .A2(n888), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G103), .A2(n703), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U991 ( .A1(n891), .A2(G115), .ZN(n892) );
  XOR2_X1 U992 ( .A(KEYINPUT117), .B(n892), .Z(n894) );
  NAND2_X1 U993 ( .A1(n707), .A2(G127), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n935) );
  XNOR2_X1 U997 ( .A(n898), .B(n935), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n905) );
  XNOR2_X1 U999 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n901), .B(G162), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1002 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G164), .B(G160), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G395) );
  XOR2_X1 U1007 ( .A(n911), .B(G286), .Z(n913) );
  XNOR2_X1 U1008 ( .A(G171), .B(n987), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(n984), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(G397) );
  XNOR2_X1 U1012 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n917), .B(n916), .ZN(n928) );
  XOR2_X1 U1015 ( .A(G2451), .B(G2430), .Z(n919) );
  XNOR2_X1 U1016 ( .A(G2438), .B(G2443), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n925) );
  XOR2_X1 U1018 ( .A(G2435), .B(G2454), .Z(n921) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G1348), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n921), .B(n920), .ZN(n923) );
  XOR2_X1 U1021 ( .A(G2446), .B(G2427), .Z(n922) );
  XNOR2_X1 U1022 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1023 ( .A(n925), .B(n924), .Z(n926) );
  NAND2_X1 U1024 ( .A1(G14), .A2(n926), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n931), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(n931), .ZN(G401) );
  INV_X1 U1031 ( .A(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1033 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1036 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n954) );
  XOR2_X1 U1038 ( .A(G2084), .B(G160), .Z(n941) );
  XNOR2_X1 U1039 ( .A(KEYINPUT120), .B(n941), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n950) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(KEYINPUT51), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n955), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT121), .B(n956), .ZN(n957) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n979) );
  NAND2_X1 U1051 ( .A1(n957), .A2(n979), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n958), .A2(G29), .ZN(n1037) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(KEYINPUT125), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(G34), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G2084), .B(n960), .ZN(n977) );
  XNOR2_X1 U1056 ( .A(G2090), .B(G35), .ZN(n975) );
  XOR2_X1 U1057 ( .A(G1991), .B(G25), .Z(n961) );
  NAND2_X1 U1058 ( .A1(n961), .A2(G28), .ZN(n972) );
  XNOR2_X1 U1059 ( .A(G27), .B(KEYINPUT123), .ZN(n963) );
  XNOR2_X1 U1060 ( .A(n963), .B(n962), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(G32), .B(G1996), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(KEYINPUT124), .B(n966), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G2067), .B(G26), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(G33), .B(G2072), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(KEYINPUT53), .B(n973), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n979), .B(n978), .ZN(n981) );
  INV_X1 U1073 ( .A(G29), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(G11), .A2(n982), .ZN(n1035) );
  INV_X1 U1076 ( .A(G16), .ZN(n1031) );
  XOR2_X1 U1077 ( .A(KEYINPUT56), .B(KEYINPUT126), .Z(n983) );
  XNOR2_X1 U1078 ( .A(n1031), .B(n983), .ZN(n1007) );
  XOR2_X1 U1079 ( .A(G1341), .B(n984), .Z(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(n987), .B(G1348), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(G1961), .B(G171), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(G1971), .A2(G303), .ZN(n988) );
  NAND2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n1005) );
  XNOR2_X1 U1088 ( .A(n996), .B(G1956), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G168), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1092 ( .A(KEYINPUT57), .B(n1001), .Z(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1033) );
  XNOR2_X1 U1096 ( .A(G20), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1981), .B(G6), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G19), .B(G1341), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(KEYINPUT59), .B(G1348), .Z(n1013) );
  XNOR2_X1 U1102 ( .A(G4), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1016), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G21), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G1961), .B(G5), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1028) );
  XNOR2_X1 U1109 ( .A(G1986), .B(G24), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G22), .B(G1971), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(G1976), .B(KEYINPUT127), .ZN(n1023) );
  XNOR2_X1 U1113 ( .A(n1023), .B(G23), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1115 ( .A(KEYINPUT58), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1038), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

