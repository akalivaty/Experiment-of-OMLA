

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U559 ( .A1(n540), .A2(n539), .ZN(G160) );
  NOR2_X1 U560 ( .A1(n547), .A2(n546), .ZN(G164) );
  BUF_X1 U561 ( .A(n558), .Z(n559) );
  XNOR2_X1 U562 ( .A(G2104), .B(KEYINPUT64), .ZN(n527) );
  NAND2_X2 U563 ( .A1(n693), .A2(n764), .ZN(n698) );
  XOR2_X1 U564 ( .A(KEYINPUT31), .B(n731), .Z(n523) );
  AND2_X1 U565 ( .A1(n979), .A2(n759), .ZN(n524) );
  XOR2_X1 U566 ( .A(n727), .B(KEYINPUT30), .Z(n525) );
  INV_X1 U567 ( .A(n698), .ZN(n720) );
  INV_X1 U568 ( .A(KEYINPUT29), .ZN(n718) );
  XNOR2_X1 U569 ( .A(n719), .B(n718), .ZN(n724) );
  NOR2_X1 U570 ( .A1(G1966), .A2(n810), .ZN(n725) );
  AND2_X1 U571 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U572 ( .A1(G8), .A2(n698), .ZN(n810) );
  INV_X1 U573 ( .A(G2105), .ZN(n526) );
  AND2_X1 U574 ( .A1(n754), .A2(n524), .ZN(n755) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U576 ( .A(n528), .B(KEYINPUT65), .ZN(n558) );
  INV_X1 U577 ( .A(KEYINPUT23), .ZN(n529) );
  NOR2_X1 U578 ( .A1(n757), .A2(n756), .ZN(n802) );
  NOR2_X1 U579 ( .A1(G651), .A2(n639), .ZN(n661) );
  XNOR2_X1 U580 ( .A(n530), .B(n529), .ZN(n533) );
  XNOR2_X1 U581 ( .A(KEYINPUT66), .B(n534), .ZN(n540) );
  NAND2_X1 U582 ( .A1(n558), .A2(G101), .ZN(n530) );
  XOR2_X1 U583 ( .A(G2104), .B(KEYINPUT64), .Z(n531) );
  AND2_X1 U584 ( .A1(G2105), .A2(n531), .ZN(n889) );
  NAND2_X1 U585 ( .A1(n889), .A2(G125), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  AND2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U588 ( .A1(G113), .A2(n888), .ZN(n538) );
  XNOR2_X1 U589 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n536) );
  NOR2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n535) );
  XNOR2_X1 U591 ( .A(n536), .B(n535), .ZN(n892) );
  NAND2_X1 U592 ( .A1(G137), .A2(n892), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U594 ( .A1(G114), .A2(n888), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G126), .A2(n889), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n558), .A2(G102), .ZN(n543) );
  XOR2_X1 U598 ( .A(KEYINPUT89), .B(n543), .Z(n545) );
  NAND2_X1 U599 ( .A1(n892), .A2(G138), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  NAND2_X1 U602 ( .A1(n661), .A2(G52), .ZN(n550) );
  XOR2_X1 U603 ( .A(G651), .B(KEYINPUT68), .Z(n551) );
  NOR2_X1 U604 ( .A1(G543), .A2(n551), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n548), .Z(n660) );
  NAND2_X1 U606 ( .A1(G64), .A2(n660), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n556) );
  NOR2_X1 U608 ( .A1(G651), .A2(G543), .ZN(n655) );
  NAND2_X1 U609 ( .A1(n655), .A2(G90), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n639), .A2(n551), .ZN(n656) );
  NAND2_X1 U611 ( .A1(G77), .A2(n656), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U616 ( .A1(G123), .A2(n889), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n557), .B(KEYINPUT18), .ZN(n566) );
  NAND2_X1 U618 ( .A1(G135), .A2(n892), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G99), .A2(n559), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n888), .A2(G111), .ZN(n562) );
  XOR2_X1 U622 ( .A(KEYINPUT80), .B(n562), .Z(n563) );
  NOR2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n936) );
  XNOR2_X1 U625 ( .A(G2096), .B(n936), .ZN(n567) );
  OR2_X1 U626 ( .A1(G2100), .A2(n567), .ZN(G156) );
  INV_X1 U627 ( .A(G57), .ZN(G237) );
  INV_X1 U628 ( .A(G82), .ZN(G220) );
  NAND2_X1 U629 ( .A1(n655), .A2(G88), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G75), .A2(n656), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n661), .A2(G50), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G62), .A2(n660), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U635 ( .A1(n573), .A2(n572), .ZN(G166) );
  NAND2_X1 U636 ( .A1(n661), .A2(G51), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G63), .A2(n660), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT6), .B(n576), .ZN(n583) );
  NAND2_X1 U640 ( .A1(G89), .A2(n655), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT76), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT4), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G76), .A2(n656), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(n581), .B(KEYINPUT5), .Z(n582) );
  NOR2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT7), .B(n584), .Z(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT77), .B(n585), .Z(G168) );
  XOR2_X1 U649 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U650 ( .A1(G7), .A2(G661), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U652 ( .A(G223), .ZN(n834) );
  NAND2_X1 U653 ( .A1(n834), .A2(G567), .ZN(n587) );
  XOR2_X1 U654 ( .A(KEYINPUT11), .B(n587), .Z(G234) );
  NAND2_X1 U655 ( .A1(G56), .A2(n660), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT14), .B(n588), .ZN(n595) );
  NAND2_X1 U657 ( .A1(G81), .A2(n655), .ZN(n589) );
  XNOR2_X1 U658 ( .A(n589), .B(KEYINPUT12), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n590), .B(KEYINPUT72), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G68), .A2(n656), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U662 ( .A(KEYINPUT13), .B(n593), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n596), .B(KEYINPUT73), .ZN(n598) );
  NAND2_X1 U665 ( .A1(G43), .A2(n661), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n997) );
  INV_X1 U667 ( .A(n997), .ZN(n599) );
  XNOR2_X1 U668 ( .A(G860), .B(KEYINPUT74), .ZN(n621) );
  NAND2_X1 U669 ( .A1(n599), .A2(n621), .ZN(G153) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n609) );
  NAND2_X1 U672 ( .A1(G54), .A2(n661), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G79), .A2(n656), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G66), .A2(n660), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G92), .A2(n655), .ZN(n602) );
  XNOR2_X1 U677 ( .A(KEYINPUT75), .B(n602), .ZN(n603) );
  NOR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT15), .ZN(n906) );
  INV_X1 U681 ( .A(n906), .ZN(n992) );
  INV_X1 U682 ( .A(G868), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n992), .A2(n617), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(G284) );
  NAND2_X1 U685 ( .A1(n655), .A2(G91), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G78), .A2(n656), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U688 ( .A(KEYINPUT70), .B(n612), .Z(n616) );
  NAND2_X1 U689 ( .A1(n660), .A2(G65), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n661), .A2(G53), .ZN(n613) );
  AND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(G299) );
  NOR2_X1 U693 ( .A1(G286), .A2(n617), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT78), .ZN(n620) );
  NOR2_X1 U695 ( .A1(G299), .A2(G868), .ZN(n619) );
  NOR2_X1 U696 ( .A1(n620), .A2(n619), .ZN(G297) );
  INV_X1 U697 ( .A(G559), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U699 ( .A1(n992), .A2(n623), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT16), .B(n624), .Z(G148) );
  NOR2_X1 U701 ( .A1(G868), .A2(n997), .ZN(n625) );
  XOR2_X1 U702 ( .A(KEYINPUT79), .B(n625), .Z(n628) );
  NAND2_X1 U703 ( .A1(G868), .A2(n906), .ZN(n626) );
  NOR2_X1 U704 ( .A1(G559), .A2(n626), .ZN(n627) );
  NOR2_X1 U705 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U706 ( .A1(n661), .A2(G55), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G67), .A2(n660), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n655), .A2(G93), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G80), .A2(n656), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n669) );
  NAND2_X1 U713 ( .A1(n906), .A2(G559), .ZN(n675) );
  XNOR2_X1 U714 ( .A(n997), .B(n675), .ZN(n635) );
  NOR2_X1 U715 ( .A1(G860), .A2(n635), .ZN(n637) );
  XNOR2_X1 U716 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n636) );
  XNOR2_X1 U717 ( .A(n637), .B(n636), .ZN(n638) );
  XOR2_X1 U718 ( .A(n669), .B(n638), .Z(G145) );
  NAND2_X1 U719 ( .A1(G87), .A2(n639), .ZN(n640) );
  XNOR2_X1 U720 ( .A(n640), .B(KEYINPUT84), .ZN(n643) );
  NAND2_X1 U721 ( .A1(G49), .A2(n661), .ZN(n641) );
  XOR2_X1 U722 ( .A(KEYINPUT83), .B(n641), .Z(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U724 ( .A1(n660), .A2(n644), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G651), .A2(G74), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G86), .A2(n655), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G48), .A2(n661), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n656), .A2(G73), .ZN(n649) );
  XNOR2_X1 U731 ( .A(n649), .B(KEYINPUT2), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n650), .B(KEYINPUT85), .ZN(n651) );
  NOR2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U734 ( .A1(G61), .A2(n660), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U736 ( .A1(n655), .A2(G85), .ZN(n658) );
  NAND2_X1 U737 ( .A1(G72), .A2(n656), .ZN(n657) );
  NAND2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U739 ( .A(KEYINPUT69), .B(n659), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n660), .A2(G60), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n661), .A2(G47), .ZN(n662) );
  AND2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(G290) );
  NOR2_X1 U744 ( .A1(G868), .A2(n669), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT87), .ZN(n678) );
  XOR2_X1 U746 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n667) );
  XNOR2_X1 U747 ( .A(G288), .B(n667), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(G305), .ZN(n672) );
  XNOR2_X1 U749 ( .A(G166), .B(n669), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n670), .B(G299), .ZN(n671) );
  XNOR2_X1 U751 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U752 ( .A(n673), .B(G290), .ZN(n674) );
  XNOR2_X1 U753 ( .A(n674), .B(n997), .ZN(n905) );
  XNOR2_X1 U754 ( .A(n905), .B(n675), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G868), .A2(n676), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n679) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U763 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U766 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U767 ( .A1(G96), .A2(n685), .ZN(n838) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n838), .ZN(n689) );
  NAND2_X1 U769 ( .A1(G108), .A2(G120), .ZN(n686) );
  NOR2_X1 U770 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G69), .A2(n687), .ZN(n839) );
  NAND2_X1 U772 ( .A1(G567), .A2(n839), .ZN(n688) );
  NAND2_X1 U773 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U774 ( .A(KEYINPUT88), .B(n690), .Z(G319) );
  INV_X1 U775 ( .A(G319), .ZN(n692) );
  NAND2_X1 U776 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n837) );
  NAND2_X1 U778 ( .A1(n837), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G166), .ZN(G303) );
  NAND2_X1 U780 ( .A1(G160), .A2(G40), .ZN(n765) );
  INV_X1 U781 ( .A(n765), .ZN(n693) );
  NOR2_X1 U782 ( .A1(G164), .A2(G1384), .ZN(n764) );
  NAND2_X1 U783 ( .A1(n720), .A2(G2067), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G1348), .A2(n698), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U786 ( .A(n696), .B(KEYINPUT100), .Z(n704) );
  OR2_X1 U787 ( .A1(n906), .A2(n704), .ZN(n703) );
  INV_X1 U788 ( .A(G1996), .ZN(n953) );
  NOR2_X1 U789 ( .A1(n698), .A2(n953), .ZN(n697) );
  XOR2_X1 U790 ( .A(n697), .B(KEYINPUT26), .Z(n700) );
  NAND2_X1 U791 ( .A1(n698), .A2(G1341), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U793 ( .A1(n997), .A2(n701), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U795 ( .A1(n704), .A2(n906), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U797 ( .A(n707), .B(KEYINPUT101), .ZN(n712) );
  NAND2_X1 U798 ( .A1(n720), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U799 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  AND2_X1 U800 ( .A1(G1956), .A2(n698), .ZN(n709) );
  NOR2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n714) );
  INV_X1 U802 ( .A(G299), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U806 ( .A(n715), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U808 ( .A(G1961), .B(KEYINPUT99), .ZN(n1024) );
  NAND2_X1 U809 ( .A1(n698), .A2(n1024), .ZN(n722) );
  XNOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U811 ( .A1(n720), .A2(n955), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n728) );
  NAND2_X1 U813 ( .A1(n728), .A2(G171), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n732) );
  XOR2_X1 U815 ( .A(KEYINPUT98), .B(n725), .Z(n743) );
  INV_X1 U816 ( .A(G8), .ZN(n738) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n698), .ZN(n742) );
  NOR2_X1 U818 ( .A1(n738), .A2(n742), .ZN(n726) );
  AND2_X1 U819 ( .A1(n743), .A2(n726), .ZN(n727) );
  NOR2_X1 U820 ( .A1(G168), .A2(n525), .ZN(n730) );
  NOR2_X1 U821 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U823 ( .A1(n732), .A2(n523), .ZN(n744) );
  AND2_X1 U824 ( .A1(G286), .A2(G8), .ZN(n733) );
  NAND2_X1 U825 ( .A1(n744), .A2(n733), .ZN(n740) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n810), .ZN(n735) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n698), .ZN(n734) );
  NOR2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U831 ( .A(n741), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U832 ( .A1(G8), .A2(n742), .ZN(n746) );
  AND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U834 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U836 ( .A(n749), .B(KEYINPUT102), .ZN(n808) );
  INV_X1 U837 ( .A(n808), .ZN(n752) );
  INV_X1 U838 ( .A(G1971), .ZN(n1016) );
  NAND2_X1 U839 ( .A1(G166), .A2(n1016), .ZN(n751) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n760) );
  INV_X1 U841 ( .A(n760), .ZN(n750) );
  NAND2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n981) );
  NOR2_X1 U843 ( .A1(n752), .A2(n981), .ZN(n753) );
  NOR2_X1 U844 ( .A1(n810), .A2(n753), .ZN(n754) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NOR2_X1 U846 ( .A1(n755), .A2(KEYINPUT33), .ZN(n757) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n989) );
  INV_X1 U848 ( .A(n989), .ZN(n756) );
  INV_X1 U849 ( .A(KEYINPUT103), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n760), .A2(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n759), .A2(n758), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n760), .A2(KEYINPUT103), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U854 ( .A1(n810), .A2(n763), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n766), .B(KEYINPUT90), .ZN(n827) );
  XNOR2_X1 U857 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U858 ( .A1(n827), .A2(n987), .ZN(n767) );
  XOR2_X1 U859 ( .A(n767), .B(KEYINPUT91), .Z(n804) );
  AND2_X1 U860 ( .A1(n768), .A2(n804), .ZN(n800) );
  NAND2_X1 U861 ( .A1(n559), .A2(G95), .ZN(n769) );
  XOR2_X1 U862 ( .A(KEYINPUT93), .B(n769), .Z(n771) );
  NAND2_X1 U863 ( .A1(n892), .A2(G131), .ZN(n770) );
  NAND2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U865 ( .A(KEYINPUT94), .B(n772), .Z(n776) );
  NAND2_X1 U866 ( .A1(G107), .A2(n888), .ZN(n774) );
  NAND2_X1 U867 ( .A1(G119), .A2(n889), .ZN(n773) );
  AND2_X1 U868 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n887) );
  NAND2_X1 U870 ( .A1(G1991), .A2(n887), .ZN(n777) );
  XNOR2_X1 U871 ( .A(n777), .B(KEYINPUT95), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n892), .A2(G141), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n559), .A2(G105), .ZN(n778) );
  XNOR2_X1 U874 ( .A(n778), .B(KEYINPUT38), .ZN(n780) );
  NAND2_X1 U875 ( .A1(G117), .A2(n888), .ZN(n779) );
  NAND2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U877 ( .A1(n889), .A2(G129), .ZN(n781) );
  XOR2_X1 U878 ( .A(KEYINPUT96), .B(n781), .Z(n782) );
  NOR2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U880 ( .A(KEYINPUT97), .B(n784), .Z(n785) );
  NAND2_X1 U881 ( .A1(n786), .A2(n785), .ZN(n882) );
  AND2_X1 U882 ( .A1(G1996), .A2(n882), .ZN(n787) );
  NOR2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n818) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NAND2_X1 U885 ( .A1(n888), .A2(G116), .ZN(n789) );
  XNOR2_X1 U886 ( .A(n789), .B(KEYINPUT92), .ZN(n791) );
  NAND2_X1 U887 ( .A1(G128), .A2(n889), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U889 ( .A(n792), .B(KEYINPUT35), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G140), .A2(n892), .ZN(n794) );
  NAND2_X1 U891 ( .A1(G104), .A2(n559), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U893 ( .A(KEYINPUT34), .B(n795), .Z(n796) );
  NAND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U895 ( .A(n798), .B(KEYINPUT36), .Z(n901) );
  OR2_X1 U896 ( .A1(n825), .A2(n901), .ZN(n941) );
  NAND2_X1 U897 ( .A1(n818), .A2(n941), .ZN(n799) );
  NAND2_X1 U898 ( .A1(n799), .A2(n827), .ZN(n803) );
  AND2_X1 U899 ( .A1(n800), .A2(n803), .ZN(n801) );
  NAND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n832) );
  INV_X1 U901 ( .A(n803), .ZN(n817) );
  INV_X1 U902 ( .A(n804), .ZN(n815) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n805) );
  XOR2_X1 U904 ( .A(n805), .B(KEYINPUT24), .Z(n806) );
  OR2_X1 U905 ( .A1(n810), .A2(n806), .ZN(n813) );
  NOR2_X1 U906 ( .A1(G2090), .A2(G303), .ZN(n807) );
  NAND2_X1 U907 ( .A1(G8), .A2(n807), .ZN(n809) );
  NAND2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n830) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n882), .ZN(n927) );
  INV_X1 U914 ( .A(n818), .ZN(n948) );
  NOR2_X1 U915 ( .A1(n887), .A2(G1991), .ZN(n819) );
  XNOR2_X1 U916 ( .A(n819), .B(KEYINPUT104), .ZN(n939) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n939), .A2(n820), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n948), .A2(n821), .ZN(n822) );
  NOR2_X1 U920 ( .A1(n927), .A2(n822), .ZN(n823) );
  XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n823), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n824), .A2(n941), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n825), .A2(n901), .ZN(n934) );
  NAND2_X1 U924 ( .A1(n826), .A2(n934), .ZN(n828) );
  AND2_X1 U925 ( .A1(n828), .A2(n827), .ZN(n829) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U931 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G188) );
  XOR2_X1 U934 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  INV_X1 U936 ( .A(G108), .ZN(G238) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(G2100), .B(G2096), .Z(n841) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(G2678), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2072), .Z(n843) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2090), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U946 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1976), .B(G1961), .Z(n849) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1966), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U952 ( .A(G1971), .B(G1956), .Z(n851) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U956 ( .A(G2474), .B(KEYINPUT107), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n857) );
  XOR2_X1 U958 ( .A(G1981), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G124), .A2(n889), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n858), .B(KEYINPUT44), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n859), .B(KEYINPUT108), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G112), .A2(n888), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G136), .A2(n892), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G100), .A2(n559), .ZN(n862) );
  NAND2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U968 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G139), .A2(n892), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G103), .A2(n559), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G115), .A2(n888), .ZN(n869) );
  NAND2_X1 U973 ( .A1(G127), .A2(n889), .ZN(n868) );
  NAND2_X1 U974 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U975 ( .A(KEYINPUT112), .B(n870), .Z(n871) );
  XNOR2_X1 U976 ( .A(KEYINPUT47), .B(n871), .ZN(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n930) );
  XOR2_X1 U978 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n875) );
  XNOR2_X1 U979 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n874) );
  XNOR2_X1 U980 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U981 ( .A(n876), .B(KEYINPUT111), .Z(n878) );
  XNOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n877) );
  XNOR2_X1 U983 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U984 ( .A(n930), .B(n879), .Z(n880) );
  XNOR2_X1 U985 ( .A(n936), .B(n880), .ZN(n881) );
  XOR2_X1 U986 ( .A(n881), .B(G162), .Z(n884) );
  XOR2_X1 U987 ( .A(G164), .B(n882), .Z(n883) );
  XNOR2_X1 U988 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U989 ( .A(G160), .B(n885), .Z(n886) );
  XNOR2_X1 U990 ( .A(n887), .B(n886), .ZN(n903) );
  NAND2_X1 U991 ( .A1(G118), .A2(n888), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G130), .A2(n889), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n899) );
  XNOR2_X1 U994 ( .A(KEYINPUT110), .B(KEYINPUT45), .ZN(n897) );
  NAND2_X1 U995 ( .A1(n892), .A2(G142), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n559), .A2(G106), .ZN(n893) );
  XOR2_X1 U997 ( .A(KEYINPUT109), .B(n893), .Z(n894) );
  NAND2_X1 U998 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U999 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n904), .ZN(G395) );
  XOR2_X1 U1004 ( .A(n905), .B(G286), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G171), .B(n906), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1008 ( .A(G2454), .B(G2435), .Z(n911) );
  XNOR2_X1 U1009 ( .A(G2438), .B(G2427), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(n918) );
  XOR2_X1 U1011 ( .A(KEYINPUT105), .B(G2446), .Z(n913) );
  XNOR2_X1 U1012 ( .A(G2443), .B(G2430), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1014 ( .A(n914), .B(G2451), .Z(n916) );
  XNOR2_X1 U1015 ( .A(G1341), .B(G1348), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n918), .B(n917), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n919), .A2(G14), .ZN(n925) );
  NAND2_X1 U1019 ( .A1(n925), .A2(G319), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G69), .ZN(G235) );
  INV_X1 U1027 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1030 ( .A(KEYINPUT118), .B(n928), .Z(n929) );
  XNOR2_X1 U1031 ( .A(KEYINPUT51), .B(n929), .ZN(n946) );
  XOR2_X1 U1032 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1033 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(n933), .B(KEYINPUT50), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G160), .B(G2084), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT117), .B(n942), .Z(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1045 ( .A(KEYINPUT119), .B(n949), .Z(n950) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n950), .ZN(n951) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n974) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n974), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n952), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G35), .ZN(n968) );
  XNOR2_X1 U1051 ( .A(G32), .B(n953), .ZN(n960) );
  XOR2_X1 U1052 ( .A(G1991), .B(G25), .Z(n954) );
  NAND2_X1 U1053 ( .A1(n954), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G27), .B(n955), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(KEYINPUT121), .B(n956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(G2072), .B(G33), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1061 ( .A(KEYINPUT120), .B(n963), .Z(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n966), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(n969), .B(KEYINPUT122), .ZN(n972) );
  XOR2_X1 U1066 ( .A(G2084), .B(G34), .Z(n970) );
  XNOR2_X1 U1067 ( .A(KEYINPUT54), .B(n970), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(n974), .B(n973), .ZN(n976) );
  INV_X1 U1070 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(G11), .A2(n977), .ZN(n1033) );
  XNOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .ZN(n1003) );
  XNOR2_X1 U1074 ( .A(G299), .B(G1956), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(G1971), .A2(G303), .ZN(n978) );
  NAND2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(KEYINPUT123), .B(n982), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1080 ( .A(KEYINPUT124), .B(n985), .Z(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1082 ( .A(KEYINPUT125), .B(n988), .Z(n1001) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G168), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n991), .B(KEYINPUT57), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G301), .B(G1961), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(n992), .B(G1348), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(G1341), .B(n997), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1031) );
  INV_X1 U1094 ( .A(G16), .ZN(n1029) );
  XNOR2_X1 U1095 ( .A(G1348), .B(KEYINPUT59), .ZN(n1004) );
  XNOR2_X1 U1096 ( .A(n1004), .B(G4), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1005) );
  NOR2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(KEYINPUT126), .B(G1956), .ZN(n1009) );
  XNOR2_X1 U1102 ( .A(G20), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G21), .ZN(n1013) );
  NOR2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1107 ( .A(KEYINPUT127), .B(n1015), .Z(n1023) );
  XOR2_X1 U1108 ( .A(G1986), .B(G24), .Z(n1018) );
  XNOR2_X1 U1109 ( .A(n1016), .B(G22), .ZN(n1017) );
  NAND2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1111 ( .A(G23), .B(G1976), .ZN(n1019) );
  NOR2_X1 U1112 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1113 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1114 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XOR2_X1 U1115 ( .A(G5), .B(n1024), .Z(n1025) );
  NOR2_X1 U1116 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

