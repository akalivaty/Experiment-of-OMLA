//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  OR4_X1    g028(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT69), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT70), .ZN(G160));
  NAND2_X1  g052(.A1(new_n469), .A2(new_n471), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT71), .B1(new_n478), .B2(new_n462), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n463), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n478), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n482), .A2(G124), .B1(G136), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT72), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n478), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n468), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G102), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n469), .A2(new_n471), .A3(G138), .A4(new_n462), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n493), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n504), .B(new_n506), .C1(new_n512), .C2(new_n513), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n511), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(new_n518), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n514), .A2(new_n525), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n523), .B1(new_n527), .B2(G51), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G168));
  AND2_X1   g107(.A1(new_n527), .A2(G52), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT75), .B(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n534), .A2(new_n502), .B1(new_n518), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(new_n527), .A2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n507), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n518), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT76), .B(G81), .Z(new_n543));
  AOI22_X1  g118(.A1(G651), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT77), .B1(new_n515), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n514), .A2(new_n555), .A3(G53), .A4(G543), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT77), .B(new_n559), .C1(new_n515), .C2(new_n553), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n542), .A2(G91), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n561), .C1(new_n502), .C2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  NAND2_X1  g141(.A1(new_n528), .A2(new_n531), .ZN(G286));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  NAND2_X1  g143(.A1(G166), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT78), .B1(new_n511), .B2(new_n519), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G303));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n502), .B1(new_n507), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(G87), .B2(new_n542), .ZN(new_n574));
  OAI211_X1 g149(.A(G49), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n507), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT80), .ZN(new_n583));
  OAI211_X1 g158(.A(G48), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n518), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n581), .A2(new_n588), .A3(G651), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n583), .A2(new_n587), .A3(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n527), .A2(G47), .B1(G85), .B2(new_n542), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT81), .B1(new_n592), .B2(new_n502), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n592), .A2(KEYINPUT81), .A3(new_n502), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(new_n527), .A2(G54), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n518), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G79), .ZN(new_n600));
  OR3_X1    g175(.A1(new_n600), .A2(new_n503), .A3(KEYINPUT82), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT82), .B1(new_n600), .B2(new_n503), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n603), .C2(new_n507), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n596), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n564), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(G868), .B2(new_n564), .ZN(G280));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n545), .A2(new_n607), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n606), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n482), .A2(G123), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n468), .B1(new_n625), .B2(G2105), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n483), .A2(G135), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n463), .A2(new_n494), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  AND2_X1   g208(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n629), .B(new_n636), .C1(new_n634), .C2(new_n632), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  AND2_X1   g225(.A1(new_n650), .A2(G14), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n652), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(new_n633), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n654), .A2(new_n655), .ZN(new_n661));
  AOI21_X1  g236(.A(KEYINPUT18), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT87), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n674), .A2(new_n665), .A3(new_n668), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n672), .B(new_n675), .C1(new_n665), .C2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G1981), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n684), .A2(G6), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G305), .B2(G16), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n686), .A2(new_n687), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(new_n689), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n684), .A2(G23), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G288), .B2(G16), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(KEYINPUT89), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n701));
  AOI211_X1 g276(.A(new_n701), .B(new_n696), .C1(G288), .C2(G16), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n699), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n684), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n684), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n700), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n698), .B2(new_n702), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n704), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT34), .B1(new_n695), .B2(new_n711), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n704), .A2(new_n710), .A3(new_n708), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT34), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n713), .A2(new_n714), .A3(new_n694), .A4(new_n691), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n482), .A2(G119), .B1(G131), .B2(new_n483), .ZN(new_n721));
  OR2_X1    g296(.A1(G95), .A2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n722), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n720), .B1(new_n725), .B2(new_n719), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT35), .B(G1991), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(G16), .A2(G24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G290), .B2(new_n684), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n717), .A2(new_n718), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n712), .A2(new_n715), .A3(new_n716), .A4(new_n729), .ZN(new_n734));
  INV_X1    g309(.A(new_n732), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT36), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT101), .B1(new_n628), .B2(new_n719), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT101), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n623), .A2(new_n739), .A3(G29), .A4(new_n627), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G5), .A2(G16), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G171), .B2(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G1961), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n719), .B1(new_n745), .B2(G28), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT102), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n745), .A2(G28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n741), .A2(new_n744), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT103), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G11), .ZN(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G21), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G168), .B2(G16), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT100), .B(G1966), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n752), .A2(new_n753), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n743), .A2(G1961), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n719), .A2(G35), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n488), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G27), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT104), .B1(new_n766), .B2(G29), .ZN(new_n767));
  OR3_X1    g342(.A1(new_n766), .A2(KEYINPUT104), .A3(G29), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(G164), .C2(new_n719), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2078), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT99), .ZN(new_n772));
  OR2_X1    g347(.A1(G29), .A2(G32), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT97), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n482), .B2(G129), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n483), .A2(G141), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n772), .B(new_n773), .C1(new_n784), .C2(new_n719), .ZN(new_n785));
  AND4_X1   g360(.A1(new_n760), .A2(new_n765), .A3(new_n770), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(G115), .A2(G2104), .ZN(new_n787));
  INV_X1    g362(.A(G127), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n478), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G2105), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT93), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n483), .A2(G139), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n494), .A2(G103), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT25), .Z(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n791), .A2(KEYINPUT94), .A3(new_n792), .A4(new_n794), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n801), .A2(new_n802), .A3(new_n719), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n719), .A2(G33), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(G2072), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G4), .B2(G16), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n807), .A2(G4), .A3(G16), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n808), .B(new_n809), .C1(new_n606), .C2(new_n684), .ZN(new_n810));
  INV_X1    g385(.A(G1348), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n719), .A2(G26), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n482), .A2(G128), .B1(G140), .B2(new_n483), .ZN(new_n816));
  OR2_X1    g391(.A1(G104), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n815), .B1(new_n819), .B2(G29), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n812), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n759), .A2(new_n786), .A3(new_n806), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n741), .A2(new_n754), .A3(new_n744), .A4(new_n751), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n756), .A2(new_n757), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n756), .A2(new_n757), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT103), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G2072), .ZN(new_n830));
  INV_X1    g405(.A(new_n802), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(new_n800), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n830), .B(new_n804), .C1(new_n832), .C2(new_n719), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n763), .A2(new_n764), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT105), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n684), .A2(KEYINPUT23), .A3(G20), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT23), .ZN(new_n837));
  INV_X1    g412(.A(G20), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(G16), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n836), .B(new_n839), .C1(new_n564), .C2(new_n684), .ZN(new_n840));
  INV_X1    g415(.A(G1956), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n834), .A2(new_n835), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n829), .A2(new_n833), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(G160), .A2(G29), .ZN(new_n845));
  AND2_X1   g420(.A1(KEYINPUT24), .A2(G34), .ZN(new_n846));
  NOR2_X1   g421(.A1(KEYINPUT24), .A2(G34), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n719), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G2084), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n684), .A2(G19), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n546), .B2(new_n684), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G1341), .ZN(new_n856));
  NOR4_X1   g431(.A1(new_n824), .A2(new_n844), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n769), .A2(G2078), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n737), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n834), .A2(new_n842), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT105), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n773), .B1(new_n784), .B2(new_n719), .ZN(new_n862));
  INV_X1    g437(.A(new_n772), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n859), .A2(KEYINPUT106), .A3(new_n861), .A4(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n737), .A2(new_n857), .A3(new_n864), .A4(new_n858), .ZN(new_n867));
  INV_X1    g442(.A(new_n861), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n869), .ZN(G311));
  NAND3_X1  g445(.A1(new_n859), .A2(new_n861), .A3(new_n864), .ZN(G150));
  NAND2_X1  g446(.A1(new_n542), .A2(G93), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(new_n502), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n527), .B2(G55), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT107), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n545), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n875), .A2(new_n545), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n614), .A2(G559), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT38), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n883), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n879), .B1(new_n886), .B2(G860), .ZN(G145));
  XNOR2_X1  g462(.A(new_n488), .B(KEYINPUT108), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(G160), .Z(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(new_n628), .Z(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n782), .A2(new_n783), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n492), .A2(G2105), .B1(G102), .B2(new_n494), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n498), .A2(new_n499), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n490), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n463), .B2(G126), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n495), .B1(new_n898), .B2(new_n462), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n498), .A2(new_n499), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT109), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n819), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n782), .B2(new_n783), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n896), .A2(new_n901), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n784), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n819), .B1(new_n909), .B2(new_n905), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n832), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n482), .A2(G130), .B1(G142), .B2(new_n483), .ZN(new_n913));
  NOR2_X1   g488(.A1(G106), .A2(G2105), .ZN(new_n914));
  OAI21_X1  g489(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(new_n631), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n724), .ZN(new_n918));
  INV_X1    g493(.A(new_n797), .ZN(new_n919));
  INV_X1    g494(.A(new_n799), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n907), .A2(new_n910), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n912), .A2(KEYINPUT110), .A3(new_n918), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n912), .A2(new_n918), .A3(new_n922), .ZN(new_n924));
  INV_X1    g499(.A(new_n918), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n907), .A2(new_n910), .A3(new_n921), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n911), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n891), .B(new_n923), .C1(new_n928), .C2(KEYINPUT110), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n927), .A3(new_n890), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g508(.A1(new_n877), .A2(new_n607), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n564), .A2(new_n606), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT111), .ZN(new_n936));
  NAND2_X1  g511(.A1(G299), .A2(new_n614), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n564), .A2(new_n938), .A3(new_n606), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n936), .A2(new_n939), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT113), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n936), .A2(new_n945), .A3(new_n939), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n937), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n940), .B(KEYINPUT112), .Z(new_n949));
  XNOR2_X1  g524(.A(new_n882), .B(new_n618), .ZN(new_n950));
  MUX2_X1   g525(.A(new_n948), .B(new_n949), .S(new_n950), .Z(new_n951));
  XNOR2_X1  g526(.A(G166), .B(KEYINPUT114), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(G305), .ZN(new_n953));
  INV_X1    g528(.A(G288), .ZN(new_n954));
  XNOR2_X1  g529(.A(G290), .B(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n953), .B(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT42), .Z(new_n957));
  XNOR2_X1  g532(.A(new_n951), .B(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n934), .B1(new_n958), .B2(new_n607), .ZN(G295));
  OAI21_X1  g534(.A(new_n934), .B1(new_n958), .B2(new_n607), .ZN(G331));
  XNOR2_X1  g535(.A(G168), .B(G171), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n882), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n880), .A3(new_n881), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n940), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n948), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n956), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n956), .B(new_n965), .C1(new_n948), .C2(new_n966), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n930), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n971), .A2(new_n930), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(KEYINPUT115), .A3(new_n970), .A4(new_n969), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n966), .A2(new_n949), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n963), .A2(new_n964), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n940), .A2(new_n941), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n978), .B(new_n979), .C1(new_n941), .C2(new_n947), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n980), .A3(new_n968), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n930), .A3(new_n971), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT44), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n970), .B1(new_n975), .B2(new_n969), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n987), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  INV_X1    g564(.A(G40), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n466), .A2(new_n990), .A3(new_n474), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n989), .B(new_n991), .C1(new_n908), .C2(G1384), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n819), .B(new_n821), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n892), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(KEYINPUT126), .B2(new_n995), .ZN(new_n996));
  OR4_X1    g571(.A1(KEYINPUT126), .A2(new_n992), .A3(new_n995), .A4(G1996), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n992), .A2(G1996), .B1(KEYINPUT126), .B2(new_n995), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT47), .ZN(new_n1000));
  INV_X1    g575(.A(new_n992), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G290), .A2(G1986), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT48), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n892), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n784), .A2(G1996), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n993), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n725), .A2(new_n728), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n724), .A2(new_n727), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1004), .B1(new_n1011), .B2(new_n992), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1008), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1013), .A2(new_n1010), .B1(new_n821), .B2(new_n904), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1014), .A2(new_n992), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1000), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT127), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT125), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n562), .A2(new_n502), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(G91), .B2(new_n542), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(KEYINPUT57), .A3(new_n557), .A4(new_n560), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n558), .B2(new_n563), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT50), .B1(new_n500), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT50), .B(new_n1026), .C1(new_n899), .C2(new_n900), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n991), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n841), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT45), .B(new_n1026), .C1(new_n896), .C2(new_n901), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n467), .A2(new_n475), .A3(G40), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1026), .B1(new_n899), .B2(new_n900), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(new_n989), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT56), .B(G2072), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1025), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1031), .A2(new_n1025), .A3(new_n1037), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1030), .A2(new_n811), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n991), .A2(new_n500), .A3(new_n1026), .A4(new_n821), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT123), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1034), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(KEYINPUT123), .A3(new_n821), .A4(new_n991), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1039), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1038), .B1(new_n1048), .B2(new_n614), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1032), .A2(new_n1005), .A3(new_n1035), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT58), .B(G1341), .Z(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n546), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(KEYINPUT59), .A3(new_n546), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1039), .A2(KEYINPUT61), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT61), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1031), .A2(new_n1025), .A3(new_n1037), .A4(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT60), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1034), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1028), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1348), .B1(new_n1066), .B2(new_n991), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1040), .A2(KEYINPUT60), .A3(new_n1046), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n614), .A3(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1040), .A2(KEYINPUT60), .A3(new_n606), .A4(new_n1046), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1049), .B1(new_n1061), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G286), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  INV_X1    g650(.A(G8), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n528), .B2(new_n531), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1075), .B1(new_n1077), .B2(KEYINPUT124), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1033), .B1(new_n1065), .B2(new_n1028), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1034), .A2(new_n989), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT45), .B(new_n1026), .C1(new_n899), .C2(new_n900), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n991), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n852), .A2(new_n1079), .B1(new_n1082), .B2(new_n757), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1074), .B(new_n1078), .C1(new_n1083), .C2(new_n1076), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT51), .B1(new_n1074), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1082), .A2(new_n757), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n852), .B(new_n991), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(G8), .B(new_n1086), .C1(new_n1089), .C2(G286), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(G8), .A3(G286), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1084), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(G2078), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1079), .A2(G1961), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1093), .A2(G2078), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1035), .A2(new_n1081), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G171), .B(KEYINPUT54), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n989), .B1(new_n908), .B2(G1384), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1103), .A2(new_n991), .A3(new_n1032), .A4(new_n1097), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1095), .A2(new_n1104), .A3(new_n1100), .A4(new_n1096), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1092), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1073), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1092), .A2(KEYINPUT62), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1084), .A2(new_n1090), .A3(new_n1091), .A4(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(G171), .A3(new_n1110), .A4(new_n1099), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1089), .A2(G8), .A3(G168), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(KEYINPUT63), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1094), .A2(new_n707), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1079), .A2(new_n764), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1094), .A2(KEYINPUT116), .A3(new_n707), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(G303), .A2(G8), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1122), .A2(KEYINPUT55), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(KEYINPUT55), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(G8), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1116), .A2(new_n1128), .A3(new_n1119), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G8), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1127), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT118), .B(G1981), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n583), .A2(new_n587), .A3(new_n589), .A4(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT119), .ZN(new_n1135));
  NAND2_X1  g710(.A1(G305), .A2(G1981), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT49), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1076), .B1(new_n1044), .B2(new_n991), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(KEYINPUT49), .A3(new_n1136), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n954), .A2(G1976), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT52), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT117), .B1(new_n954), .B2(G1976), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1144), .B(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(KEYINPUT121), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1126), .B(new_n1132), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1115), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1140), .ZN(new_n1155));
  INV_X1    g730(.A(G1976), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1142), .A2(new_n1156), .A3(new_n954), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1157), .B2(new_n1135), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1148), .A2(new_n1127), .B1(KEYINPUT122), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1121), .A2(G8), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(KEYINPUT122), .A3(new_n1127), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1112), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1148), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI221_X4 g741(.A(new_n1158), .B1(new_n1160), .B2(new_n1162), .C1(new_n1166), .C2(KEYINPUT63), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1154), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(G290), .A2(G1986), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1011), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1001), .B1(new_n1170), .B2(new_n1002), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1019), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1113), .B1(new_n1073), .B2(new_n1106), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1152), .B1(new_n1173), .B2(new_n1111), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1158), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1125), .B1(new_n1121), .B2(G8), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1112), .B(new_n1148), .C1(new_n1177), .C2(KEYINPUT122), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1175), .B(new_n1176), .C1(new_n1178), .C2(new_n1159), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1019), .B(new_n1171), .C1(new_n1174), .C2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1018), .B1(new_n1172), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g757(.A(G319), .B(new_n682), .C1(new_n985), .C2(new_n986), .ZN(new_n1184));
  AOI21_X1  g758(.A(G227), .B1(new_n650), .B2(G14), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n932), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n1184), .A2(new_n1186), .ZN(G308));
  INV_X1    g761(.A(new_n969), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n971), .A2(new_n930), .ZN(new_n1189));
  OAI21_X1  g763(.A(KEYINPUT43), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n975), .A2(new_n970), .A3(new_n981), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n460), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g766(.A1(new_n1192), .A2(new_n682), .A3(new_n932), .A4(new_n1185), .ZN(G225));
endmodule


