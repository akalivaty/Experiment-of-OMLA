//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n461), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n465), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n467), .A2(new_n468), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT65), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n479), .A2(new_n461), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n478), .B(new_n482), .C1(G124), .C2(new_n483), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n470), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n480), .A2(KEYINPUT4), .A3(G138), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(G126), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT66), .A3(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(G50), .A3(G543), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n503), .B(KEYINPUT67), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT68), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  AND2_X1   g085(.A1(G75), .A2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n502), .A2(new_n509), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n504), .A2(new_n515), .ZN(G166));
  INV_X1    g091(.A(new_n509), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n501), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G89), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n501), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  AND3_X1   g098(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT5), .B1(KEYINPUT68), .B2(G543), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n507), .A2(KEYINPUT69), .A3(new_n508), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n519), .A2(new_n522), .A3(new_n529), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n499), .A2(new_n509), .A3(G90), .A4(new_n500), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n499), .A2(G52), .A3(G543), .A4(new_n500), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n536), .A3(new_n534), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n526), .A2(new_n527), .A3(G64), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n538), .A2(new_n539), .B1(G651), .B2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(new_n521), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(new_n513), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n528), .A2(G56), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n495), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n521), .A2(G53), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n556), .A2(KEYINPUT71), .A3(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n521), .A2(G53), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n517), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(G91), .A2(new_n518), .B1(new_n563), .B2(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G299));
  NAND2_X1  g140(.A1(new_n542), .A2(G651), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n535), .A2(new_n536), .A3(new_n534), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n567), .B2(new_n537), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT72), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n566), .B(new_n570), .C1(new_n567), .C2(new_n537), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G301));
  INV_X1    g148(.A(G166), .ZN(G303));
  AOI22_X1  g149(.A1(G49), .A2(new_n521), .B1(new_n518), .B2(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n518), .A2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n521), .A2(G48), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n509), .A2(G61), .ZN(new_n580));
  AND2_X1   g155(.A1(G73), .A2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n528), .A2(G60), .ZN(new_n584));
  INV_X1    g159(.A(G72), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n520), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n495), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(new_n587), .B2(new_n586), .ZN(new_n589));
  AOI22_X1  g164(.A1(G47), .A2(new_n521), .B1(new_n518), .B2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(new_n518), .A2(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n517), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(G54), .A2(new_n521), .B1(new_n597), .B2(G651), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(G868), .B2(new_n572), .ZN(G284));
  AOI21_X1  g176(.A(new_n600), .B1(G868), .B2(new_n572), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  XNOR2_X1  g180(.A(G280), .B(KEYINPUT74), .ZN(G297));
  INV_X1    g181(.A(new_n599), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(KEYINPUT75), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(KEYINPUT75), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n612), .B(new_n613), .C1(G868), .C2(new_n550), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n464), .A2(new_n469), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT76), .B(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT77), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n480), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n483), .A2(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n461), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  OAI211_X1 g202(.A(new_n621), .B(new_n627), .C1(new_n619), .C2(new_n618), .ZN(G156));
  XOR2_X1   g203(.A(KEYINPUT15), .B(G2435), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT78), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n630), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(new_n643), .A3(G14), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT79), .ZN(G401));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT17), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n649), .B2(new_n646), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  INV_X1    g230(.A(new_n646), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n656), .A2(new_n652), .A3(new_n648), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n647), .A2(new_n652), .A3(new_n649), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT81), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n665), .A2(new_n666), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(new_n668), .ZN(new_n674));
  MUX2_X1   g249(.A(new_n674), .B(new_n673), .S(new_n664), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(G288), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT33), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1976), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(G22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT85), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n683), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1971), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT32), .B(G1981), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT84), .Z(new_n696));
  AOI21_X1  g271(.A(new_n692), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n688), .B(new_n697), .C1(new_n694), .C2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G24), .B(G290), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT83), .Z(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G1986), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(G1986), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n480), .A2(G131), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n483), .A2(G119), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n461), .A2(G107), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT82), .ZN(new_n710));
  MUX2_X1   g285(.A(G25), .B(new_n710), .S(G29), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n703), .A2(new_n704), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n700), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT36), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G164), .A2(new_n718), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G27), .B2(new_n718), .ZN(new_n725));
  INV_X1    g300(.A(G2078), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G34), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(KEYINPUT24), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n728), .B2(KEYINPUT24), .ZN(new_n730));
  AOI22_X1  g305(.A1(G160), .A2(G29), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G2084), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n718), .A2(G33), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT25), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n469), .A2(G127), .ZN(new_n736));
  NAND2_X1  g311(.A1(G115), .A2(G2104), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n461), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n735), .B(new_n738), .C1(G139), .C2(new_n480), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n718), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G2072), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n727), .A2(new_n732), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n718), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n745), .A2(G104), .A3(G2105), .ZN(new_n746));
  INV_X1    g321(.A(G104), .ZN(new_n747));
  AOI21_X1  g322(.A(KEYINPUT86), .B1(new_n747), .B2(new_n461), .ZN(new_n748));
  OAI221_X1 g323(.A(G2104), .B1(G116), .B2(new_n461), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G140), .ZN(new_n750));
  INV_X1    g325(.A(G128), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n469), .A2(G2105), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n749), .B1(new_n470), .B2(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n744), .B1(new_n754), .B2(new_n718), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n726), .B2(new_n725), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n723), .A2(new_n742), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n683), .A2(G19), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n550), .B2(new_n683), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G1341), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n599), .A2(G16), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n683), .A2(G4), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n766), .B2(new_n765), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n721), .A2(new_n722), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n761), .A2(G1341), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n759), .A2(new_n768), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n718), .A2(G32), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n464), .A2(G105), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n480), .A2(G141), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n483), .A2(G129), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT26), .Z(new_n777));
  NAND4_X1  g352(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n772), .B1(new_n779), .B2(new_n718), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n683), .A2(G5), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G171), .B2(new_n683), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n783), .B1(new_n731), .B2(G2084), .C1(new_n785), .C2(G1961), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT89), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT30), .B(G28), .ZN(new_n788));
  OR2_X1    g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  NAND2_X1  g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n788), .A2(new_n718), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n626), .B2(new_n718), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT88), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n740), .A2(G2072), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G168), .A2(new_n683), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n683), .B2(G21), .ZN(new_n796));
  INV_X1    g371(.A(G1966), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI211_X1 g373(.A(new_n794), .B(new_n798), .C1(new_n793), .C2(new_n792), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n780), .A2(new_n782), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT87), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n797), .B2(new_n796), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n785), .A2(G1961), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n683), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT23), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G299), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1956), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n799), .A2(new_n802), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n771), .A2(new_n787), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n717), .A2(new_n809), .ZN(G311));
  NAND2_X1  g385(.A1(new_n717), .A2(new_n809), .ZN(G150));
  XNOR2_X1  g386(.A(KEYINPUT90), .B(G55), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n502), .A2(G543), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n513), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n526), .A2(new_n527), .A3(G67), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n495), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT92), .B(G860), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n608), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT91), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n547), .A2(new_n548), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G651), .ZN(new_n829));
  AOI22_X1  g404(.A1(G43), .A2(new_n521), .B1(new_n518), .B2(G81), .ZN(new_n830));
  INV_X1    g405(.A(new_n818), .ZN(new_n831));
  AOI22_X1  g406(.A1(G93), .A2(new_n518), .B1(new_n521), .B2(new_n812), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n546), .A2(new_n549), .B1(new_n815), .B2(new_n818), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n827), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT39), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n824), .B1(new_n838), .B2(new_n821), .ZN(G145));
  XOR2_X1   g414(.A(G160), .B(new_n626), .Z(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(G162), .Z(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n492), .B(new_n753), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n778), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n739), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n483), .A2(G130), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n461), .A2(G118), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(G142), .B2(new_n480), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n617), .B(new_n850), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n710), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT94), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n845), .A2(KEYINPUT94), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(KEYINPUT95), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n845), .A2(new_n852), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n857), .B2(KEYINPUT95), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n842), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n857), .B(new_n842), .C1(new_n852), .C2(new_n845), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(G395));
  INV_X1    g442(.A(G868), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n820), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G290), .B(G166), .ZN(new_n870));
  XOR2_X1   g445(.A(G288), .B(G305), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(KEYINPUT42), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT97), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(KEYINPUT42), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n599), .A2(G299), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n594), .A2(new_n598), .B1(new_n560), .B2(new_n564), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n607), .A2(new_n604), .ZN(new_n882));
  INV_X1    g457(.A(new_n880), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n879), .B2(new_n880), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n610), .B(new_n835), .ZN(new_n889));
  MUX2_X1   g464(.A(new_n881), .B(new_n888), .S(new_n889), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n878), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n869), .B1(new_n891), .B2(new_n868), .ZN(G295));
  OAI21_X1  g467(.A(new_n869), .B1(new_n891), .B2(new_n868), .ZN(G331));
  XNOR2_X1  g468(.A(KEYINPUT98), .B(KEYINPUT43), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n569), .A2(G168), .A3(new_n571), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT99), .B1(G171), .B2(G286), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n569), .A2(G168), .A3(KEYINPUT99), .A4(new_n571), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n835), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n899), .A2(new_n835), .A3(new_n900), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(KEYINPUT100), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n835), .A3(new_n900), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n903), .A2(KEYINPUT101), .A3(new_n881), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n899), .A2(new_n900), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n836), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n899), .A2(new_n835), .A3(KEYINPUT100), .A4(new_n900), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n906), .A2(new_n909), .A3(new_n881), .A4(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n902), .A2(new_n901), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n887), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n870), .A2(new_n871), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n870), .A2(new_n871), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n896), .B1(new_n922), .B2(new_n863), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n916), .B1(new_n907), .B2(new_n913), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n896), .B(new_n863), .C1(new_n924), .C2(new_n872), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n872), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n895), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n906), .A2(new_n909), .A3(new_n910), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n929), .A2(new_n888), .B1(new_n915), .B2(new_n881), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(new_n872), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT103), .B1(new_n930), .B2(new_n872), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n933), .A2(new_n894), .A3(new_n926), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT104), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n887), .B1(new_n903), .B2(new_n906), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n915), .A2(new_n881), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n921), .B(new_n932), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n940), .A2(new_n934), .A3(new_n863), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n894), .A4(new_n926), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n928), .A2(new_n936), .A3(new_n937), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n872), .B1(new_n914), .B2(new_n917), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT102), .B1(new_n945), .B2(G37), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n894), .A3(new_n926), .A4(new_n925), .ZN(new_n947));
  INV_X1    g522(.A(new_n926), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n940), .A2(new_n934), .A3(new_n863), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT44), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n944), .A2(new_n952), .ZN(G397));
  XNOR2_X1  g528(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n492), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n958), .B2(new_n957), .ZN(new_n960));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n471), .A2(new_n474), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n778), .B(G1996), .Z(new_n966));
  XNOR2_X1  g541(.A(new_n753), .B(new_n756), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n713), .B2(new_n710), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n710), .A2(new_n713), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n965), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(G290), .A2(G1986), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n965), .B1(new_n973), .B2(KEYINPUT107), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n973), .A2(KEYINPUT107), .ZN(new_n975));
  NOR2_X1   g550(.A1(G290), .A2(G1986), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n978), .B2(new_n977), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT109), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n492), .A2(new_n956), .A3(new_n955), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT45), .B1(new_n492), .B2(new_n956), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n982), .A2(new_n963), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT113), .B1(new_n984), .B2(G1966), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n986));
  INV_X1    g561(.A(new_n957), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n962), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n986), .B(new_n797), .C1(new_n988), .C2(new_n982), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n957), .A2(KEYINPUT50), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n492), .A2(new_n991), .A3(new_n956), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n962), .A3(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(G2084), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n985), .A2(new_n989), .A3(new_n994), .A4(G168), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT51), .B1(new_n995), .B2(G8), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT121), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n985), .A2(new_n994), .A3(new_n989), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n998), .A2(G8), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n996), .A2(new_n997), .B1(new_n999), .B2(G286), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(G8), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n995), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(KEYINPUT121), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1007));
  OAI21_X1  g582(.A(G8), .B1(new_n963), .B2(new_n957), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G288), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT52), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G305), .A2(G1981), .ZN(new_n1016));
  INV_X1    g591(.A(G1981), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n578), .A2(new_n579), .A3(new_n582), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT49), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1019), .A2(KEYINPUT111), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(KEYINPUT111), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1018), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1008), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G166), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT55), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n962), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n955), .B1(new_n492), .B2(new_n956), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT110), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1971), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n957), .A2(new_n954), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n962), .A4(new_n1031), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n993), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n722), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1028), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1015), .B(new_n1027), .C1(new_n1030), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1030), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT124), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1040), .A2(G1961), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT122), .B(new_n1048), .C1(new_n1049), .C2(G2078), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  AOI21_X1  g626(.A(G2078), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(KEYINPUT53), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1047), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n984), .A2(KEYINPUT53), .A3(new_n726), .ZN(new_n1055));
  AOI21_X1  g630(.A(G301), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1042), .A2(new_n1030), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1008), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n1025), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .A4(new_n1044), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1046), .A2(new_n1056), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1000), .A2(new_n1005), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1007), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT125), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1007), .A2(new_n1063), .A3(new_n1068), .A4(new_n1065), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1045), .A2(new_n1060), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1018), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G288), .A2(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1027), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1008), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n998), .A2(G8), .A3(G168), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(KEYINPUT114), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(KEYINPUT63), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1077), .B(new_n1078), .C1(new_n1080), .C2(KEYINPUT63), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1075), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n560), .B2(new_n564), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(G2072), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1036), .A2(new_n962), .A3(new_n1031), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT117), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1031), .A2(new_n962), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n1036), .A4(new_n1090), .ZN(new_n1095));
  INV_X1    g670(.A(G1956), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n993), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1088), .A2(new_n1092), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT118), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n963), .A2(new_n957), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n993), .A2(new_n766), .B1(new_n1100), .B2(new_n756), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(new_n599), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1092), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1088), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1099), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT58), .B(G1341), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1032), .A2(G1996), .A3(new_n1033), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n550), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT59), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1101), .A2(new_n599), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1102), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1106), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1101), .A2(new_n1116), .A3(new_n607), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1106), .B(KEYINPUT119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(new_n1099), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1121), .B2(KEYINPUT120), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(new_n1119), .C1(new_n1120), .C2(new_n1099), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1107), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1047), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1032), .A2(new_n1048), .A3(G2078), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n960), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT123), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(new_n572), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1126), .B1(new_n1133), .B2(new_n1056), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1046), .A2(new_n1062), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(G171), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1054), .A2(G301), .A3(new_n1055), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(KEYINPUT54), .A3(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .A4(new_n1006), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1084), .B1(new_n1125), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n981), .B1(new_n1070), .B2(new_n1140), .ZN(new_n1141));
  OR3_X1    g716(.A1(new_n965), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT46), .B1(new_n965), .B2(G1996), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n967), .A2(new_n779), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1142), .A2(new_n1143), .B1(new_n964), .B2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT47), .Z(new_n1146));
  INV_X1    g721(.A(new_n968), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n970), .B1(new_n965), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(G2067), .B2(new_n753), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(KEYINPUT126), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n964), .B1(new_n1149), .B2(KEYINPUT126), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n976), .A2(new_n964), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT127), .Z(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT48), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(KEYINPUT48), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(new_n972), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1152), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1141), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g734(.A1(G229), .A2(new_n459), .A3(new_n644), .A4(G227), .ZN(new_n1161));
  OAI21_X1  g735(.A(new_n1161), .B1(new_n861), .B2(new_n864), .ZN(new_n1162));
  AND2_X1   g736(.A1(new_n936), .A2(new_n943), .ZN(new_n1163));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n1163), .B2(new_n928), .ZN(G308));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n928), .ZN(new_n1165));
  INV_X1    g739(.A(new_n1162), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1166), .ZN(G225));
endmodule


