

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U551 ( .A1(n750), .A2(n749), .ZN(n752) );
  AND2_X2 U552 ( .A1(n534), .A2(G2104), .ZN(n879) );
  XOR2_X1 U553 ( .A(KEYINPUT99), .B(n740), .Z(n514) );
  OR2_X1 U554 ( .A1(n759), .A2(n748), .ZN(n515) );
  XOR2_X1 U555 ( .A(KEYINPUT75), .B(n525), .Z(n516) );
  XNOR2_X1 U556 ( .A(KEYINPUT90), .B(n718), .ZN(n702) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n700) );
  XNOR2_X1 U558 ( .A(n701), .B(n700), .ZN(n707) );
  OR2_X1 U559 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U560 ( .A1(n792), .A2(n794), .ZN(n718) );
  NAND2_X1 U561 ( .A1(n955), .A2(n515), .ZN(n749) );
  INV_X1 U562 ( .A(KEYINPUT101), .ZN(n751) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n794) );
  INV_X1 U564 ( .A(G651), .ZN(n522) );
  NOR2_X1 U565 ( .A1(n626), .A2(n522), .ZN(n632) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n634) );
  NOR2_X2 U567 ( .A1(G2104), .A2(n534), .ZN(n882) );
  NOR2_X1 U568 ( .A1(G651), .A2(n626), .ZN(n641) );
  XNOR2_X1 U569 ( .A(n530), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U570 ( .A1(G89), .A2(n634), .ZN(n517) );
  XNOR2_X1 U571 ( .A(n517), .B(KEYINPUT4), .ZN(n518) );
  XNOR2_X1 U572 ( .A(n518), .B(KEYINPUT74), .ZN(n520) );
  XOR2_X1 U573 ( .A(G543), .B(KEYINPUT0), .Z(n626) );
  NAND2_X1 U574 ( .A1(G76), .A2(n632), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U576 ( .A(n521), .B(KEYINPUT5), .ZN(n529) );
  NOR2_X1 U577 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U578 ( .A(KEYINPUT66), .B(n523), .Z(n524) );
  XNOR2_X2 U579 ( .A(KEYINPUT1), .B(n524), .ZN(n635) );
  NAND2_X1 U580 ( .A1(G63), .A2(n635), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n641), .A2(G51), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n516), .A2(n526), .ZN(n527) );
  XOR2_X1 U583 ( .A(KEYINPUT6), .B(n527), .Z(n528) );
  NAND2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  XOR2_X2 U586 ( .A(n531), .B(KEYINPUT17), .Z(n878) );
  NAND2_X1 U587 ( .A1(n878), .A2(G138), .ZN(n538) );
  INV_X1 U588 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U589 ( .A1(G126), .A2(n882), .ZN(n533) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U591 ( .A1(G114), .A2(n883), .ZN(n532) );
  AND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U593 ( .A1(G102), .A2(n879), .ZN(n535) );
  AND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n537) );
  AND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U596 ( .A1(G85), .A2(n634), .ZN(n540) );
  NAND2_X1 U597 ( .A1(G60), .A2(n635), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G72), .A2(n632), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G47), .A2(n641), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U602 ( .A1(n544), .A2(n543), .ZN(G290) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U604 ( .A1(n641), .A2(G53), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G65), .A2(n635), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G91), .A2(n634), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G78), .A2(n632), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n963) );
  INV_X1 U611 ( .A(n963), .ZN(G299) );
  INV_X1 U612 ( .A(G57), .ZN(G237) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  NAND2_X1 U614 ( .A1(n641), .A2(G52), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G64), .A2(n635), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT67), .B(n553), .Z(n558) );
  NAND2_X1 U618 ( .A1(G90), .A2(n634), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G77), .A2(n632), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U622 ( .A1(n558), .A2(n557), .ZN(G171) );
  NAND2_X1 U623 ( .A1(G88), .A2(n634), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G75), .A2(n632), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n641), .A2(G50), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G62), .A2(n635), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(G166) );
  XOR2_X1 U630 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n566) );
  NAND2_X1 U631 ( .A1(G101), .A2(n879), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G113), .A2(n883), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT65), .B(n567), .Z(n568) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G137), .A2(n878), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G125), .A2(n882), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(G160) );
  XOR2_X1 U640 ( .A(G168), .B(KEYINPUT8), .Z(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT76), .B(n574), .ZN(G286) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U644 ( .A(G223), .B(KEYINPUT69), .ZN(n815) );
  NAND2_X1 U645 ( .A1(n815), .A2(G567), .ZN(n576) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  XOR2_X1 U647 ( .A(G860), .B(KEYINPUT72), .Z(n600) );
  NAND2_X1 U648 ( .A1(G81), .A2(n634), .ZN(n577) );
  XNOR2_X1 U649 ( .A(n577), .B(KEYINPUT12), .ZN(n578) );
  XNOR2_X1 U650 ( .A(n578), .B(KEYINPUT70), .ZN(n580) );
  NAND2_X1 U651 ( .A1(G68), .A2(n632), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U653 ( .A(KEYINPUT13), .B(n581), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n635), .A2(G56), .ZN(n582) );
  XOR2_X1 U655 ( .A(KEYINPUT14), .B(n582), .Z(n585) );
  NAND2_X1 U656 ( .A1(G43), .A2(n641), .ZN(n583) );
  XNOR2_X1 U657 ( .A(KEYINPUT71), .B(n583), .ZN(n584) );
  NOR2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n959) );
  OR2_X1 U660 ( .A1(n600), .A2(n959), .ZN(G153) );
  INV_X1 U661 ( .A(G868), .ZN(n653) );
  NOR2_X1 U662 ( .A1(n653), .A2(G171), .ZN(n588) );
  XNOR2_X1 U663 ( .A(n588), .B(KEYINPUT73), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G92), .A2(n634), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G79), .A2(n632), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n641), .A2(G54), .ZN(n592) );
  NAND2_X1 U668 ( .A1(G66), .A2(n635), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U671 ( .A(KEYINPUT15), .B(n595), .ZN(n894) );
  NAND2_X1 U672 ( .A1(n653), .A2(n894), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(G284) );
  NAND2_X1 U674 ( .A1(G868), .A2(G286), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G299), .A2(n653), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n600), .A2(G559), .ZN(n601) );
  INV_X1 U678 ( .A(n894), .ZN(n973) );
  NAND2_X1 U679 ( .A1(n601), .A2(n973), .ZN(n602) );
  XNOR2_X1 U680 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n959), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G868), .A2(n973), .ZN(n603) );
  NOR2_X1 U683 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U684 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n882), .ZN(n606) );
  XOR2_X1 U686 ( .A(KEYINPUT18), .B(n606), .Z(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT77), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G135), .A2(n878), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U690 ( .A(KEYINPUT78), .B(n610), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G111), .A2(n883), .ZN(n612) );
  NAND2_X1 U692 ( .A1(G99), .A2(n879), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n915) );
  XOR2_X1 U695 ( .A(G2096), .B(n915), .Z(n615) );
  NOR2_X1 U696 ( .A1(G2100), .A2(n615), .ZN(n616) );
  XNOR2_X1 U697 ( .A(KEYINPUT79), .B(n616), .ZN(G156) );
  NAND2_X1 U698 ( .A1(n641), .A2(G55), .ZN(n618) );
  NAND2_X1 U699 ( .A1(G67), .A2(n635), .ZN(n617) );
  NAND2_X1 U700 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n634), .A2(G93), .ZN(n619) );
  XOR2_X1 U702 ( .A(KEYINPUT80), .B(n619), .Z(n620) );
  NOR2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n632), .A2(G80), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n654) );
  NAND2_X1 U706 ( .A1(n973), .A2(G559), .ZN(n651) );
  XNOR2_X1 U707 ( .A(n959), .B(n651), .ZN(n624) );
  NOR2_X1 U708 ( .A1(G860), .A2(n624), .ZN(n625) );
  XOR2_X1 U709 ( .A(n654), .B(n625), .Z(G145) );
  NAND2_X1 U710 ( .A1(G87), .A2(n626), .ZN(n628) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U713 ( .A1(n635), .A2(n629), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n641), .A2(G49), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G73), .A2(n632), .ZN(n633) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n633), .Z(n640) );
  NAND2_X1 U718 ( .A1(G86), .A2(n634), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G61), .A2(n635), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U721 ( .A(KEYINPUT81), .B(n638), .Z(n639) );
  NOR2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n641), .A2(G48), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(G305) );
  XOR2_X1 U725 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n644) );
  XNOR2_X1 U726 ( .A(n959), .B(n644), .ZN(n645) );
  XNOR2_X1 U727 ( .A(G288), .B(n645), .ZN(n647) );
  XOR2_X1 U728 ( .A(G299), .B(G166), .Z(n646) );
  XNOR2_X1 U729 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U730 ( .A(n648), .B(G290), .ZN(n649) );
  XNOR2_X1 U731 ( .A(n649), .B(n654), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n650), .B(G305), .ZN(n896) );
  XNOR2_X1 U733 ( .A(n896), .B(n651), .ZN(n652) );
  NOR2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n656) );
  NOR2_X1 U735 ( .A1(G868), .A2(n654), .ZN(n655) );
  NOR2_X1 U736 ( .A1(n656), .A2(n655), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n657) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n658), .ZN(n660) );
  XOR2_X1 U740 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n659) );
  XNOR2_X1 U741 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U742 ( .A1(G2072), .A2(n661), .ZN(G158) );
  XOR2_X1 U743 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  XNOR2_X1 U744 ( .A(KEYINPUT84), .B(G44), .ZN(n662) );
  XNOR2_X1 U745 ( .A(n662), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n663) );
  XNOR2_X1 U747 ( .A(KEYINPUT22), .B(n663), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n664), .A2(G96), .ZN(n665) );
  NOR2_X1 U749 ( .A1(n665), .A2(G218), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n666), .B(KEYINPUT85), .ZN(n820) );
  NAND2_X1 U751 ( .A1(n820), .A2(G2106), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G120), .A2(G69), .ZN(n667) );
  NOR2_X1 U753 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U754 ( .A1(G108), .A2(n668), .ZN(n819) );
  NAND2_X1 U755 ( .A1(G567), .A2(n819), .ZN(n669) );
  XNOR2_X1 U756 ( .A(KEYINPUT86), .B(n669), .ZN(n670) );
  NAND2_X1 U757 ( .A1(n671), .A2(n670), .ZN(n832) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U759 ( .A1(n832), .A2(n672), .ZN(n818) );
  NAND2_X1 U760 ( .A1(n818), .A2(G36), .ZN(G176) );
  INV_X1 U761 ( .A(G166), .ZN(G303) );
  INV_X1 U762 ( .A(G171), .ZN(G301) );
  NAND2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n962) );
  INV_X1 U764 ( .A(n962), .ZN(n674) );
  AND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n792) );
  NAND2_X1 U766 ( .A1(n718), .A2(G8), .ZN(n759) );
  INV_X1 U767 ( .A(KEYINPUT100), .ZN(n743) );
  OR2_X1 U768 ( .A1(n759), .A2(n743), .ZN(n673) );
  NOR2_X1 U769 ( .A1(n674), .A2(n673), .ZN(n741) );
  NOR2_X1 U770 ( .A1(G1976), .A2(G288), .ZN(n744) );
  NOR2_X1 U771 ( .A1(G1971), .A2(G303), .ZN(n675) );
  NOR2_X1 U772 ( .A1(n744), .A2(n675), .ZN(n966) );
  XNOR2_X1 U773 ( .A(KEYINPUT98), .B(n966), .ZN(n739) );
  XOR2_X1 U774 ( .A(KEYINPUT27), .B(KEYINPUT91), .Z(n677) );
  INV_X1 U775 ( .A(n702), .ZN(n689) );
  NAND2_X1 U776 ( .A1(G2072), .A2(n689), .ZN(n676) );
  XNOR2_X1 U777 ( .A(n677), .B(n676), .ZN(n680) );
  NAND2_X1 U778 ( .A1(n702), .A2(G1956), .ZN(n678) );
  XOR2_X1 U779 ( .A(KEYINPUT92), .B(n678), .Z(n679) );
  NOR2_X2 U780 ( .A1(n680), .A2(n679), .ZN(n683) );
  NOR2_X1 U781 ( .A1(n963), .A2(n683), .ZN(n682) );
  XNOR2_X1 U782 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n681) );
  XNOR2_X1 U783 ( .A(n682), .B(n681), .ZN(n699) );
  NAND2_X1 U784 ( .A1(n963), .A2(n683), .ZN(n697) );
  XNOR2_X1 U785 ( .A(G1996), .B(KEYINPUT94), .ZN(n932) );
  INV_X1 U786 ( .A(n718), .ZN(n703) );
  NAND2_X1 U787 ( .A1(n932), .A2(n703), .ZN(n684) );
  XNOR2_X1 U788 ( .A(n684), .B(KEYINPUT26), .ZN(n686) );
  NAND2_X1 U789 ( .A1(n718), .A2(G1341), .ZN(n685) );
  NAND2_X1 U790 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U791 ( .A1(n959), .A2(n687), .ZN(n688) );
  OR2_X1 U792 ( .A1(n973), .A2(n688), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n973), .A2(n688), .ZN(n693) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n689), .ZN(n691) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n718), .ZN(n690) );
  NAND2_X1 U796 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U797 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U798 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U799 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U800 ( .A1(n699), .A2(n698), .ZN(n701) );
  XOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .Z(n937) );
  NOR2_X1 U802 ( .A1(n937), .A2(n702), .ZN(n705) );
  NOR2_X1 U803 ( .A1(n703), .A2(G1961), .ZN(n704) );
  NOR2_X1 U804 ( .A1(n705), .A2(n704), .ZN(n712) );
  OR2_X1 U805 ( .A1(n712), .A2(G301), .ZN(n706) );
  NAND2_X1 U806 ( .A1(n707), .A2(n706), .ZN(n731) );
  XNOR2_X1 U807 ( .A(KEYINPUT30), .B(KEYINPUT95), .ZN(n710) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n759), .ZN(n733) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n718), .ZN(n732) );
  NOR2_X1 U810 ( .A1(n733), .A2(n732), .ZN(n708) );
  NAND2_X1 U811 ( .A1(n708), .A2(G8), .ZN(n709) );
  XOR2_X1 U812 ( .A(n710), .B(n709), .Z(n711) );
  NOR2_X1 U813 ( .A1(G168), .A2(n711), .ZN(n715) );
  NAND2_X1 U814 ( .A1(n712), .A2(G301), .ZN(n713) );
  XOR2_X1 U815 ( .A(KEYINPUT96), .B(n713), .Z(n714) );
  NOR2_X1 U816 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U817 ( .A(KEYINPUT31), .B(n716), .Z(n730) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n759), .ZN(n717) );
  XNOR2_X1 U819 ( .A(KEYINPUT97), .B(n717), .ZN(n721) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n718), .ZN(n719) );
  NOR2_X1 U821 ( .A1(G166), .A2(n719), .ZN(n720) );
  NAND2_X1 U822 ( .A1(n721), .A2(n720), .ZN(n723) );
  AND2_X1 U823 ( .A1(n730), .A2(n723), .ZN(n722) );
  NAND2_X1 U824 ( .A1(n731), .A2(n722), .ZN(n728) );
  INV_X1 U825 ( .A(n723), .ZN(n724) );
  NOR2_X1 U826 ( .A1(n724), .A2(G286), .ZN(n726) );
  INV_X1 U827 ( .A(G8), .ZN(n725) );
  NOR2_X1 U828 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U829 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U830 ( .A(n729), .B(KEYINPUT32), .ZN(n738) );
  AND2_X1 U831 ( .A1(n731), .A2(n730), .ZN(n736) );
  AND2_X1 U832 ( .A1(G8), .A2(n732), .ZN(n734) );
  OR2_X1 U833 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U834 ( .A1(n738), .A2(n737), .ZN(n757) );
  NAND2_X1 U835 ( .A1(n739), .A2(n757), .ZN(n740) );
  AND2_X1 U836 ( .A1(n741), .A2(n514), .ZN(n742) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n742), .ZN(n750) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n955) );
  NAND2_X1 U839 ( .A1(n743), .A2(n744), .ZN(n747) );
  NAND2_X1 U840 ( .A1(n744), .A2(KEYINPUT33), .ZN(n745) );
  NAND2_X1 U841 ( .A1(n745), .A2(KEYINPUT100), .ZN(n746) );
  NAND2_X1 U842 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U843 ( .A(n752), .B(n751), .ZN(n763) );
  NOR2_X1 U844 ( .A1(G1981), .A2(G305), .ZN(n753) );
  XOR2_X1 U845 ( .A(n753), .B(KEYINPUT24), .Z(n754) );
  NOR2_X1 U846 ( .A1(n759), .A2(n754), .ZN(n761) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U848 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U853 ( .A(n764), .B(KEYINPUT102), .ZN(n797) );
  XOR2_X1 U854 ( .A(G2067), .B(KEYINPUT37), .Z(n765) );
  XNOR2_X1 U855 ( .A(KEYINPUT87), .B(n765), .ZN(n808) );
  NAND2_X1 U856 ( .A1(G140), .A2(n878), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G104), .A2(n879), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n768), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G128), .A2(n882), .ZN(n770) );
  NAND2_X1 U861 ( .A1(G116), .A2(n883), .ZN(n769) );
  NAND2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U863 ( .A(KEYINPUT35), .B(n771), .Z(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U865 ( .A(KEYINPUT36), .B(n774), .ZN(n863) );
  NOR2_X1 U866 ( .A1(n808), .A2(n863), .ZN(n804) );
  NAND2_X1 U867 ( .A1(G129), .A2(n882), .ZN(n776) );
  NAND2_X1 U868 ( .A1(G141), .A2(n878), .ZN(n775) );
  NAND2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n879), .A2(G105), .ZN(n777) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(n777), .Z(n778) );
  NOR2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n883), .A2(G117), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n867) );
  NAND2_X1 U875 ( .A1(G1996), .A2(n867), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G119), .A2(n882), .ZN(n782) );
  XNOR2_X1 U877 ( .A(n782), .B(KEYINPUT88), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G107), .A2(n883), .ZN(n784) );
  NAND2_X1 U879 ( .A1(G95), .A2(n879), .ZN(n783) );
  NAND2_X1 U880 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U881 ( .A1(G131), .A2(n878), .ZN(n785) );
  XNOR2_X1 U882 ( .A(KEYINPUT89), .B(n785), .ZN(n786) );
  NOR2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n859) );
  NAND2_X1 U885 ( .A1(G1991), .A2(n859), .ZN(n790) );
  NAND2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n800) );
  NOR2_X1 U887 ( .A1(n804), .A2(n800), .ZN(n917) );
  XOR2_X1 U888 ( .A(G1986), .B(G290), .Z(n970) );
  NAND2_X1 U889 ( .A1(n917), .A2(n970), .ZN(n795) );
  INV_X1 U890 ( .A(n792), .ZN(n793) );
  NOR2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n810) );
  NAND2_X1 U892 ( .A1(n795), .A2(n810), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n813) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n867), .ZN(n912) );
  NOR2_X1 U895 ( .A1(G1991), .A2(n859), .ZN(n918) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n798) );
  XOR2_X1 U897 ( .A(n798), .B(KEYINPUT103), .Z(n799) );
  NOR2_X1 U898 ( .A1(n918), .A2(n799), .ZN(n801) );
  NOR2_X1 U899 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U900 ( .A1(n912), .A2(n802), .ZN(n803) );
  XNOR2_X1 U901 ( .A(n803), .B(KEYINPUT39), .ZN(n806) );
  INV_X1 U902 ( .A(n804), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U904 ( .A(n807), .B(KEYINPUT104), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n808), .A2(n863), .ZN(n926) );
  NAND2_X1 U906 ( .A1(n809), .A2(n926), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U909 ( .A(KEYINPUT40), .B(n814), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n815), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n816) );
  NAND2_X1 U912 ( .A1(G661), .A2(n816), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(G188) );
  XOR2_X1 U915 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  XNOR2_X1 U916 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  XOR2_X1 U917 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U919 ( .A(G96), .ZN(G221) );
  NOR2_X1 U920 ( .A1(n820), .A2(n819), .ZN(G325) );
  INV_X1 U921 ( .A(G325), .ZN(G261) );
  XOR2_X1 U922 ( .A(G2454), .B(G2435), .Z(n822) );
  XNOR2_X1 U923 ( .A(G2438), .B(G2427), .ZN(n821) );
  XNOR2_X1 U924 ( .A(n822), .B(n821), .ZN(n829) );
  XOR2_X1 U925 ( .A(KEYINPUT105), .B(G2446), .Z(n824) );
  XNOR2_X1 U926 ( .A(G2443), .B(G2430), .ZN(n823) );
  XNOR2_X1 U927 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U928 ( .A(n825), .B(G2451), .Z(n827) );
  XNOR2_X1 U929 ( .A(G1341), .B(G1348), .ZN(n826) );
  XNOR2_X1 U930 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U931 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U932 ( .A1(n830), .A2(G14), .ZN(n831) );
  XOR2_X1 U933 ( .A(KEYINPUT106), .B(n831), .Z(n903) );
  XOR2_X1 U934 ( .A(KEYINPUT107), .B(n903), .Z(G401) );
  INV_X1 U935 ( .A(n832), .ZN(G319) );
  XOR2_X1 U936 ( .A(G2100), .B(G2096), .Z(n834) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n833) );
  XNOR2_X1 U938 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2090), .Z(n836) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n835) );
  XNOR2_X1 U941 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U942 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n839) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U945 ( .A(KEYINPUT111), .B(G1956), .Z(n842) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1961), .ZN(n841) );
  XNOR2_X1 U947 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U948 ( .A(n843), .B(KEYINPUT41), .Z(n845) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U950 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U951 ( .A(G1976), .B(G1981), .Z(n847) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1971), .ZN(n846) );
  XNOR2_X1 U953 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U954 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U955 ( .A(KEYINPUT110), .B(G2474), .ZN(n850) );
  XNOR2_X1 U956 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U957 ( .A1(n882), .A2(G124), .ZN(n852) );
  XNOR2_X1 U958 ( .A(n852), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U959 ( .A1(G100), .A2(n879), .ZN(n853) );
  NAND2_X1 U960 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G112), .A2(n883), .ZN(n856) );
  NAND2_X1 U962 ( .A1(G136), .A2(n878), .ZN(n855) );
  NAND2_X1 U963 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U964 ( .A1(n858), .A2(n857), .ZN(G162) );
  XNOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n859), .B(G164), .ZN(n860) );
  XNOR2_X1 U967 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U968 ( .A(KEYINPUT113), .B(n862), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n863), .B(KEYINPUT48), .ZN(n864) );
  XNOR2_X1 U970 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n915), .B(n866), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n867), .B(G160), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n869), .B(n868), .ZN(n892) );
  NAND2_X1 U974 ( .A1(G142), .A2(n878), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G106), .A2(n879), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n872), .B(KEYINPUT45), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G130), .A2(n882), .ZN(n874) );
  NAND2_X1 U979 ( .A1(G118), .A2(n883), .ZN(n873) );
  NAND2_X1 U980 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U981 ( .A(KEYINPUT112), .B(n875), .Z(n876) );
  NAND2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G139), .A2(n878), .ZN(n881) );
  NAND2_X1 U984 ( .A1(G103), .A2(n879), .ZN(n880) );
  NAND2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G127), .A2(n882), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G115), .A2(n883), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n886), .Z(n887) );
  NOR2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n906) );
  XNOR2_X1 U991 ( .A(n889), .B(n906), .ZN(n890) );
  XNOR2_X1 U992 ( .A(G162), .B(n890), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U994 ( .A1(G37), .A2(n893), .ZN(G395) );
  XOR2_X1 U995 ( .A(G301), .B(n894), .Z(n895) );
  XNOR2_X1 U996 ( .A(n895), .B(G286), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U998 ( .A1(G37), .A2(n898), .ZN(G397) );
  XNOR2_X1 U999 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n900) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n901), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1007 ( .A(G2072), .B(n906), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(G164), .B(G2078), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n907), .B(KEYINPUT118), .ZN(n908) );
  NAND2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(n910), .B(KEYINPUT50), .ZN(n924) );
  XOR2_X1 U1012 ( .A(G2090), .B(G162), .Z(n911) );
  NOR2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1014 ( .A(KEYINPUT51), .B(n913), .Z(n922) );
  XOR2_X1 U1015 ( .A(G160), .B(G2084), .Z(n914) );
  NOR2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1019 ( .A(KEYINPUT117), .B(n920), .Z(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n927), .B(KEYINPUT119), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(KEYINPUT52), .B(n928), .ZN(n930) );
  INV_X1 U1025 ( .A(KEYINPUT55), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n931), .A2(G29), .ZN(n1012) );
  XNOR2_X1 U1028 ( .A(G2090), .B(G35), .ZN(n946) );
  XOR2_X1 U1029 ( .A(G2072), .B(G33), .Z(n936) );
  XNOR2_X1 U1030 ( .A(n932), .B(G32), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(G26), .B(G2067), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(G27), .B(n937), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(KEYINPUT120), .B(n940), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n941), .A2(G28), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G25), .B(G1991), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(KEYINPUT53), .B(n944), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1042 ( .A(G2084), .B(G34), .Z(n947) );
  XNOR2_X1 U1043 ( .A(KEYINPUT54), .B(n947), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1045 ( .A(KEYINPUT55), .B(n950), .Z(n952) );
  INV_X1 U1046 ( .A(G29), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(G11), .A2(n953), .ZN(n1010) );
  XNOR2_X1 U1049 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n954) );
  XOR2_X1 U1050 ( .A(G16), .B(n954), .Z(n982) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT122), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT57), .B(n958), .ZN(n980) );
  XNOR2_X1 U1055 ( .A(G1341), .B(KEYINPUT124), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(n960), .B(n959), .ZN(n972) );
  NAND2_X1 U1057 ( .A1(G1971), .A2(G303), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G1956), .B(KEYINPUT123), .ZN(n964) );
  XOR2_X1 U1060 ( .A(n964), .B(n963), .Z(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n977) );
  XOR2_X1 U1065 ( .A(G171), .B(G1961), .Z(n975) );
  XOR2_X1 U1066 ( .A(n973), .B(G1348), .Z(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(KEYINPUT125), .B(n978), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n1008) );
  INV_X1 U1072 ( .A(G16), .ZN(n1006) );
  XNOR2_X1 U1073 ( .A(G1986), .B(G24), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1976), .B(G23), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT127), .B(n985), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(KEYINPUT58), .B(n988), .Z(n1003) );
  XOR2_X1 U1080 ( .A(G1961), .B(G5), .Z(n998) );
  XNOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(G4), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(G6), .B(G1981), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(G20), .B(G1956), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(KEYINPUT60), .B(n996), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G21), .B(G1966), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1093 ( .A(KEYINPUT126), .B(n1001), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(KEYINPUT61), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT62), .B(n1013), .ZN(G150) );
  INV_X1 U1101 ( .A(G150), .ZN(G311) );
endmodule

