//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G902), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT64), .A2(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT64), .A2(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(G146), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n195), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT78), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n195), .A2(KEYINPUT78), .A3(new_n198), .A4(new_n200), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G143), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n197), .B1(new_n205), .B2(G146), .ZN(new_n206));
  INV_X1    g020(.A(new_n194), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT64), .A2(G143), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n199), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n203), .B(new_n204), .C1(new_n206), .C2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G104), .B(G107), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(G104), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT77), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(G104), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n219), .B1(new_n217), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n215), .B1(new_n226), .B2(new_n214), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n212), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n217), .ZN(new_n229));
  INV_X1    g043(.A(new_n217), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n222), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n214), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n215), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n208), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n210), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  OAI21_X1  g052(.A(G128), .B1(new_n197), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n234), .A2(new_n240), .A3(new_n201), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n228), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT11), .A3(G134), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(G137), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  INV_X1    g065(.A(G131), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n245), .A2(new_n247), .A3(new_n252), .A4(new_n248), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(KEYINPUT66), .A3(G131), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT12), .B1(new_n242), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n259), .B(new_n256), .C1(new_n228), .C2(new_n241), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT80), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT10), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n228), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n230), .B1(new_n213), .B2(new_n221), .ZN(new_n264));
  OAI21_X1  g078(.A(G101), .B1(new_n264), .B2(new_n219), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT4), .A3(new_n232), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n210), .B2(new_n236), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n195), .A2(new_n267), .A3(new_n198), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n195), .A2(KEYINPUT65), .A3(new_n267), .A4(new_n198), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(G101), .C1(new_n264), .C2(new_n219), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n266), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n193), .A2(new_n194), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n235), .B1(new_n279), .B2(new_n208), .ZN(new_n280));
  INV_X1    g094(.A(new_n239), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n201), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n263), .A2(new_n256), .A3(new_n278), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G110), .B(G140), .ZN(new_n285));
  INV_X1    g099(.A(G953), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n286), .A2(G227), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n285), .B(new_n287), .Z(new_n288));
  AND2_X1   g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n193), .A2(new_n194), .A3(G146), .ZN(new_n290));
  OAI21_X1  g104(.A(G128), .B1(new_n290), .B2(new_n238), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n195), .A2(new_n198), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n291), .A2(new_n292), .B1(new_n201), .B2(new_n202), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n234), .B1(new_n204), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n227), .A2(new_n282), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n257), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n259), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n242), .A2(KEYINPUT12), .A3(new_n257), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT80), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n261), .A2(new_n289), .A3(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n278), .B(new_n283), .C1(new_n294), .C2(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT79), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT79), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n263), .A2(new_n304), .A3(new_n278), .A4(new_n283), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n257), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n288), .B1(new_n306), .B2(new_n284), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n191), .B(new_n192), .C1(new_n301), .C2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n191), .A2(new_n192), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n284), .B1(new_n258), .B2(new_n260), .ZN(new_n310));
  INV_X1    g124(.A(new_n288), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n306), .A2(new_n289), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n309), .B1(new_n312), .B2(G469), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n190), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G214), .B1(G237), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G210), .B1(G237), .B2(G902), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OR2_X1    g132(.A1(KEYINPUT2), .A2(G113), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT2), .A2(G113), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G116), .ZN(new_n323));
  INV_X1    g137(.A(G116), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n319), .A2(new_n323), .A3(new_n325), .A4(new_n320), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(KEYINPUT67), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n321), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n266), .A2(new_n332), .A3(new_n277), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n322), .A3(G116), .ZN(new_n335));
  OAI211_X1 g149(.A(G113), .B(new_n335), .C1(new_n326), .C2(new_n334), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n336), .A2(KEYINPUT81), .ZN(new_n337));
  INV_X1    g151(.A(new_n328), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n336), .B2(KEYINPUT81), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n227), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G122), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n333), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n333), .A2(new_n340), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(KEYINPUT82), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n333), .B2(new_n340), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT6), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT84), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n282), .B2(G125), .ZN(new_n352));
  INV_X1    g166(.A(G125), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n240), .A2(KEYINPUT84), .A3(new_n353), .A4(new_n201), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n356));
  INV_X1    g170(.A(new_n270), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT65), .B1(new_n206), .B2(new_n267), .ZN(new_n358));
  INV_X1    g172(.A(new_n274), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n356), .B1(new_n360), .B2(G125), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n275), .A2(KEYINPUT83), .A3(new_n353), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n355), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G224), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G953), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n360), .A2(new_n356), .A3(G125), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT83), .B1(new_n275), .B2(new_n353), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n365), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n355), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n348), .A2(new_n350), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n369), .A2(KEYINPUT7), .A3(new_n370), .A4(new_n355), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n333), .A2(new_n340), .A3(new_n341), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n234), .A2(new_n337), .A3(new_n339), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n341), .B(KEYINPUT8), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n336), .A2(new_n328), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n376), .B(new_n377), .C1(new_n234), .C2(new_n378), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n352), .A2(new_n354), .B1(new_n360), .B2(G125), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n370), .B1(new_n381), .B2(KEYINPUT7), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n381), .B2(KEYINPUT7), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n375), .B(new_n379), .C1(new_n380), .C2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n192), .B1(new_n374), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n318), .B1(new_n372), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n384), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n387), .B2(new_n373), .ZN(new_n388));
  INV_X1    g202(.A(new_n371), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n370), .B1(new_n369), .B2(new_n355), .ZN(new_n390));
  INV_X1    g204(.A(new_n350), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n375), .B1(new_n349), .B2(KEYINPUT6), .ZN(new_n392));
  OAI22_X1  g206(.A1(new_n389), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n393), .A3(new_n317), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n316), .B1(new_n386), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G237), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n396), .A2(new_n286), .A3(G214), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n279), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n286), .A3(G214), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n196), .ZN(new_n400));
  OAI21_X1  g214(.A(G131), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT17), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n205), .A2(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n397), .A2(G143), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n252), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n252), .B1(new_n403), .B2(new_n404), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT17), .ZN(new_n408));
  INV_X1    g222(.A(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n353), .A2(G140), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n353), .A2(KEYINPUT16), .A3(G140), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(G146), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT72), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(G146), .B1(new_n412), .B2(new_n413), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n413), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT72), .A3(new_n208), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n406), .B(new_n408), .C1(new_n418), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n407), .A2(KEYINPUT18), .ZN(new_n423));
  OR3_X1    g237(.A1(new_n398), .A2(KEYINPUT18), .A3(new_n400), .ZN(new_n424));
  XNOR2_X1  g238(.A(G125), .B(G140), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(new_n208), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n423), .A2(new_n424), .A3(new_n426), .A4(new_n405), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT90), .B(G104), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n428), .B(new_n429), .Z(new_n430));
  AND3_X1   g244(.A1(new_n422), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n430), .B1(new_n422), .B2(new_n427), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n192), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT91), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(new_n192), .C1(new_n431), .C2(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(G475), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(G475), .A2(G902), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT89), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT88), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT19), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n425), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n439), .B(new_n414), .C1(new_n444), .C2(G146), .ZN(new_n445));
  INV_X1    g259(.A(new_n405), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT87), .B1(new_n446), .B2(new_n407), .ZN(new_n447));
  AOI21_X1  g261(.A(G146), .B1(new_n442), .B2(new_n443), .ZN(new_n448));
  INV_X1    g262(.A(new_n414), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT89), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n401), .A2(new_n451), .A3(new_n405), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n445), .A2(new_n447), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n430), .B1(new_n453), .B2(new_n427), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n438), .B1(new_n454), .B2(new_n431), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n458), .B(new_n438), .C1(new_n454), .C2(new_n431), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n437), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n205), .A2(G128), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n196), .A2(G128), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G134), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n244), .A3(new_n464), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT92), .B1(new_n324), .B2(G122), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n324), .A2(KEYINPUT92), .A3(G122), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n324), .A2(G122), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n218), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n466), .A2(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(KEYINPUT14), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT14), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n477), .A3(new_n470), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G107), .ZN(new_n480));
  INV_X1    g294(.A(new_n473), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT93), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n462), .A2(KEYINPUT13), .A3(new_n464), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n484), .B(G134), .C1(KEYINPUT13), .C2(new_n462), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n218), .B1(new_n471), .B2(new_n472), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n485), .B(new_n467), .C1(new_n486), .C2(new_n481), .ZN(new_n487));
  INV_X1    g301(.A(G217), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n188), .A2(new_n488), .A3(G953), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n483), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n483), .B2(new_n487), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n192), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI221_X1 g309(.A(new_n192), .B1(KEYINPUT15), .B2(new_n493), .C1(new_n490), .C2(new_n491), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(G234), .A2(G237), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n498), .A2(G952), .A3(new_n286), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT21), .B(G898), .Z(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n498), .A2(G902), .A3(G953), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n461), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n314), .A2(new_n395), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n248), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n244), .A2(G137), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n282), .A2(new_n253), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n329), .A2(new_n331), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n509), .B(new_n510), .C1(new_n360), .C2(new_n256), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT28), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n513), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT71), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(KEYINPUT70), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n275), .A2(new_n255), .A3(new_n254), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n510), .B1(new_n519), .B2(new_n509), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI211_X1 g335(.A(KEYINPUT70), .B(new_n510), .C1(new_n519), .C2(new_n509), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n514), .B(new_n516), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT26), .B(G101), .Z(new_n524));
  NAND3_X1  g338(.A1(new_n396), .A2(new_n286), .A3(G210), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n509), .B1(new_n360), .B2(new_n256), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n519), .A2(KEYINPUT30), .A3(new_n509), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n332), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n535), .A2(new_n511), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n528), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT29), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n516), .A2(new_n514), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n531), .A2(new_n332), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n511), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT28), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT29), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n528), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n192), .ZN(new_n546));
  OAI21_X1  g360(.A(G472), .B1(new_n538), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n535), .A2(new_n511), .A3(new_n529), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT31), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n535), .A2(KEYINPUT31), .A3(new_n511), .A4(new_n529), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n551), .A2(new_n552), .B1(new_n523), .B2(new_n528), .ZN(new_n553));
  NOR2_X1   g367(.A1(G472), .A2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n548), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n523), .A2(new_n528), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(KEYINPUT32), .A3(new_n554), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n547), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n286), .A2(G221), .A3(G234), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT74), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT22), .B(G137), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n419), .A2(new_n208), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n415), .A3(new_n414), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n322), .A2(G128), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n199), .A2(G119), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT24), .B(G110), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT23), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(G119), .B2(new_n199), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n322), .A2(KEYINPUT23), .A3(G128), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n569), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n573), .B1(G110), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n568), .A2(new_n420), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G110), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n569), .C1(new_n575), .C2(new_n576), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n571), .A2(new_n572), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n425), .A2(new_n208), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n414), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n566), .B1(new_n579), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n585), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n414), .A4(new_n586), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n568), .A2(new_n420), .A3(new_n578), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n565), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n488), .B1(G234), .B2(new_n192), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n595), .A2(G902), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n589), .A2(new_n594), .A3(new_n192), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT75), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT25), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n589), .A2(new_n594), .A3(KEYINPUT75), .A4(new_n192), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT76), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT76), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n600), .A2(new_n605), .A3(new_n601), .A4(new_n602), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n598), .A2(new_n601), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n597), .B1(new_n608), .B2(new_n596), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n505), .A2(new_n561), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  NAND2_X1  g425(.A1(new_n559), .A2(new_n554), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n553), .B2(G902), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n314), .A2(new_n612), .A3(new_n609), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT94), .Z(new_n615));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n386), .A2(new_n394), .ZN(new_n617));
  INV_X1    g431(.A(new_n503), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n315), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n490), .B2(new_n491), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n483), .A2(new_n487), .ZN(new_n622));
  INV_X1    g436(.A(new_n489), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n483), .A2(new_n487), .A3(new_n489), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(KEYINPUT33), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n493), .A2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n492), .A2(new_n493), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n461), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n616), .B1(new_n619), .B2(new_n631), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n316), .B(new_n503), .C1(new_n386), .C2(new_n394), .ZN(new_n633));
  INV_X1    g447(.A(new_n631), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(KEYINPUT95), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n615), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT96), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n456), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(new_n438), .C1(new_n454), .C2(new_n431), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n457), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n437), .A2(new_n644), .A3(new_n497), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n619), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n615), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NAND2_X1  g463(.A1(new_n613), .A2(new_n612), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n608), .A2(new_n596), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n592), .A2(new_n593), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n566), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n596), .A2(G902), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n505), .A2(new_n651), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  NAND2_X1  g477(.A1(new_n308), .A2(new_n313), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n664), .A2(new_n395), .A3(new_n189), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n502), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n499), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n437), .A2(new_n644), .A3(new_n497), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n665), .A2(new_n561), .A3(new_n671), .A4(new_n658), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NOR2_X1   g487(.A1(new_n536), .A2(new_n528), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n192), .B1(new_n541), .B2(new_n529), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n556), .A2(new_n560), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n556), .A2(new_n560), .A3(KEYINPUT100), .A4(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n658), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n669), .B(KEYINPUT39), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n314), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n617), .B(KEYINPUT38), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n461), .A2(new_n497), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n689), .A2(new_n316), .A3(new_n690), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n683), .A2(new_n687), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n205), .ZN(G45));
  INV_X1    g507(.A(new_n669), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n631), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n665), .A2(new_n561), .A3(new_n658), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  OAI21_X1  g511(.A(new_n192), .B1(new_n301), .B2(new_n307), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n699), .A2(new_n189), .A3(new_n308), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n561), .A2(new_n700), .A3(new_n609), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n636), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT41), .B(G113), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  AND4_X1   g518(.A1(new_n395), .A2(new_n699), .A3(new_n189), .A4(new_n308), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n561), .A3(new_n646), .A4(new_n609), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NAND4_X1  g521(.A1(new_n705), .A2(new_n561), .A3(new_n504), .A4(new_n658), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NOR2_X1   g523(.A1(new_n619), .A2(new_n690), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n542), .A2(new_n514), .A3(new_n516), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n551), .A2(new_n552), .B1(new_n711), .B2(new_n528), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n555), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n559), .A2(new_n192), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT101), .B(G472), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n710), .A2(new_n700), .A3(new_n609), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  AOI21_X1  g532(.A(G902), .B1(new_n557), .B2(new_n558), .ZN(new_n719));
  INV_X1    g533(.A(new_n715), .ZN(new_n720));
  OAI22_X1  g534(.A1(new_n719), .A2(new_n720), .B1(new_n555), .B2(new_n712), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n608), .A2(new_n596), .B1(new_n656), .B2(new_n655), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n705), .A2(new_n723), .A3(new_n695), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n561), .A2(new_n609), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n386), .A2(new_n394), .A3(new_n315), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n695), .A2(new_n314), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n695), .A2(new_n314), .A3(new_n728), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(KEYINPUT102), .A3(new_n561), .A4(new_n609), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(G472), .ZN(new_n735));
  INV_X1    g549(.A(new_n537), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n540), .A2(KEYINPUT70), .A3(new_n511), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n518), .A2(new_n520), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n517), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n528), .B1(new_n539), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n543), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n546), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n735), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n556), .A2(new_n560), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(KEYINPUT103), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(KEYINPUT103), .B2(new_n744), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(KEYINPUT42), .A3(new_n609), .A4(new_n732), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n734), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  AND3_X1   g563(.A1(new_n728), .A2(new_n664), .A3(new_n189), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n561), .A3(new_n671), .A4(new_n609), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n628), .A2(new_n629), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n461), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n755), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  INV_X1    g571(.A(G475), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n422), .A2(new_n427), .ZN(new_n759));
  INV_X1    g573(.A(new_n430), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n422), .A2(new_n427), .A3(new_n430), .ZN(new_n762));
  AOI21_X1  g576(.A(G902), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n758), .B1(new_n763), .B2(new_n435), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n764), .A2(new_n434), .B1(new_n457), .B2(new_n459), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n630), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n757), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  OR3_X1    g583(.A1(new_n766), .A2(KEYINPUT105), .A3(new_n767), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT105), .B1(new_n766), .B2(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(KEYINPUT106), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n651), .A2(new_n722), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT106), .B1(new_n769), .B2(new_n772), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n753), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n776), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n773), .A4(new_n774), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n312), .A2(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n312), .A2(KEYINPUT45), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(G469), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n309), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n308), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n782), .B2(new_n783), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n189), .B(new_n685), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n728), .B(KEYINPUT107), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n777), .A2(new_n779), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  OAI21_X1  g605(.A(new_n189), .B1(new_n785), .B2(new_n786), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n695), .A2(new_n728), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n561), .A2(new_n795), .A3(new_n609), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NOR2_X1   g612(.A1(G952), .A2(G953), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT117), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n769), .A2(new_n772), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n609), .A3(new_n499), .A4(new_n716), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n689), .A2(new_n700), .A3(new_n316), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT50), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n700), .A2(new_n499), .A3(new_n728), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n723), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n682), .A2(new_n609), .A3(new_n806), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n765), .A3(new_n754), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n805), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n699), .A2(new_n308), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n189), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n793), .A2(new_n794), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n802), .A2(new_n788), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n816), .B2(new_n817), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n811), .B(KEYINPUT51), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n807), .A2(new_n609), .A3(new_n746), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n809), .A2(new_n634), .ZN(new_n826));
  INV_X1    g640(.A(new_n705), .ZN(new_n827));
  OAI211_X1 g641(.A(G952), .B(new_n286), .C1(new_n802), .C2(new_n827), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n819), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n816), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n811), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n821), .B(new_n829), .C1(new_n832), .C2(KEYINPUT51), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n765), .B2(new_n754), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n461), .A2(KEYINPUT109), .A3(new_n630), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n633), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT110), .B1(new_n837), .B2(new_n633), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n838), .A2(new_n839), .A3(new_n614), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n561), .A2(new_n665), .A3(new_n609), .A4(new_n504), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT111), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n633), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT110), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n614), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n843), .B(new_n610), .C1(new_n848), .C2(new_n838), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n751), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n658), .A2(new_n314), .A3(new_n669), .A4(new_n728), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n437), .A2(new_n644), .A3(new_n496), .A4(new_n495), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n744), .B2(new_n743), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n716), .A2(new_n634), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT112), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n561), .A2(new_n853), .B1(new_n716), .B2(new_n634), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n751), .B(new_n858), .C1(new_n859), .C2(new_n852), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n659), .B(new_n706), .C1(new_n636), .C2(new_n701), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n633), .A2(new_n765), .A3(new_n497), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n614), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n717), .A3(new_n708), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n850), .A2(new_n861), .A3(new_n748), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n664), .A2(new_n189), .ZN(new_n869));
  INV_X1    g683(.A(new_n395), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n869), .A2(new_n870), .A3(new_n694), .A4(new_n690), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n681), .A2(new_n871), .A3(new_n722), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n672), .A2(new_n696), .A3(new_n724), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n672), .A2(new_n724), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n681), .A2(new_n871), .A3(new_n722), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n696), .A4(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  OR4_X1    g693(.A1(KEYINPUT113), .A2(new_n867), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n867), .B2(new_n878), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n865), .B(new_n862), .C1(new_n842), .C2(new_n849), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n874), .A2(new_n877), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n857), .A2(new_n860), .B1(new_n734), .B2(new_n747), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n882), .A2(KEYINPUT53), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT113), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n880), .A2(KEYINPUT54), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n881), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n800), .B1(new_n833), .B2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n766), .A2(new_n316), .A3(new_n190), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT49), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n609), .B(new_n892), .C1(new_n812), .C2(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT108), .Z(new_n895));
  NAND2_X1  g709(.A1(new_n812), .A2(new_n893), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n682), .A2(new_n689), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n891), .B1(new_n895), .B2(new_n897), .ZN(G75));
  NAND2_X1  g712(.A1(new_n881), .A2(new_n885), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(G902), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT56), .B1(new_n901), .B2(G210), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n389), .A2(new_n391), .A3(new_n392), .A4(new_n390), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n372), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n902), .A2(new_n905), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n286), .A2(G952), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G51));
  NAND2_X1  g723(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n889), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n899), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n309), .B(KEYINPUT57), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n301), .A2(new_n307), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n900), .A2(new_n782), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n908), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(KEYINPUT119), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n918), .B1(new_n915), .B2(new_n916), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n908), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(G54));
  NAND2_X1  g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT120), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n900), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n454), .A2(new_n431), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n921), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n930), .B2(new_n929), .ZN(G60));
  AND2_X1   g746(.A1(new_n621), .A2(new_n626), .ZN(new_n933));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT59), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n890), .B2(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n912), .A2(new_n913), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n933), .A2(new_n935), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n908), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(G63));
  OAI21_X1  g753(.A(new_n921), .B1(KEYINPUT122), .B2(KEYINPUT61), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n488), .A2(new_n192), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n881), .B2(new_n885), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n940), .B1(new_n944), .B2(new_n655), .ZN(new_n945));
  INV_X1    g759(.A(new_n595), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(new_n944), .ZN(new_n947));
  NAND2_X1  g761(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G66));
  OAI21_X1  g763(.A(G953), .B1(new_n501), .B2(new_n364), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n882), .B2(G953), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT123), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n348), .B(new_n350), .C1(G898), .C2(new_n286), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  NAND2_X1  g768(.A1(new_n533), .A2(new_n534), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT124), .Z(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(new_n444), .Z(new_n957));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n790), .A2(new_n797), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n960));
  AOI211_X1 g774(.A(new_n851), .B(new_n873), .C1(new_n734), .C2(new_n747), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n870), .A2(new_n690), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n746), .A2(new_n609), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n964));
  OR3_X1    g778(.A1(new_n963), .A2(new_n964), .A3(new_n787), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n963), .B2(new_n787), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n790), .A3(new_n797), .A4(new_n961), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n286), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n286), .A2(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n958), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(G953), .B1(new_n968), .B2(new_n970), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n976), .A2(KEYINPUT127), .A3(new_n973), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n957), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(G227), .A2(G900), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(G953), .ZN(new_n980));
  INV_X1    g794(.A(new_n957), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n692), .A2(new_n873), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT62), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n837), .B1(new_n765), .B2(new_n497), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n984), .A2(new_n316), .A3(new_n617), .ZN(new_n985));
  INV_X1    g799(.A(new_n727), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n986), .A3(new_n314), .A4(new_n685), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n983), .A2(new_n959), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n981), .B1(new_n988), .B2(G953), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n978), .A2(new_n980), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n972), .A2(new_n958), .A3(new_n974), .ZN(new_n991));
  OAI21_X1  g805(.A(KEYINPUT127), .B1(new_n976), .B2(new_n973), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(G953), .B(new_n979), .C1(new_n993), .C2(new_n981), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n990), .A2(new_n994), .ZN(G72));
  NAND2_X1  g809(.A1(new_n988), .A2(new_n882), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  AOI211_X1 g812(.A(new_n536), .B(new_n528), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n880), .A2(new_n886), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n537), .A2(new_n998), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n1000), .A2(new_n674), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n968), .A2(new_n882), .A3(new_n970), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n537), .B1(new_n1003), .B2(new_n998), .ZN(new_n1004));
  NOR4_X1   g818(.A1(new_n999), .A2(new_n908), .A3(new_n1002), .A4(new_n1004), .ZN(G57));
endmodule


