//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  AND2_X1   g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT67), .B1(new_n188), .B2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT66), .B1(new_n190), .B2(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(new_n190), .A3(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n188), .A3(G143), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n193), .A4(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n187), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n188), .A2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n190), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n203), .A2(new_n187), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT69), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n208), .A2(new_n210), .A3(new_n214), .A4(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G131), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT68), .B(G131), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n196), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n226), .A2(new_n201), .A3(new_n202), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT68), .A2(G131), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT68), .A2(G131), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n209), .A2(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n211), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n230), .A2(new_n233), .B1(G131), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n229), .A2(KEYINPUT70), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n227), .B1(new_n196), .B2(new_n223), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(G131), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n212), .B2(new_n218), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n238), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n205), .A2(new_n221), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  XOR2_X1   g057(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT71), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G119), .ZN(new_n249));
  INV_X1    g063(.A(G119), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT72), .A3(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT2), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G113), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n257), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n260), .A2(new_n251), .A3(new_n252), .A4(new_n249), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n217), .A2(new_n263), .A3(new_n220), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n213), .B2(new_n215), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT73), .B1(new_n266), .B2(new_n219), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n205), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n239), .A2(new_n241), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT74), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n239), .B2(new_n241), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n268), .A2(KEYINPUT30), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT70), .B1(new_n229), .B2(new_n236), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n239), .A2(new_n241), .A3(new_n238), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n266), .A2(new_n219), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n200), .A2(new_n204), .ZN(new_n278));
  OAI22_X1  g092(.A1(new_n275), .A2(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n244), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n246), .A2(new_n262), .A3(new_n274), .A4(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G237), .A2(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G210), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n284), .B(KEYINPUT27), .Z(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G101), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g101(.A(new_n262), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n268), .A2(new_n288), .A3(new_n273), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n282), .A2(KEYINPUT31), .A3(new_n287), .A4(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n268), .A2(new_n288), .A3(new_n273), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n243), .A2(new_n288), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT28), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n269), .A2(new_n262), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n268), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n287), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT75), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n302), .B1(new_n292), .B2(new_n293), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(new_n306), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n301), .B(KEYINPUT77), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n288), .B1(new_n268), .B2(new_n273), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n289), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n315), .B1(new_n318), .B2(KEYINPUT28), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n315), .B(KEYINPUT28), .C1(new_n295), .C2(new_n316), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n314), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n297), .A2(new_n323), .A3(new_n301), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n287), .ZN(new_n325));
  INV_X1    g139(.A(new_n287), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n282), .A2(new_n323), .A3(new_n326), .A4(new_n289), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n322), .A2(KEYINPUT29), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G472), .B1(new_n328), .B2(G902), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n304), .A2(KEYINPUT78), .A3(KEYINPUT32), .A4(new_n307), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n310), .A2(new_n313), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G217), .ZN(new_n332));
  INV_X1    g146(.A(G902), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(G234), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n225), .A2(KEYINPUT23), .A3(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n250), .A2(G128), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT23), .B1(new_n225), .B2(G119), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT80), .B(G110), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n250), .B2(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n225), .A2(KEYINPUT79), .A3(G119), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n336), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n339), .A2(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT16), .ZN(new_n349));
  INV_X1    g163(.A(G140), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(G125), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(G125), .ZN(new_n352));
  INV_X1    g166(.A(G125), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(G146), .B(new_n351), .C1(new_n355), .C2(new_n349), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n346), .A2(new_n347), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n354), .A3(new_n188), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n348), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n351), .B1(new_n355), .B2(new_n349), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n188), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n356), .ZN(new_n362));
  INV_X1    g176(.A(G110), .ZN(new_n363));
  OAI221_X1 g177(.A(new_n362), .B1(new_n363), .B2(new_n339), .C1(new_n344), .C2(new_n345), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT22), .B(G137), .ZN(new_n366));
  INV_X1    g180(.A(G953), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n367), .A2(G221), .A3(G234), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n366), .B(new_n368), .Z(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n369), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n359), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n373), .A2(KEYINPUT25), .A3(new_n333), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT25), .B1(new_n373), .B2(new_n333), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n334), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n334), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n333), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT82), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n373), .A2(new_n380), .A3(new_n333), .A4(new_n377), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G221), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT9), .B(G234), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n387), .B2(new_n333), .ZN(new_n388));
  XNOR2_X1  g202(.A(G110), .B(G140), .ZN(new_n389));
  INV_X1    g203(.A(G227), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n389), .B(new_n391), .Z(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G101), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n395), .A2(new_n398), .A3(new_n402), .A4(new_n399), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n405), .A3(G101), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n404), .B(new_n406), .C1(new_n200), .C2(new_n204), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n394), .A2(G107), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n397), .A2(G104), .ZN(new_n409));
  OAI21_X1  g223(.A(G101), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n229), .A2(KEYINPUT10), .A3(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT84), .B(KEYINPUT1), .C1(new_n190), .C2(G146), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT84), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n416));
  OAI21_X1  g230(.A(G128), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n203), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n411), .B1(new_n418), .B2(new_n228), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n407), .B(new_n413), .C1(new_n419), .C2(KEYINPUT10), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n263), .B1(new_n217), .B2(new_n220), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n266), .A2(KEYINPUT73), .A3(new_n219), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT85), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n264), .A2(new_n424), .A3(new_n267), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n420), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n264), .A2(new_n267), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n419), .A2(KEYINPUT10), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n407), .A2(new_n413), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n393), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(KEYINPUT88), .B(new_n393), .C1(new_n426), .C2(new_n430), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n239), .A2(new_n411), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n227), .B1(new_n417), .B2(new_n203), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(new_n411), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n264), .A3(new_n267), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT86), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n438), .A2(KEYINPUT12), .A3(new_n221), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT87), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n442), .A2(new_n448), .A3(new_n444), .A4(new_n445), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n426), .A2(new_n393), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n435), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G469), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n333), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n423), .A2(new_n425), .ZN(new_n455));
  INV_X1    g269(.A(new_n420), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n392), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n430), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n446), .A2(new_n457), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n392), .B(KEYINPUT83), .Z(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G469), .B1(new_n462), .B2(G902), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n388), .B1(new_n454), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G214), .B1(G237), .B2(G902), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G122), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n404), .A2(KEYINPUT89), .A3(new_n262), .A4(new_n406), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT90), .B(KEYINPUT5), .Z(new_n469));
  NOR2_X1   g283(.A1(new_n248), .A2(G119), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n254), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n253), .A2(new_n469), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n412), .B(new_n261), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n400), .A2(G101), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n476), .A2(new_n405), .B1(new_n259), .B2(new_n261), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT89), .B1(new_n477), .B2(new_n404), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n467), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(KEYINPUT6), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n205), .A2(new_n353), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n229), .A2(G125), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G224), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G953), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n483), .B(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n404), .A2(new_n262), .A3(new_n406), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n468), .A3(new_n474), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT91), .B1(new_n490), .B2(new_n467), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n489), .A2(new_n468), .A3(new_n474), .A4(new_n466), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT6), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n490), .A2(KEYINPUT91), .A3(new_n467), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT92), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n492), .A2(KEYINPUT6), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n479), .A2(new_n498), .ZN(new_n499));
  AND4_X1   g313(.A1(KEYINPUT92), .A2(new_n497), .A3(new_n499), .A4(new_n495), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n480), .B(new_n486), .C1(new_n496), .C2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G210), .B1(G237), .B2(G902), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n503));
  OR4_X1    g317(.A1(new_n503), .A2(new_n481), .A3(new_n485), .A4(new_n482), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n483), .B1(new_n503), .B2(new_n485), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n261), .B(new_n411), .C1(new_n472), .C2(new_n473), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n466), .B(KEYINPUT8), .ZN(new_n507));
  INV_X1    g321(.A(new_n261), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT5), .A4(new_n252), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(new_n471), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n506), .B(new_n507), .C1(new_n510), .C2(new_n411), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n504), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n512), .B2(new_n492), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n501), .A2(new_n502), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n502), .B1(new_n501), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n465), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n517));
  INV_X1    g331(.A(G237), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n367), .A3(G214), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n190), .ZN(new_n520));
  AOI21_X1  g334(.A(G143), .B1(new_n283), .B2(G214), .ZN(new_n521));
  OAI211_X1 g335(.A(KEYINPUT18), .B(G131), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n190), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n283), .A2(G143), .A3(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n355), .A2(G146), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n358), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n522), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n233), .B1(new_n523), .B2(new_n524), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n361), .A3(new_n356), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n520), .A2(new_n521), .A3(new_n218), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n533), .A2(new_n530), .A3(KEYINPUT17), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n529), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G113), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(new_n394), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n352), .A2(new_n354), .A3(KEYINPUT19), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT19), .B1(new_n352), .B2(new_n354), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n188), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n542), .A2(new_n356), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n533), .B2(new_n530), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n218), .B1(new_n520), .B2(new_n521), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n523), .A2(new_n233), .A3(new_n524), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT93), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT94), .A3(new_n529), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n538), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT94), .B1(new_n549), .B2(new_n529), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n539), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G475), .A2(G902), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT95), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n517), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n517), .A3(new_n555), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT96), .ZN(new_n558));
  INV_X1    g372(.A(new_n555), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n549), .A2(new_n529), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n538), .A3(new_n550), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n559), .B1(new_n563), .B2(new_n539), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n517), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n556), .B1(new_n558), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G475), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n535), .B(new_n538), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n568), .B1(new_n569), .B2(new_n333), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G478), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT102), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n190), .A2(G128), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n190), .B2(G128), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n225), .A2(KEYINPUT99), .A3(G143), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n579), .A2(new_n580), .B1(new_n575), .B2(new_n576), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n581), .B2(KEYINPUT100), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n580), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n575), .A2(new_n576), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n207), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n583), .A2(new_n207), .A3(new_n575), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n590));
  INV_X1    g404(.A(G122), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(G116), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n248), .A2(KEYINPUT98), .A3(G122), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(KEYINPUT97), .A2(G122), .ZN(new_n595));
  NOR2_X1   g409(.A1(KEYINPUT97), .A2(G122), .ZN(new_n596));
  OAI21_X1  g410(.A(G116), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n594), .A2(new_n597), .A3(new_n397), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n397), .B1(new_n594), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n589), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n594), .A2(new_n597), .A3(new_n397), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n583), .A2(new_n207), .A3(new_n575), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n207), .B1(new_n583), .B2(new_n575), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT97), .B(G122), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n594), .A2(KEYINPUT14), .B1(new_n605), .B2(G116), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT14), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n592), .A2(new_n607), .A3(new_n593), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n397), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI22_X1  g423(.A1(new_n588), .A2(new_n600), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n386), .A2(new_n332), .A3(G953), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n225), .A2(KEYINPUT99), .A3(G143), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT99), .B1(new_n225), .B2(G143), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n584), .B(KEYINPUT100), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n577), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n581), .A2(KEYINPUT100), .ZN(new_n619));
  OAI21_X1  g433(.A(G134), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n594), .A2(new_n597), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G107), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n602), .B1(new_n622), .B2(new_n601), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n248), .A2(KEYINPUT98), .A3(G122), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT98), .B1(new_n248), .B2(G122), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT14), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n597), .A3(new_n608), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G107), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n575), .B1(new_n614), .B2(new_n615), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G134), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n589), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(new_n601), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n624), .A2(KEYINPUT101), .A3(new_n633), .A4(new_n611), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n613), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n605), .A2(G116), .B1(new_n592), .B2(new_n593), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n631), .A2(new_n589), .B1(new_n397), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n620), .A2(new_n623), .B1(new_n637), .B2(new_n629), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT101), .B1(new_n638), .B2(new_n611), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n574), .B(new_n333), .C1(new_n635), .C2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n610), .B2(new_n612), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n634), .A3(new_n613), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n574), .B1(new_n644), .B2(new_n333), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n573), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n573), .B1(new_n644), .B2(new_n333), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n367), .A2(G952), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(G234), .B2(G237), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT21), .B(G898), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT103), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n333), .B(new_n367), .C1(G234), .C2(G237), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n571), .A2(new_n649), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n516), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n331), .A2(new_n384), .A3(new_n464), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G101), .ZN(G3));
  OAI211_X1 g475(.A(new_n657), .B(new_n465), .C1(new_n514), .C2(new_n515), .ZN(new_n662));
  INV_X1    g476(.A(new_n556), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n565), .B1(new_n564), .B2(new_n517), .ZN(new_n664));
  AND4_X1   g478(.A1(new_n565), .A2(new_n553), .A3(new_n517), .A4(new_n555), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n570), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n644), .A2(new_n333), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT102), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n572), .A3(new_n640), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT33), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n644), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n638), .A2(new_n611), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n613), .A3(KEYINPUT33), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n572), .A2(G902), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n673), .A2(KEYINPUT105), .A3(new_n675), .A4(new_n676), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n671), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n662), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n312), .A2(new_n306), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n312), .B2(G902), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g501(.A(KEYINPUT104), .B(G472), .C1(new_n312), .C2(G902), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n388), .B(new_n383), .C1(new_n454), .C2(new_n463), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n683), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT34), .B(G104), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G6));
  NAND2_X1  g507(.A1(new_n687), .A2(new_n688), .ZN(new_n694));
  INV_X1    g508(.A(new_n684), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n690), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n557), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n570), .B1(new_n698), .B2(new_n556), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n663), .A2(new_n697), .A3(new_n557), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n670), .A2(new_n640), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n647), .B1(new_n702), .B2(new_n573), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n662), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n696), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT35), .B(G107), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G9));
  INV_X1    g522(.A(new_n465), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n501), .A2(new_n513), .ZN(new_n710));
  INV_X1    g524(.A(new_n502), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n501), .A2(new_n502), .A3(new_n513), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n668), .A2(new_n703), .A3(new_n656), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n371), .A2(KEYINPUT36), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n365), .B(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n333), .A3(new_n377), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n376), .A2(new_n718), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n464), .A2(new_n714), .A3(new_n715), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n689), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT37), .B(G110), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G12));
  INV_X1    g537(.A(G900), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n651), .B1(new_n655), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n703), .A2(new_n699), .A3(new_n700), .A4(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n727), .B(new_n465), .C1(new_n515), .C2(new_n514), .ZN(new_n728));
  INV_X1    g542(.A(new_n388), .ZN(new_n729));
  AOI211_X1 g543(.A(G469), .B(G902), .C1(new_n435), .C2(new_n451), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n460), .A2(new_n461), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n450), .B1(new_n427), .B2(new_n456), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n453), .B1(new_n733), .B2(new_n333), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n729), .B(new_n719), .C1(new_n730), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n331), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G128), .ZN(G30));
  XOR2_X1   g552(.A(new_n725), .B(KEYINPUT39), .Z(new_n739));
  NAND2_X1  g553(.A1(new_n464), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT40), .ZN(new_n741));
  INV_X1    g555(.A(new_n330), .ZN(new_n742));
  INV_X1    g556(.A(G472), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n318), .A2(new_n326), .ZN(new_n744));
  AOI21_X1  g558(.A(G902), .B1(new_n290), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n313), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT78), .B1(new_n684), .B2(KEYINPUT32), .ZN(new_n747));
  OR3_X1    g561(.A1(new_n742), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n514), .A2(new_n515), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT38), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n649), .B1(new_n666), .B2(new_n667), .ZN(new_n752));
  INV_X1    g566(.A(new_n719), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n465), .ZN(new_n754));
  OR4_X1    g568(.A1(new_n741), .A2(new_n749), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G143), .ZN(G45));
  OAI211_X1 g570(.A(new_n681), .B(new_n726), .C1(new_n567), .C2(new_n570), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n735), .A2(new_n516), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n331), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G146), .ZN(G48));
  AOI21_X1  g574(.A(new_n453), .B1(new_n452), .B2(new_n333), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n730), .A3(new_n388), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n331), .A2(new_n683), .A3(new_n384), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT41), .B(G113), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G15));
  NAND2_X1  g579(.A1(new_n331), .A2(new_n384), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n705), .A3(new_n762), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G116), .ZN(G18));
  NAND2_X1  g583(.A1(new_n433), .A2(new_n434), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n458), .B1(new_n446), .B2(KEYINPUT87), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n449), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n772), .B2(G902), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n729), .A3(new_n454), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n516), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n658), .A2(new_n753), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n331), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G119), .ZN(G21));
  OAI211_X1 g592(.A(new_n752), .B(new_n465), .C1(new_n514), .C2(new_n515), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n292), .A2(new_n293), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT28), .B1(new_n295), .B2(new_n316), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT76), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n320), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n287), .B1(new_n784), .B2(new_n314), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n307), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n786), .A2(new_n685), .A3(new_n384), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n780), .A2(new_n787), .A3(new_n762), .A4(new_n657), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT107), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n774), .A2(new_n656), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(KEYINPUT107), .A3(new_n787), .A4(new_n780), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G122), .ZN(G24));
  INV_X1    g608(.A(new_n757), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n786), .A2(new_n685), .A3(new_n719), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n775), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G125), .ZN(G27));
  NAND2_X1  g612(.A1(new_n322), .A2(KEYINPUT29), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n325), .A2(new_n327), .ZN(new_n800));
  AOI21_X1  g614(.A(G902), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n308), .B(new_n313), .C1(new_n801), .C2(new_n743), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n384), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n464), .A2(new_n750), .A3(new_n795), .A4(new_n465), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT42), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n729), .B1(new_n730), .B2(new_n734), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n712), .A2(new_n465), .A3(new_n713), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n757), .A2(KEYINPUT42), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n331), .A2(new_n808), .A3(new_n384), .A4(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G131), .ZN(G33));
  NAND3_X1  g626(.A1(new_n767), .A2(new_n727), .A3(new_n808), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G134), .ZN(G36));
  XNOR2_X1  g628(.A(new_n733), .B(KEYINPUT45), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(G469), .ZN(new_n816));
  NAND2_X1  g630(.A1(G469), .A2(G902), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n816), .A2(KEYINPUT46), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT46), .B1(new_n816), .B2(new_n817), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n818), .A2(new_n819), .A3(new_n730), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n820), .A2(new_n729), .A3(new_n739), .ZN(new_n821));
  INV_X1    g635(.A(new_n689), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n571), .A2(new_n681), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT43), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n825), .A3(new_n719), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT44), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n807), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n821), .B(new_n828), .C1(new_n827), .C2(new_n826), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G137), .ZN(G39));
  NOR4_X1   g644(.A1(new_n331), .A2(new_n384), .A3(new_n757), .A4(new_n807), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT108), .Z(new_n832));
  AND3_X1   g646(.A1(new_n820), .A2(KEYINPUT47), .A3(new_n729), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT47), .B1(new_n820), .B2(new_n729), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G140), .ZN(G42));
  NOR2_X1   g650(.A1(new_n761), .A2(new_n730), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n388), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n833), .A2(new_n834), .A3(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n825), .A2(new_n651), .A3(new_n787), .ZN(new_n841));
  INV_X1    g655(.A(new_n807), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT116), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT51), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n841), .A2(new_n709), .A3(new_n751), .A4(new_n762), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(KEYINPUT118), .A3(KEYINPUT50), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n651), .A2(new_n825), .A3(new_n762), .A4(new_n842), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n796), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n762), .A2(new_n842), .A3(new_n384), .A4(new_n651), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n748), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n668), .A2(new_n681), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n849), .A2(new_n850), .A3(new_n852), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT119), .B1(new_n845), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n843), .B(KEYINPUT116), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n820), .A2(new_n729), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT47), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n820), .A2(KEYINPUT47), .A3(new_n729), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(new_n838), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n859), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n849), .A2(new_n852), .A3(new_n856), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n850), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n858), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT117), .B1(new_n833), .B2(new_n834), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n863), .A2(new_n872), .A3(new_n864), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n844), .B1(new_n874), .B2(new_n838), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n859), .B1(new_n875), .B2(new_n857), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n851), .A2(new_n384), .A3(new_n802), .ZN(new_n877));
  XOR2_X1   g691(.A(KEYINPUT120), .B(KEYINPUT48), .Z(new_n878));
  XNOR2_X1  g692(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n682), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n854), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n650), .B1(new_n841), .B2(new_n775), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n870), .A2(new_n876), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n870), .A2(new_n876), .A3(KEYINPUT121), .A4(new_n883), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n649), .A2(KEYINPUT111), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n649), .A2(KEYINPUT111), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(new_n701), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n786), .A2(new_n685), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n331), .A2(new_n892), .B1(new_n880), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n808), .A2(new_n719), .A3(new_n726), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n813), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT113), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT112), .B1(new_n891), .B2(new_n668), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT112), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n899), .B(new_n571), .C1(new_n889), .C2(new_n890), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n662), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n696), .A2(new_n901), .B1(new_n720), .B2(new_n689), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT110), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n660), .A2(new_n903), .A3(new_n691), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n660), .B2(new_n691), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n660), .A2(new_n691), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT110), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(KEYINPUT113), .A3(new_n904), .A4(new_n902), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n896), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n779), .A2(new_n806), .A3(new_n719), .A4(new_n725), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n748), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n759), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT52), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n737), .A2(new_n797), .ZN(new_n916));
  OR3_X1    g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n914), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n763), .A2(new_n777), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n811), .A2(new_n920), .A3(new_n768), .A4(new_n793), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n911), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n915), .B1(new_n912), .B2(new_n748), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n737), .A2(KEYINPUT114), .A3(new_n797), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT114), .B1(new_n737), .B2(new_n797), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n759), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n924), .B1(new_n930), .B2(new_n918), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n921), .A2(KEYINPUT115), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n921), .A2(KEYINPUT115), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n911), .A2(new_n931), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n925), .A2(new_n926), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n923), .A2(KEYINPUT53), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n896), .B(new_n921), .C1(new_n907), .C2(new_n910), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT53), .B1(new_n930), .B2(new_n918), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n935), .B1(new_n940), .B2(new_n926), .ZN(new_n941));
  OAI22_X1  g755(.A1(new_n888), .A2(new_n941), .B1(G952), .B2(G953), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n837), .B(KEYINPUT49), .ZN(new_n943));
  NOR4_X1   g757(.A1(new_n823), .A2(new_n383), .A3(new_n388), .A4(new_n709), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n749), .A2(new_n751), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT109), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n942), .A2(new_n946), .ZN(G75));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n925), .A2(new_n934), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(G902), .ZN(new_n950));
  INV_X1    g764(.A(G210), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n480), .B1(new_n496), .B2(new_n500), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(new_n486), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT55), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n952), .A2(new_n956), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n367), .A2(G952), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G51));
  NOR2_X1   g774(.A1(new_n950), .A2(new_n816), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT53), .B1(new_n937), .B2(new_n919), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n911), .A2(new_n931), .A3(new_n932), .A4(new_n933), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT54), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n935), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n817), .B(KEYINPUT57), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n772), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n968), .B2(KEYINPUT122), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT122), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n964), .B2(new_n935), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n772), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n959), .B1(new_n969), .B2(new_n972), .ZN(G54));
  NAND4_X1  g787(.A1(new_n949), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n974));
  INV_X1    g788(.A(new_n553), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n959), .ZN(G60));
  AND2_X1   g792(.A1(new_n673), .A2(new_n675), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT59), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n941), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n979), .A2(new_n981), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n959), .B(new_n982), .C1(new_n965), .C2(new_n983), .ZN(G63));
  XNOR2_X1  g798(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n332), .A2(new_n333), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n962), .B2(new_n963), .ZN(new_n988));
  INV_X1    g802(.A(new_n373), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n959), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n717), .B(new_n987), .C1(new_n962), .C2(new_n963), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n992), .A2(KEYINPUT124), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT124), .ZN(new_n994));
  INV_X1    g808(.A(new_n987), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n925), .B2(new_n934), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n996), .B2(new_n717), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n990), .B(new_n991), .C1(new_n993), .C2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n992), .A2(KEYINPUT124), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n996), .A2(new_n994), .A3(new_n717), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n991), .B1(new_n1002), .B2(new_n990), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n999), .A2(new_n1003), .ZN(G66));
  OAI21_X1  g818(.A(G953), .B1(new_n654), .B2(new_n484), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n907), .A2(new_n910), .ZN(new_n1006));
  AND4_X1   g820(.A1(new_n768), .A2(new_n1006), .A3(new_n793), .A4(new_n920), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n953), .B1(G898), .B2(new_n367), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(G69));
  NAND3_X1  g824(.A1(new_n246), .A2(new_n274), .A3(new_n281), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n540), .A2(new_n541), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1011), .B(new_n1012), .Z(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n928), .A2(new_n929), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n331), .B2(new_n758), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n755), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT62), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n898), .A2(new_n900), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n740), .B(new_n807), .C1(new_n1020), .C2(new_n682), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n767), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n835), .A2(new_n829), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1014), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n821), .A2(new_n384), .A3(new_n780), .A4(new_n802), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n835), .A2(new_n811), .A3(new_n813), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n829), .A2(new_n1016), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT126), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n829), .A2(new_n1016), .A3(KEYINPUT126), .ZN(new_n1030));
  AOI211_X1 g844(.A(new_n1013), .B(new_n1026), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n367), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(G953), .B1(new_n390), .B2(new_n724), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT127), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n1013), .A2(new_n724), .A3(new_n367), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1036), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1035), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  NAND2_X1  g854(.A1(new_n282), .A2(new_n289), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n287), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1019), .A2(new_n1007), .A3(new_n1023), .ZN(new_n1043));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  AOI21_X1  g859(.A(new_n1042), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1041), .A2(new_n287), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1026), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n1007), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1048), .B1(new_n1050), .B2(new_n1045), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1048), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n940), .A2(new_n1052), .ZN(new_n1053));
  NOR4_X1   g867(.A1(new_n1046), .A2(new_n1051), .A3(new_n959), .A4(new_n1053), .ZN(G57));
endmodule


