

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747;

  AND2_X1 U365 ( .A1(n379), .A2(n391), .ZN(n390) );
  XNOR2_X1 U366 ( .A(n378), .B(n725), .ZN(n469) );
  XNOR2_X1 U367 ( .A(n443), .B(KEYINPUT71), .ZN(n378) );
  XOR2_X1 U368 ( .A(KEYINPUT70), .B(G140), .Z(n435) );
  XNOR2_X1 U369 ( .A(KEYINPUT3), .B(G116), .ZN(n447) );
  XNOR2_X2 U370 ( .A(n595), .B(n407), .ZN(n585) );
  XNOR2_X2 U371 ( .A(n393), .B(n502), .ZN(n733) );
  XNOR2_X2 U372 ( .A(n381), .B(n455), .ZN(n703) );
  NOR2_X2 U373 ( .A1(n534), .A2(n533), .ZN(n535) );
  INV_X2 U374 ( .A(G146), .ZN(n434) );
  NAND2_X4 U375 ( .A1(n390), .A2(n387), .ZN(n375) );
  NAND2_X1 U376 ( .A1(n613), .A2(n616), .ZN(n670) );
  XNOR2_X1 U377 ( .A(n355), .B(KEYINPUT40), .ZN(n746) );
  NAND2_X1 U378 ( .A1(n576), .A2(n575), .ZN(n589) );
  XNOR2_X1 U379 ( .A(n401), .B(n453), .ZN(n580) );
  XNOR2_X1 U380 ( .A(n431), .B(n430), .ZN(n549) );
  XNOR2_X1 U381 ( .A(n403), .B(n402), .ZN(n503) );
  XNOR2_X1 U382 ( .A(n447), .B(G113), .ZN(n468) );
  XNOR2_X1 U383 ( .A(n395), .B(G131), .ZN(n485) );
  INV_X2 U384 ( .A(KEYINPUT68), .ZN(n354) );
  XNOR2_X1 U385 ( .A(G143), .B(G128), .ZN(n458) );
  INV_X2 U386 ( .A(G953), .ZN(n456) );
  AND2_X2 U387 ( .A1(n672), .A2(n416), .ZN(n346) );
  AND2_X2 U388 ( .A1(n672), .A2(n416), .ZN(n711) );
  AND2_X1 U389 ( .A1(n582), .A2(n375), .ZN(n586) );
  NAND2_X1 U390 ( .A1(n674), .A2(n675), .ZN(n442) );
  NOR2_X2 U391 ( .A1(n703), .A2(n517), .ZN(n380) );
  XNOR2_X2 U392 ( .A(n733), .B(n434), .ZN(n376) );
  XNOR2_X1 U393 ( .A(n406), .B(n405), .ZN(n404) );
  INV_X1 U394 ( .A(KEYINPUT74), .ZN(n405) );
  NAND2_X1 U395 ( .A1(n368), .A2(n365), .ZN(n406) );
  AND2_X1 U396 ( .A1(n367), .A2(n366), .ZN(n365) );
  NOR2_X1 U397 ( .A1(n400), .A2(n397), .ZN(n581) );
  NOR2_X1 U398 ( .A1(n657), .A2(n369), .ZN(n368) );
  NAND2_X1 U399 ( .A1(n371), .A2(n374), .ZN(n370) );
  AND2_X1 U400 ( .A1(n634), .A2(n410), .ZN(n551) );
  NAND2_X1 U401 ( .A1(n364), .A2(n348), .ZN(n363) );
  NOR2_X1 U402 ( .A1(n746), .A2(n745), .ZN(n584) );
  INV_X1 U403 ( .A(n485), .ZN(n394) );
  XOR2_X1 U404 ( .A(KEYINPUT12), .B(G122), .Z(n493) );
  XNOR2_X1 U405 ( .A(KEYINPUT102), .B(KEYINPUT11), .ZN(n488) );
  NAND2_X1 U406 ( .A1(n620), .A2(n471), .ZN(n401) );
  XNOR2_X1 U407 ( .A(n464), .B(n463), .ZN(n382) );
  XNOR2_X1 U408 ( .A(n469), .B(n727), .ZN(n383) );
  XNOR2_X1 U409 ( .A(n578), .B(KEYINPUT41), .ZN(n704) );
  INV_X1 U410 ( .A(n589), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n497), .B(n498), .ZN(n528) );
  NAND2_X1 U412 ( .A1(n389), .A2(n471), .ZN(n388) );
  NAND2_X1 U413 ( .A1(n693), .A2(KEYINPUT47), .ZN(n366) );
  INV_X1 U414 ( .A(n667), .ZN(n600) );
  INV_X1 U415 ( .A(KEYINPUT69), .ZN(n395) );
  INV_X1 U416 ( .A(KEYINPUT8), .ZN(n402) );
  NAND2_X1 U417 ( .A1(n456), .A2(G234), .ZN(n403) );
  XNOR2_X1 U418 ( .A(n434), .B(G125), .ZN(n462) );
  XOR2_X1 U419 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n459) );
  XOR2_X1 U420 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n479) );
  AND2_X1 U421 ( .A1(n375), .A2(n570), .ZN(n572) );
  NAND2_X1 U422 ( .A1(n398), .A2(n549), .ZN(n397) );
  NOR2_X1 U423 ( .A1(n579), .A2(n399), .ZN(n398) );
  INV_X1 U424 ( .A(n679), .ZN(n399) );
  INV_X1 U425 ( .A(G469), .ZN(n389) );
  NAND2_X1 U426 ( .A1(G902), .A2(G469), .ZN(n391) );
  NOR2_X1 U427 ( .A1(n549), .A2(n531), .ZN(n569) );
  XNOR2_X1 U428 ( .A(G137), .B(G128), .ZN(n417) );
  XOR2_X1 U429 ( .A(KEYINPUT23), .B(KEYINPUT98), .Z(n418) );
  INV_X1 U430 ( .A(G134), .ZN(n392) );
  XOR2_X1 U431 ( .A(KEYINPUT7), .B(G122), .Z(n500) );
  XNOR2_X1 U432 ( .A(n494), .B(n412), .ZN(n495) );
  XNOR2_X1 U433 ( .A(n380), .B(KEYINPUT34), .ZN(n512) );
  XNOR2_X1 U434 ( .A(n534), .B(KEYINPUT96), .ZN(n517) );
  XNOR2_X1 U435 ( .A(KEYINPUT16), .B(G122), .ZN(n465) );
  NOR2_X1 U436 ( .A1(n704), .A2(n360), .ZN(n583) );
  AND2_X1 U437 ( .A1(n609), .A2(n661), .ZN(n355) );
  XNOR2_X1 U438 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n520) );
  AND2_X1 U439 ( .A1(n373), .A2(n372), .ZN(n657) );
  INV_X1 U440 ( .A(n591), .ZN(n372) );
  NAND2_X1 U441 ( .A1(n409), .A2(n549), .ZN(n634) );
  INV_X1 U442 ( .A(KEYINPUT66), .ZN(n411) );
  XNOR2_X1 U443 ( .A(KEYINPUT106), .B(n539), .ZN(n747) );
  AND2_X1 U444 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U445 ( .A(n384), .B(KEYINPUT85), .ZN(n538) );
  XNOR2_X1 U446 ( .A(n713), .B(n712), .ZN(n714) );
  AND2_X1 U447 ( .A1(n357), .A2(n358), .ZN(n347) );
  AND2_X1 U448 ( .A1(n404), .A2(n600), .ZN(n348) );
  AND2_X1 U449 ( .A1(n359), .A2(n358), .ZN(n349) );
  XOR2_X1 U450 ( .A(n606), .B(KEYINPUT38), .Z(n350) );
  AND2_X1 U451 ( .A1(n536), .A2(n602), .ZN(n351) );
  XNOR2_X1 U452 ( .A(n383), .B(n382), .ZN(n637) );
  XNOR2_X1 U453 ( .A(n645), .B(KEYINPUT59), .ZN(n352) );
  XNOR2_X1 U454 ( .A(KEYINPUT119), .B(n635), .ZN(n353) );
  INV_X1 U455 ( .A(KEYINPUT47), .ZN(n374) );
  INV_X1 U456 ( .A(n717), .ZN(n358) );
  XNOR2_X1 U457 ( .A(n535), .B(KEYINPUT22), .ZN(n542) );
  INV_X1 U458 ( .A(n528), .ZN(n529) );
  NOR2_X1 U459 ( .A1(n744), .A2(KEYINPUT65), .ZN(n410) );
  XNOR2_X1 U460 ( .A(n496), .B(n495), .ZN(n645) );
  XNOR2_X1 U461 ( .A(n487), .B(n488), .ZN(n489) );
  XNOR2_X2 U462 ( .A(n354), .B(G101), .ZN(n443) );
  XNOR2_X1 U463 ( .A(n584), .B(KEYINPUT46), .ZN(n364) );
  NAND2_X1 U464 ( .A1(n356), .A2(n350), .ZN(n577) );
  XNOR2_X1 U465 ( .A(n413), .B(n419), .ZN(n423) );
  XNOR2_X1 U466 ( .A(n646), .B(n352), .ZN(n357) );
  XNOR2_X1 U467 ( .A(n636), .B(n353), .ZN(n359) );
  NAND2_X1 U468 ( .A1(n628), .A2(G469), .ZN(n379) );
  XNOR2_X2 U469 ( .A(n376), .B(n439), .ZN(n628) );
  INV_X1 U470 ( .A(n586), .ZN(n360) );
  NAND2_X1 U471 ( .A1(n361), .A2(n611), .ZN(n734) );
  XNOR2_X1 U472 ( .A(n363), .B(n362), .ZN(n361) );
  INV_X1 U473 ( .A(KEYINPUT48), .ZN(n362) );
  XNOR2_X1 U474 ( .A(n590), .B(KEYINPUT110), .ZN(n373) );
  NAND2_X1 U475 ( .A1(n659), .A2(KEYINPUT47), .ZN(n367) );
  NOR2_X1 U476 ( .A1(n659), .A2(n370), .ZN(n369) );
  INV_X1 U477 ( .A(n693), .ZN(n371) );
  XNOR2_X2 U478 ( .A(n587), .B(KEYINPUT82), .ZN(n659) );
  NAND2_X1 U479 ( .A1(n675), .A2(n375), .ZN(n516) );
  XNOR2_X2 U480 ( .A(n375), .B(n441), .ZN(n674) );
  XNOR2_X1 U481 ( .A(n376), .B(n451), .ZN(n620) );
  XNOR2_X2 U482 ( .A(n377), .B(KEYINPUT0), .ZN(n534) );
  NAND2_X1 U483 ( .A1(n585), .A2(n414), .ZN(n377) );
  XNOR2_X2 U484 ( .A(n408), .B(n477), .ZN(n595) );
  NAND2_X1 U485 ( .A1(n519), .A2(n593), .ZN(n381) );
  AND2_X1 U486 ( .A1(n542), .A2(n602), .ZN(n547) );
  NAND2_X1 U487 ( .A1(n542), .A2(n351), .ZN(n384) );
  NAND2_X1 U488 ( .A1(n560), .A2(n559), .ZN(n561) );
  OR2_X2 U489 ( .A1(n385), .A2(n541), .ZN(n527) );
  NAND2_X1 U490 ( .A1(n385), .A2(n541), .ZN(n552) );
  XNOR2_X1 U491 ( .A(n385), .B(n742), .ZN(G24) );
  XNOR2_X2 U492 ( .A(n514), .B(n513), .ZN(n385) );
  NAND2_X1 U493 ( .A1(n386), .A2(n617), .ZN(n618) );
  XNOR2_X2 U494 ( .A(n561), .B(KEYINPUT45), .ZN(n386) );
  NAND2_X1 U495 ( .A1(n386), .A2(n612), .ZN(n613) );
  NAND2_X1 U496 ( .A1(n386), .A2(n456), .ZN(n721) );
  OR2_X1 U497 ( .A1(n628), .A2(n388), .ZN(n387) );
  XNOR2_X1 U498 ( .A(n458), .B(n392), .ZN(n502) );
  XNOR2_X1 U499 ( .A(n396), .B(n394), .ZN(n393) );
  XNOR2_X1 U500 ( .A(n461), .B(G137), .ZN(n396) );
  XNOR2_X2 U501 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n461) );
  INV_X1 U502 ( .A(n549), .ZN(n537) );
  INV_X1 U503 ( .A(n397), .ZN(n592) );
  INV_X1 U504 ( .A(n580), .ZN(n400) );
  INV_X1 U505 ( .A(KEYINPUT19), .ZN(n407) );
  NAND2_X2 U506 ( .A1(n562), .A2(n689), .ZN(n408) );
  XNOR2_X1 U507 ( .A(n548), .B(n411), .ZN(n409) );
  NAND2_X1 U508 ( .A1(n634), .A2(n550), .ZN(n556) );
  NOR2_X1 U509 ( .A1(n734), .A2(n616), .ZN(n617) );
  AND2_X2 U510 ( .A1(n670), .A2(n615), .ZN(n416) );
  XOR2_X1 U511 ( .A(n493), .B(n492), .Z(n412) );
  XOR2_X1 U512 ( .A(n418), .B(n417), .Z(n413) );
  XOR2_X1 U513 ( .A(n484), .B(KEYINPUT95), .Z(n414) );
  NOR2_X1 U514 ( .A1(n526), .A2(n525), .ZN(n415) );
  BUF_X1 U515 ( .A(n569), .Z(n675) );
  XNOR2_X1 U516 ( .A(n423), .B(n422), .ZN(n425) );
  BUF_X1 U517 ( .A(n562), .Z(n606) );
  XNOR2_X1 U518 ( .A(n521), .B(n520), .ZN(n665) );
  XNOR2_X1 U519 ( .A(n715), .B(n714), .ZN(n716) );
  XOR2_X1 U520 ( .A(KEYINPUT88), .B(KEYINPUT33), .Z(n455) );
  NAND2_X1 U521 ( .A1(G221), .A2(n503), .ZN(n419) );
  XNOR2_X2 U522 ( .A(G119), .B(G110), .ZN(n466) );
  XOR2_X1 U523 ( .A(KEYINPUT24), .B(n466), .Z(n421) );
  XOR2_X1 U524 ( .A(KEYINPUT80), .B(KEYINPUT97), .Z(n420) );
  XNOR2_X1 U525 ( .A(n421), .B(n420), .ZN(n422) );
  INV_X1 U526 ( .A(n462), .ZN(n424) );
  XNOR2_X1 U527 ( .A(KEYINPUT10), .B(n424), .ZN(n487) );
  XNOR2_X1 U528 ( .A(n487), .B(n435), .ZN(n732) );
  XNOR2_X1 U529 ( .A(n425), .B(n732), .ZN(n713) );
  NOR2_X1 U530 ( .A1(G902), .A2(n713), .ZN(n431) );
  XOR2_X1 U531 ( .A(KEYINPUT99), .B(KEYINPUT20), .Z(n427) );
  XNOR2_X1 U532 ( .A(G902), .B(KEYINPUT15), .ZN(n614) );
  NAND2_X1 U533 ( .A1(G234), .A2(n614), .ZN(n426) );
  XNOR2_X1 U534 ( .A(n427), .B(n426), .ZN(n432) );
  NAND2_X1 U535 ( .A1(G217), .A2(n432), .ZN(n429) );
  INV_X1 U536 ( .A(KEYINPUT25), .ZN(n428) );
  XNOR2_X1 U537 ( .A(n429), .B(n428), .ZN(n430) );
  NAND2_X1 U538 ( .A1(n432), .A2(G221), .ZN(n433) );
  XOR2_X1 U539 ( .A(KEYINPUT21), .B(n433), .Z(n679) );
  XOR2_X1 U540 ( .A(n679), .B(KEYINPUT100), .Z(n531) );
  XOR2_X1 U541 ( .A(G107), .B(G104), .Z(n725) );
  XOR2_X1 U542 ( .A(G110), .B(n435), .Z(n437) );
  NAND2_X1 U543 ( .A1(G227), .A2(n456), .ZN(n436) );
  XOR2_X1 U544 ( .A(n437), .B(n436), .Z(n438) );
  XNOR2_X1 U545 ( .A(n469), .B(n438), .ZN(n439) );
  INV_X1 U546 ( .A(KEYINPUT67), .ZN(n440) );
  XNOR2_X1 U547 ( .A(n440), .B(KEYINPUT1), .ZN(n441) );
  XNOR2_X2 U548 ( .A(n442), .B(KEYINPUT75), .ZN(n519) );
  XOR2_X1 U549 ( .A(KEYINPUT5), .B(n443), .Z(n446) );
  NOR2_X1 U550 ( .A1(G953), .A2(G237), .ZN(n444) );
  XOR2_X1 U551 ( .A(KEYINPUT77), .B(n444), .Z(n491) );
  NAND2_X1 U552 ( .A1(G210), .A2(n491), .ZN(n445) );
  XNOR2_X1 U553 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U554 ( .A(G119), .B(KEYINPUT76), .ZN(n448) );
  XNOR2_X1 U555 ( .A(n468), .B(n448), .ZN(n449) );
  XNOR2_X1 U556 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U557 ( .A(G902), .ZN(n471) );
  INV_X1 U558 ( .A(KEYINPUT73), .ZN(n452) );
  XNOR2_X1 U559 ( .A(n452), .B(G472), .ZN(n453) );
  INV_X1 U560 ( .A(KEYINPUT6), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n580), .B(n454), .ZN(n593) );
  NAND2_X1 U562 ( .A1(G224), .A2(n456), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U564 ( .A(n460), .B(n459), .ZN(n464) );
  XNOR2_X1 U565 ( .A(n461), .B(n462), .ZN(n463) );
  XNOR2_X1 U566 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n467), .B(n468), .ZN(n727) );
  NAND2_X1 U568 ( .A1(n637), .A2(n614), .ZN(n474) );
  INV_X1 U569 ( .A(G237), .ZN(n470) );
  NAND2_X1 U570 ( .A1(n471), .A2(n470), .ZN(n475) );
  NAND2_X1 U571 ( .A1(n475), .A2(G210), .ZN(n472) );
  XNOR2_X1 U572 ( .A(n472), .B(KEYINPUT89), .ZN(n473) );
  XNOR2_X2 U573 ( .A(n474), .B(n473), .ZN(n562) );
  NAND2_X1 U574 ( .A1(n475), .A2(G214), .ZN(n476) );
  XNOR2_X1 U575 ( .A(n476), .B(KEYINPUT90), .ZN(n689) );
  INV_X1 U576 ( .A(KEYINPUT86), .ZN(n477) );
  NAND2_X1 U577 ( .A1(G234), .A2(G237), .ZN(n478) );
  XNOR2_X1 U578 ( .A(n479), .B(n478), .ZN(n481) );
  NAND2_X1 U579 ( .A1(n481), .A2(G952), .ZN(n480) );
  XNOR2_X1 U580 ( .A(n480), .B(KEYINPUT92), .ZN(n701) );
  NOR2_X1 U581 ( .A1(G953), .A2(n701), .ZN(n567) );
  NAND2_X1 U582 ( .A1(n481), .A2(G902), .ZN(n482) );
  XNOR2_X1 U583 ( .A(KEYINPUT94), .B(n482), .ZN(n563) );
  XNOR2_X1 U584 ( .A(G898), .B(KEYINPUT93), .ZN(n720) );
  NAND2_X1 U585 ( .A1(G953), .A2(n720), .ZN(n728) );
  NOR2_X1 U586 ( .A1(n563), .A2(n728), .ZN(n483) );
  OR2_X1 U587 ( .A1(n567), .A2(n483), .ZN(n484) );
  XNOR2_X1 U588 ( .A(KEYINPUT13), .B(G475), .ZN(n498) );
  XNOR2_X1 U589 ( .A(G143), .B(n485), .ZN(n486) );
  XNOR2_X1 U590 ( .A(n486), .B(G140), .ZN(n490) );
  XNOR2_X1 U591 ( .A(n490), .B(n489), .ZN(n496) );
  AND2_X1 U592 ( .A1(G214), .A2(n491), .ZN(n494) );
  XNOR2_X1 U593 ( .A(G113), .B(G104), .ZN(n492) );
  NOR2_X1 U594 ( .A1(G902), .A2(n645), .ZN(n497) );
  XNOR2_X1 U595 ( .A(G116), .B(G107), .ZN(n499) );
  XNOR2_X1 U596 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U597 ( .A(n502), .B(n501), .ZN(n507) );
  NAND2_X1 U598 ( .A1(G217), .A2(n503), .ZN(n505) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n504) );
  XNOR2_X1 U600 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U601 ( .A(n507), .B(n506), .ZN(n635) );
  NOR2_X1 U602 ( .A1(G902), .A2(n635), .ZN(n509) );
  XNOR2_X1 U603 ( .A(KEYINPUT104), .B(G478), .ZN(n508) );
  XNOR2_X1 U604 ( .A(n509), .B(n508), .ZN(n530) );
  INV_X1 U605 ( .A(n530), .ZN(n510) );
  NAND2_X1 U606 ( .A1(n528), .A2(n510), .ZN(n591) );
  XNOR2_X1 U607 ( .A(n591), .B(KEYINPUT81), .ZN(n511) );
  NAND2_X1 U608 ( .A1(n512), .A2(n511), .ZN(n514) );
  INV_X1 U609 ( .A(KEYINPUT35), .ZN(n513) );
  INV_X1 U610 ( .A(KEYINPUT44), .ZN(n515) );
  AND2_X1 U611 ( .A1(n515), .A2(KEYINPUT72), .ZN(n541) );
  NAND2_X1 U612 ( .A1(n528), .A2(n530), .ZN(n658) );
  INV_X1 U613 ( .A(n658), .ZN(n661) );
  NOR2_X1 U614 ( .A1(n528), .A2(n530), .ZN(n664) );
  NOR2_X1 U615 ( .A1(n661), .A2(n664), .ZN(n693) );
  INV_X1 U616 ( .A(n400), .ZN(n678) );
  OR2_X1 U617 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U618 ( .A1(n678), .A2(n518), .ZN(n649) );
  NAND2_X1 U619 ( .A1(n519), .A2(n678), .ZN(n683) );
  NOR2_X1 U620 ( .A1(n683), .A2(n534), .ZN(n521) );
  NOR2_X1 U621 ( .A1(n649), .A2(n665), .ZN(n522) );
  NOR2_X1 U622 ( .A1(n693), .A2(n522), .ZN(n526) );
  NOR2_X1 U623 ( .A1(KEYINPUT44), .A2(KEYINPUT65), .ZN(n524) );
  AND2_X1 U624 ( .A1(KEYINPUT72), .A2(KEYINPUT44), .ZN(n523) );
  NOR2_X1 U625 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U626 ( .A1(n527), .A2(n415), .ZN(n540) );
  NAND2_X1 U627 ( .A1(n530), .A2(n529), .ZN(n691) );
  NOR2_X1 U628 ( .A1(n691), .A2(n531), .ZN(n532) );
  XNOR2_X1 U629 ( .A(n532), .B(KEYINPUT105), .ZN(n533) );
  INV_X1 U630 ( .A(n674), .ZN(n602) );
  INV_X1 U631 ( .A(n593), .ZN(n536) );
  NOR2_X1 U632 ( .A1(n540), .A2(n747), .ZN(n560) );
  NAND2_X1 U633 ( .A1(n674), .A2(n549), .ZN(n543) );
  NOR2_X1 U634 ( .A1(n543), .A2(n593), .ZN(n544) );
  NAND2_X1 U635 ( .A1(n542), .A2(n544), .ZN(n546) );
  INV_X1 U636 ( .A(KEYINPUT32), .ZN(n545) );
  XNOR2_X1 U637 ( .A(n546), .B(n545), .ZN(n744) );
  INV_X1 U638 ( .A(n744), .ZN(n550) );
  NAND2_X1 U639 ( .A1(n547), .A2(n400), .ZN(n548) );
  NAND2_X1 U640 ( .A1(n552), .A2(n551), .ZN(n558) );
  INV_X1 U641 ( .A(KEYINPUT65), .ZN(n553) );
  NAND2_X1 U642 ( .A1(n553), .A2(KEYINPUT44), .ZN(n554) );
  AND2_X1 U643 ( .A1(n554), .A2(KEYINPUT72), .ZN(n555) );
  NAND2_X1 U644 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U645 ( .A1(n558), .A2(n557), .ZN(n559) );
  OR2_X1 U646 ( .A1(n456), .A2(n563), .ZN(n564) );
  XOR2_X1 U647 ( .A(KEYINPUT107), .B(n564), .Z(n565) );
  NOR2_X1 U648 ( .A1(G900), .A2(n565), .ZN(n566) );
  NOR2_X1 U649 ( .A1(n567), .A2(n566), .ZN(n579) );
  INV_X1 U650 ( .A(n579), .ZN(n568) );
  AND2_X1 U651 ( .A1(n569), .A2(n568), .ZN(n570) );
  INV_X1 U652 ( .A(KEYINPUT79), .ZN(n571) );
  XNOR2_X1 U653 ( .A(n572), .B(n571), .ZN(n576) );
  NAND2_X1 U654 ( .A1(n689), .A2(n580), .ZN(n574) );
  XNOR2_X1 U655 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n573) );
  XNOR2_X1 U656 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U657 ( .A(n577), .B(KEYINPUT39), .ZN(n609) );
  NAND2_X1 U658 ( .A1(n350), .A2(n689), .ZN(n692) );
  NOR2_X1 U659 ( .A1(n692), .A2(n691), .ZN(n578) );
  XNOR2_X1 U660 ( .A(n581), .B(KEYINPUT28), .ZN(n582) );
  XNOR2_X1 U661 ( .A(n583), .B(KEYINPUT42), .ZN(n745) );
  NAND2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U663 ( .A(n606), .ZN(n588) );
  NOR2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n658), .A2(n594), .ZN(n601) );
  INV_X1 U667 ( .A(n601), .ZN(n597) );
  INV_X1 U668 ( .A(n595), .ZN(n596) );
  NOR2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U670 ( .A(KEYINPUT36), .B(n598), .Z(n599) );
  NOR2_X1 U671 ( .A1(n602), .A2(n599), .ZN(n667) );
  INV_X1 U672 ( .A(n689), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n605), .B(KEYINPUT43), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U677 ( .A(n608), .B(KEYINPUT108), .ZN(n743) );
  NAND2_X1 U678 ( .A1(n664), .A2(n609), .ZN(n669) );
  INV_X1 U679 ( .A(n669), .ZN(n610) );
  NOR2_X1 U680 ( .A1(n743), .A2(n610), .ZN(n611) );
  INV_X1 U681 ( .A(n734), .ZN(n612) );
  INV_X1 U682 ( .A(KEYINPUT2), .ZN(n616) );
  INV_X1 U683 ( .A(n614), .ZN(n615) );
  XNOR2_X2 U684 ( .A(n618), .B(KEYINPUT78), .ZN(n672) );
  NAND2_X1 U685 ( .A1(n711), .A2(G472), .ZN(n622) );
  XNOR2_X1 U686 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n619) );
  XNOR2_X1 U687 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U688 ( .A(n622), .B(n621), .ZN(n623) );
  INV_X1 U689 ( .A(n623), .ZN(n625) );
  INV_X1 U690 ( .A(G952), .ZN(n624) );
  AND2_X1 U691 ( .A1(n624), .A2(G953), .ZN(n717) );
  NAND2_X1 U692 ( .A1(n625), .A2(n358), .ZN(n626) );
  XNOR2_X1 U693 ( .A(n626), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U694 ( .A1(n346), .A2(G469), .ZN(n630) );
  XOR2_X1 U695 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n627) );
  XNOR2_X1 U696 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U698 ( .A1(n631), .A2(n717), .ZN(n633) );
  INV_X1 U699 ( .A(KEYINPUT117), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n633), .B(n632), .ZN(G54) );
  XNOR2_X1 U701 ( .A(n634), .B(G110), .ZN(G12) );
  NAND2_X1 U702 ( .A1(n711), .A2(G478), .ZN(n636) );
  XNOR2_X1 U703 ( .A(n349), .B(KEYINPUT120), .ZN(G63) );
  NAND2_X1 U704 ( .A1(n346), .A2(G210), .ZN(n641) );
  XNOR2_X1 U705 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n638) );
  XOR2_X1 U706 ( .A(n638), .B(KEYINPUT55), .Z(n639) );
  XNOR2_X1 U707 ( .A(n637), .B(n639), .ZN(n640) );
  XNOR2_X1 U708 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X2 U709 ( .A1(n642), .A2(n717), .ZN(n644) );
  XNOR2_X1 U710 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n644), .B(n643), .ZN(G51) );
  NAND2_X1 U712 ( .A1(n711), .A2(G475), .ZN(n646) );
  XNOR2_X1 U713 ( .A(KEYINPUT118), .B(KEYINPUT60), .ZN(n647) );
  XNOR2_X1 U714 ( .A(n347), .B(n647), .ZN(G60) );
  NAND2_X1 U715 ( .A1(n649), .A2(n661), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n648), .B(G104), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n651) );
  NAND2_X1 U718 ( .A1(n649), .A2(n664), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U720 ( .A(G107), .B(n652), .ZN(G9) );
  INV_X1 U721 ( .A(n664), .ZN(n653) );
  NOR2_X1 U722 ( .A1(n659), .A2(n653), .ZN(n655) );
  XNOR2_X1 U723 ( .A(KEYINPUT112), .B(KEYINPUT29), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U725 ( .A(G128), .B(n656), .ZN(G30) );
  XOR2_X1 U726 ( .A(G143), .B(n657), .Z(G45) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U728 ( .A(G146), .B(n660), .Z(G48) );
  XOR2_X1 U729 ( .A(G113), .B(KEYINPUT113), .Z(n663) );
  NAND2_X1 U730 ( .A1(n665), .A2(n661), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(G15) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n666), .B(G116), .ZN(G18) );
  XNOR2_X1 U734 ( .A(G125), .B(n667), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U736 ( .A(G134), .B(n669), .ZN(G36) );
  INV_X1 U737 ( .A(n670), .ZN(n671) );
  XNOR2_X1 U738 ( .A(n671), .B(KEYINPUT83), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n708) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n686) );
  NOR2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U742 ( .A(n676), .B(KEYINPUT50), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n679), .A2(n537), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n680), .B(KEYINPUT49), .ZN(n681) );
  NAND2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U748 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U749 ( .A(n687), .B(KEYINPUT114), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n704), .A2(n688), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n350), .A2(n689), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U755 ( .A1(n703), .A2(n696), .ZN(n697) );
  NOR2_X1 U756 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n699), .B(KEYINPUT52), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n702), .B(KEYINPUT116), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U761 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U763 ( .A1(n709), .A2(G953), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n710), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U765 ( .A1(n346), .A2(G217), .ZN(n715) );
  XOR2_X1 U766 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n712) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U768 ( .A1(G953), .A2(G224), .ZN(n718) );
  XOR2_X1 U769 ( .A(KEYINPUT61), .B(n718), .Z(n719) );
  NOR2_X1 U770 ( .A1(n720), .A2(n719), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n721), .B(KEYINPUT123), .ZN(n722) );
  NOR2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U773 ( .A(KEYINPUT124), .B(n724), .Z(n731) );
  XNOR2_X1 U774 ( .A(G101), .B(n725), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U777 ( .A(n731), .B(n730), .Z(G69) );
  XNOR2_X1 U778 ( .A(n733), .B(n732), .ZN(n736) );
  XNOR2_X1 U779 ( .A(n734), .B(n736), .ZN(n735) );
  NAND2_X1 U780 ( .A1(n735), .A2(n456), .ZN(n741) );
  XNOR2_X1 U781 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U782 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U783 ( .A1(n738), .A2(G953), .ZN(n739) );
  XOR2_X1 U784 ( .A(KEYINPUT125), .B(n739), .Z(n740) );
  NAND2_X1 U785 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U786 ( .A(G122), .B(KEYINPUT126), .ZN(n742) );
  XOR2_X1 U787 ( .A(G140), .B(n743), .Z(G42) );
  XOR2_X1 U788 ( .A(G119), .B(n744), .Z(G21) );
  XOR2_X1 U789 ( .A(G137), .B(n745), .Z(G39) );
  XOR2_X1 U790 ( .A(n746), .B(G131), .Z(G33) );
  XOR2_X1 U791 ( .A(G101), .B(n747), .Z(G3) );
endmodule

