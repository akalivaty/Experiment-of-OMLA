//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G107), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT80), .A3(G104), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n192), .A2(KEYINPUT80), .A3(KEYINPUT3), .A4(G104), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n191), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n190), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G101), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(KEYINPUT81), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G101), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(new_n190), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n195), .B2(new_n196), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT4), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n199), .B1(new_n202), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G116), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT69), .B1(new_n211), .B2(G119), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n213));
  INV_X1    g027(.A(G119), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G116), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G119), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT68), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n219));
  INV_X1    g033(.A(G113), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT67), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(KEYINPUT2), .B2(G113), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n221), .A2(new_n223), .B1(KEYINPUT2), .B2(G113), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT2), .A2(G113), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n222), .A2(KEYINPUT2), .A3(G113), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n219), .B2(new_n220), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n188), .B1(new_n210), .B2(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n203), .A2(new_n205), .A3(new_n190), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n200), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n234), .B(KEYINPUT4), .C1(new_n198), .C2(new_n197), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n201), .A2(new_n208), .A3(G101), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n235), .A2(new_n231), .A3(new_n188), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n192), .A2(G104), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n198), .B1(new_n238), .B2(new_n190), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n200), .B2(new_n233), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT83), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT83), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n207), .B2(new_n239), .ZN(new_n243));
  XOR2_X1   g057(.A(KEYINPUT87), .B(KEYINPUT5), .Z(new_n244));
  NOR2_X1   g058(.A1(new_n211), .A2(G119), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n220), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT87), .B(KEYINPUT5), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(new_n212), .A3(new_n215), .A4(new_n216), .ZN(new_n248));
  INV_X1    g062(.A(new_n217), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n246), .A2(new_n248), .B1(new_n249), .B2(new_n224), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n241), .A2(new_n243), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n237), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n187), .B1(new_n232), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n235), .A2(new_n231), .A3(new_n236), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT86), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n255), .A2(KEYINPUT88), .A3(new_n251), .A4(new_n237), .ZN(new_n256));
  XNOR2_X1  g070(.A(G110), .B(G122), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n255), .A2(new_n251), .A3(new_n237), .A4(new_n257), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n260), .A2(KEYINPUT6), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n253), .A2(new_n263), .A3(new_n256), .A4(new_n258), .ZN(new_n264));
  INV_X1    g078(.A(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n267), .A2(G146), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT65), .B1(new_n265), .B2(G143), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n267), .A3(G146), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n270), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G125), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n266), .A2(new_n268), .A3(new_n281), .A4(G128), .ZN(new_n282));
  INV_X1    g096(.A(G128), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n266), .B2(KEYINPUT1), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n275), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n280), .B1(G125), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G224), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G953), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n286), .B(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n262), .A2(new_n264), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n240), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n250), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n257), .B(KEYINPUT8), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n294), .A2(new_n246), .B1(new_n224), .B2(new_n249), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n292), .B(new_n293), .C1(new_n295), .C2(new_n291), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n286), .B1(new_n297), .B2(new_n288), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n286), .A2(new_n297), .A3(new_n288), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n301), .B2(new_n260), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n290), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n290), .B2(new_n302), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT89), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT89), .B(new_n303), .C1(new_n290), .C2(new_n302), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  OAI21_X1  g126(.A(G221), .B1(new_n312), .B2(G902), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n313), .B(KEYINPUT79), .Z(new_n314));
  NAND4_X1  g128(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT10), .A4(new_n285), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n316));
  INV_X1    g130(.A(new_n282), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT1), .B1(new_n267), .B2(G146), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT82), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n266), .A2(new_n320), .A3(KEYINPUT1), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(G128), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n266), .A2(new_n268), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n316), .B1(new_n291), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n273), .B1(new_n267), .B2(G146), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n265), .A2(KEYINPUT65), .A3(G143), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n266), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n326), .B1(new_n329), .B2(new_n277), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n235), .A2(new_n330), .A3(new_n236), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n315), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT11), .ZN(new_n335));
  INV_X1    g149(.A(G134), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(G137), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(G137), .ZN(new_n338));
  INV_X1    g152(.A(G137), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT11), .A3(G134), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G131), .ZN(new_n342));
  INV_X1    g156(.A(G131), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n337), .A2(new_n340), .A3(new_n343), .A4(new_n338), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n315), .A2(new_n331), .A3(KEYINPUT84), .A4(new_n325), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n334), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n345), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n315), .A2(new_n331), .A3(new_n348), .A4(new_n325), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G140), .ZN(new_n350));
  INV_X1    g164(.A(G953), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(G227), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n350), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n291), .A2(new_n324), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n240), .A2(new_n285), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n345), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT12), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n281), .B1(G143), .B2(new_n265), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n283), .B1(new_n362), .B2(new_n320), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n363), .A2(new_n319), .B1(new_n266), .B2(new_n268), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n240), .B1(new_n364), .B2(new_n317), .ZN(new_n365));
  INV_X1    g179(.A(new_n284), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n329), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n367), .B(new_n282), .C1(new_n207), .C2(new_n239), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT12), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n345), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n361), .A2(new_n349), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n353), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n357), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G469), .B1(new_n375), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n361), .A2(new_n371), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n377), .B1(new_n378), .B2(new_n355), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n370), .B1(new_n369), .B2(new_n345), .ZN(new_n380));
  AOI211_X1 g194(.A(KEYINPUT12), .B(new_n348), .C1(new_n365), .C2(new_n368), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n382), .A2(KEYINPUT85), .A3(new_n349), .A4(new_n354), .ZN(new_n383));
  INV_X1    g197(.A(new_n349), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n348), .B1(new_n332), .B2(new_n333), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(new_n346), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n379), .B(new_n383), .C1(new_n386), .C2(new_n354), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT73), .B(G902), .Z(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n314), .B1(new_n376), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G952), .ZN(new_n392));
  AOI211_X1 g206(.A(G953), .B(new_n392), .C1(G234), .C2(G237), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n351), .B(new_n389), .C1(G234), .C2(G237), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n267), .A2(G128), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n283), .A2(G143), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n336), .ZN(new_n401));
  XNOR2_X1  g215(.A(G116), .B(G122), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n192), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n211), .A2(KEYINPUT14), .A3(G122), .ZN(new_n404));
  INV_X1    g218(.A(new_n402), .ZN(new_n405));
  OAI211_X1 g219(.A(G107), .B(new_n404), .C1(new_n405), .C2(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n398), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n399), .B1(new_n408), .B2(KEYINPUT13), .ZN(new_n410));
  OAI21_X1  g224(.A(G134), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n400), .A2(new_n336), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n402), .B(new_n192), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G217), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n312), .A2(new_n415), .A3(G953), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n416), .B1(new_n407), .B2(new_n414), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n389), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT93), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(new_n389), .C1(new_n418), .C2(new_n419), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n420), .A2(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G902), .ZN(new_n429));
  INV_X1    g243(.A(G237), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n351), .A3(G214), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n267), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n430), .A2(new_n351), .A3(G143), .A4(G214), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n343), .A3(new_n433), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(KEYINPUT75), .A2(G125), .ZN(new_n439));
  INV_X1    g253(.A(G140), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(KEYINPUT16), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT16), .ZN(new_n444));
  INV_X1    g258(.A(G125), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(G140), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n265), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n265), .B1(new_n443), .B2(new_n446), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n434), .A2(KEYINPUT17), .A3(G131), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n438), .A2(new_n447), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n441), .A2(G146), .A3(new_n442), .ZN(new_n452));
  XNOR2_X1  g266(.A(G125), .B(G140), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT76), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n453), .A2(new_n454), .A3(new_n265), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(new_n453), .B2(new_n265), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT18), .A2(G131), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n434), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n432), .A2(new_n433), .A3(new_n458), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n457), .B(new_n460), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G113), .B(G122), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(new_n189), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n451), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n451), .B2(new_n464), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n429), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G475), .ZN(new_n470));
  NOR2_X1   g284(.A1(G475), .A2(G902), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT19), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n453), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n441), .A2(KEYINPUT19), .A3(new_n442), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n265), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT91), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n473), .A2(new_n474), .A3(new_n477), .A4(new_n265), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n448), .B1(new_n435), .B2(new_n437), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n466), .B1(new_n481), .B2(new_n464), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n471), .B1(new_n467), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT20), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n451), .A2(new_n464), .A3(new_n466), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n457), .A2(new_n460), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n461), .B(KEYINPUT90), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n487), .A2(new_n488), .B1(new_n479), .B2(new_n480), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n486), .B1(new_n489), .B2(new_n466), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n485), .B1(new_n490), .B2(new_n471), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n470), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(KEYINPUT92), .B(new_n470), .C1(new_n484), .C2(new_n491), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n428), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n391), .A2(new_n397), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n311), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n453), .A2(new_n265), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT76), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n453), .A2(new_n454), .A3(new_n265), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n214), .B2(G128), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n283), .A2(KEYINPUT23), .A3(G119), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n505), .C1(G119), .C2(new_n283), .ZN(new_n506));
  XNOR2_X1  g320(.A(G119), .B(G128), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  OAI22_X1  g322(.A1(new_n506), .A2(G110), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n502), .A2(new_n449), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n506), .A2(G110), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  INV_X1    g325(.A(new_n447), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n448), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n351), .A2(G221), .A3(G234), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT77), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT22), .B(G137), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n510), .A3(new_n513), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n415), .B1(new_n389), .B2(G234), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(G902), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT78), .ZN(new_n525));
  INV_X1    g339(.A(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(new_n389), .A3(new_n521), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n520), .A2(KEYINPUT25), .A3(new_n389), .A4(new_n521), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G472), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n279), .B1(new_n344), .B2(new_n342), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n339), .A2(G134), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n336), .A2(G137), .ZN(new_n537));
  OAI21_X1  g351(.A(G131), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n344), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n367), .B2(new_n282), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n535), .A2(new_n540), .A3(new_n231), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n330), .A2(new_n345), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n344), .A2(new_n538), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n285), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n542), .A2(new_n544), .B1(new_n225), .B2(new_n230), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT28), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT26), .B(G101), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n430), .A2(new_n351), .A3(G210), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n550), .B(KEYINPUT71), .Z(new_n551));
  XNOR2_X1  g365(.A(new_n549), .B(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n345), .A2(new_n330), .B1(new_n543), .B2(new_n285), .ZN(new_n553));
  INV_X1    g367(.A(new_n231), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT28), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n546), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT29), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n389), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n553), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n542), .A2(new_n544), .ZN(new_n563));
  INV_X1    g377(.A(new_n561), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT66), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n554), .B1(new_n553), .B2(KEYINPUT30), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n541), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n558), .B(new_n557), .C1(new_n568), .C2(new_n552), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT72), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n559), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n552), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT30), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n231), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n562), .B2(new_n565), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n572), .B1(new_n575), .B2(new_n541), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n576), .A2(KEYINPUT72), .A3(new_n558), .A4(new_n557), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n534), .B1(new_n571), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n568), .A2(KEYINPUT31), .A3(new_n552), .ZN(new_n579));
  NOR2_X1   g393(.A1(G472), .A2(G902), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n563), .A2(new_n231), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n553), .A2(new_n554), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n555), .B1(new_n584), .B2(KEYINPUT28), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n581), .B1(new_n585), .B2(new_n552), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n575), .A2(new_n541), .A3(new_n572), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n579), .B(new_n580), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT32), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n546), .A2(new_n556), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT31), .B1(new_n590), .B2(new_n572), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n568), .A2(new_n552), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT32), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n579), .A4(new_n580), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n578), .A2(KEYINPUT74), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n557), .A2(new_n558), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT66), .B1(new_n563), .B2(new_n564), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n560), .B(new_n561), .C1(new_n542), .C2(new_n544), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n567), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n552), .B1(new_n600), .B2(new_n583), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n570), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n559), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n577), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT74), .B1(new_n604), .B2(G472), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n533), .B1(new_n596), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n498), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n203), .A2(new_n205), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n609), .B(new_n610), .Z(G3));
  NAND2_X1  g425(.A1(new_n290), .A2(new_n302), .ZN(new_n612));
  INV_X1    g426(.A(new_n303), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n290), .A2(new_n302), .A3(new_n303), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n309), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n494), .A2(new_n495), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  INV_X1    g433(.A(new_n419), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n417), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n418), .A2(KEYINPUT33), .A3(new_n419), .ZN(new_n622));
  OAI211_X1 g436(.A(G478), .B(new_n389), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n616), .A2(new_n397), .A3(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n579), .B(new_n389), .C1(new_n586), .C2(new_n587), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G472), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n588), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n391), .A2(new_n631), .A3(new_n532), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G104), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n614), .A2(new_n615), .ZN(new_n637));
  INV_X1    g451(.A(new_n428), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n492), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n637), .A2(new_n308), .A3(new_n397), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n632), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT95), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n531), .ZN(new_n645));
  INV_X1    g459(.A(new_n523), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(new_n514), .Z(new_n648));
  OAI21_X1  g462(.A(new_n645), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n629), .A2(new_n588), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n498), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT37), .B(G110), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  NAND3_X1  g467(.A1(new_n604), .A2(KEYINPUT74), .A3(G472), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n589), .A2(new_n595), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n616), .B1(new_n605), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n391), .ZN(new_n658));
  INV_X1    g472(.A(new_n649), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n639), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n393), .B1(new_n394), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  NAND4_X1  g480(.A1(new_n494), .A2(new_n308), .A3(new_n495), .A4(new_n428), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n649), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT96), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n663), .B(KEYINPUT39), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n391), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n568), .A2(new_n572), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n429), .B1(new_n584), .B2(new_n552), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n655), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n669), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n614), .A2(KEYINPUT89), .A3(new_n615), .ZN(new_n678));
  INV_X1    g492(.A(new_n310), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n677), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n267), .ZN(G45));
  INV_X1    g498(.A(new_n663), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n494), .A2(new_n495), .A3(new_n624), .A4(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n660), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  INV_X1    g503(.A(KEYINPUT97), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n387), .A2(new_n389), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n387), .B2(new_n389), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n314), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n694), .B(new_n532), .C1(new_n656), .C2(new_n605), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n627), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT41), .B(G113), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  OAI211_X1 g512(.A(new_n308), .B(new_n397), .C1(new_n304), .C2(new_n305), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n661), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT98), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n607), .A2(new_n700), .A3(new_n701), .A4(new_n694), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT98), .B1(new_n695), .B2(new_n640), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  OAI21_X1  g519(.A(new_n308), .B1(new_n304), .B2(new_n305), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n596), .B2(new_n606), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n496), .A2(new_n397), .A3(new_n649), .ZN(new_n708));
  INV_X1    g522(.A(new_n693), .ZN(new_n709));
  INV_X1    g523(.A(new_n314), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n387), .A2(new_n389), .A3(new_n691), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  AOI21_X1  g529(.A(new_n667), .B1(new_n614), .B2(new_n615), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT99), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT78), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n524), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n645), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT99), .B1(new_n525), .B2(new_n531), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n629), .A3(new_n588), .A4(new_n397), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n716), .A2(new_n694), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR2_X1   g540(.A1(new_n650), .A2(new_n686), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n616), .A2(new_n727), .A3(new_n694), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT100), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n706), .A2(new_n712), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT100), .A3(new_n727), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n347), .A2(new_n356), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(new_n347), .B2(new_n356), .ZN(new_n737));
  OAI211_X1 g551(.A(G469), .B(new_n373), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(G469), .A2(G902), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT101), .Z(new_n740));
  NAND3_X1  g554(.A1(new_n390), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(new_n710), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n742), .B(new_n308), .C1(new_n307), .C2(new_n310), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n687), .B(new_n722), .C1(new_n656), .C2(new_n605), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT42), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n309), .B1(new_n678), .B2(new_n679), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n607), .A2(new_n746), .A3(new_n742), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT103), .B(G131), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G33));
  NAND4_X1  g565(.A1(new_n607), .A2(new_n746), .A3(new_n664), .A4(new_n742), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  INV_X1    g567(.A(new_n740), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT45), .B(new_n373), .C1(new_n736), .C2(new_n737), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n388), .B1(new_n374), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT104), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n755), .A2(new_n757), .A3(KEYINPUT104), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n754), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT46), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n390), .B1(new_n762), .B2(KEYINPUT46), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n710), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n617), .A2(new_n624), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT105), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT43), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n625), .B1(new_n494), .B2(new_n495), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(KEYINPUT105), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n770), .A2(new_n773), .A3(new_n630), .A4(new_n649), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n746), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n670), .A2(new_n767), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n339), .ZN(G39));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n766), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT47), .B(new_n710), .C1(new_n764), .C2(new_n765), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n596), .A2(new_n606), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n777), .A2(new_n785), .A3(new_n532), .A4(new_n686), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  NOR2_X1   g603(.A1(G952), .A2(G953), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n655), .A2(new_n532), .A3(new_n393), .A4(new_n675), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n624), .B1(new_n494), .B2(new_n495), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n308), .B(new_n694), .C1(new_n307), .C2(new_n310), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT108), .B1(new_n746), .B2(new_n694), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n793), .B(new_n794), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n796), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n746), .A2(KEYINPUT108), .A3(new_n694), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n792), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n801), .B1(new_n804), .B2(new_n794), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n770), .A2(new_n773), .A3(new_n393), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n797), .B2(new_n798), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n802), .A2(new_n803), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(KEYINPUT109), .A3(new_n808), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n650), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n791), .B1(new_n806), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n650), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT109), .B1(new_n812), .B2(new_n808), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n810), .B(new_n807), .C1(new_n802), .C2(new_n803), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n804), .A2(new_n801), .A3(new_n794), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n822), .A3(KEYINPUT112), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n631), .A2(new_n722), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n694), .A2(new_n309), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n807), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n681), .A2(new_n826), .A3(KEYINPUT50), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT50), .B1(new_n681), .B2(new_n826), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT51), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n692), .A2(new_n693), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT106), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n314), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n782), .A2(new_n783), .A3(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n777), .A2(new_n807), .A3(new_n824), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n829), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n815), .A2(new_n823), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n804), .A2(new_n626), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n807), .A2(new_n824), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n392), .B(G953), .C1(new_n838), .C2(new_n731), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n722), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n596), .B2(new_n606), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n817), .B2(new_n818), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT48), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT48), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n845), .B(new_n842), .C1(new_n817), .C2(new_n818), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n840), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n836), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n658), .A2(new_n659), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n707), .B(new_n850), .C1(new_n664), .C2(new_n687), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n649), .A2(new_n663), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT107), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n716), .A3(new_n742), .A4(new_n676), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n733), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n733), .A2(new_n851), .A3(KEYINPUT52), .A4(new_n854), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n695), .A2(new_n627), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n311), .B(new_n497), .C1(new_n607), .C2(new_n816), .ZN(new_n861));
  INV_X1    g675(.A(new_n632), .ZN(new_n862));
  INV_X1    g676(.A(new_n496), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n494), .A2(new_n625), .A3(new_n495), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n311), .A2(new_n862), .A3(new_n397), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n712), .A2(new_n723), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n707), .A2(new_n713), .B1(new_n716), .B2(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n860), .A2(new_n861), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n745), .A2(new_n748), .A3(new_n752), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n492), .A2(new_n428), .A3(new_n663), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n850), .A2(new_n785), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n742), .A2(new_n727), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n777), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n869), .A2(new_n704), .A3(new_n870), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n849), .B1(new_n859), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n694), .A2(new_n397), .A3(new_n496), .A4(new_n649), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n725), .B1(new_n657), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n696), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n704), .A3(new_n866), .A4(new_n861), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n745), .A2(new_n748), .A3(new_n752), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n874), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n857), .A2(new_n858), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(KEYINPUT53), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT54), .B1(new_n877), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n877), .A2(KEYINPUT54), .A3(new_n885), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n848), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n819), .B(new_n822), .C1(new_n828), .C2(new_n827), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(KEYINPUT111), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n890), .A2(KEYINPUT111), .B1(new_n833), .B2(new_n834), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT51), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n790), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT49), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n831), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n831), .A2(new_n896), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n722), .A2(new_n308), .A3(new_n710), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n676), .A2(new_n899), .A3(new_n768), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n897), .A2(new_n681), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n789), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n888), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n836), .B(new_n847), .C1(new_n904), .C2(new_n886), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n893), .ZN(new_n906));
  OAI211_X1 g720(.A(KEYINPUT113), .B(new_n901), .C1(new_n906), .C2(new_n790), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n907), .ZN(G75));
  NAND2_X1  g722(.A1(new_n392), .A2(G953), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT115), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n877), .A2(new_n885), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n912), .A2(new_n389), .A3(new_n303), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n262), .A2(new_n264), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n289), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT55), .Z(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT56), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n910), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT114), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n913), .A2(new_n919), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n918), .B1(new_n923), .B2(new_n916), .ZN(G51));
  INV_X1    g738(.A(new_n910), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n904), .A2(new_n886), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n740), .B(KEYINPUT57), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(KEYINPUT116), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n887), .A2(new_n888), .A3(new_n927), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT116), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n928), .A2(new_n931), .A3(new_n387), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n912), .A2(new_n389), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n760), .A3(new_n761), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n925), .B1(new_n932), .B2(new_n934), .ZN(G54));
  NAND2_X1  g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT117), .Z(new_n937));
  AND3_X1   g751(.A1(new_n933), .A2(new_n490), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n490), .B1(new_n933), .B2(new_n937), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n939), .A3(new_n925), .ZN(G60));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT59), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n621), .A2(new_n622), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT118), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n926), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n926), .B2(new_n942), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n925), .ZN(G63));
  INV_X1    g761(.A(new_n648), .ZN(new_n948));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT119), .B1(new_n911), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n953), .B(new_n950), .C1(new_n877), .C2(new_n885), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n948), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n861), .A2(new_n866), .A3(new_n868), .A4(new_n860), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n702), .A2(new_n703), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n874), .ZN(new_n958));
  AND4_X1   g772(.A1(KEYINPUT53), .A2(new_n884), .A3(new_n958), .A4(new_n870), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT53), .B1(new_n883), .B2(new_n884), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n951), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n953), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n911), .A2(KEYINPUT119), .A3(new_n951), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n520), .A2(new_n521), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT120), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n955), .A2(new_n966), .A3(new_n910), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n648), .B1(new_n962), .B2(new_n963), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(KEYINPUT121), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT61), .B1(new_n955), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n955), .A2(new_n966), .A3(new_n910), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n971), .A2(new_n975), .ZN(G66));
  XNOR2_X1  g790(.A(new_n881), .B(KEYINPUT122), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n351), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n395), .B2(new_n287), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT123), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n914), .B1(G898), .B2(new_n351), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT124), .Z(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT125), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n981), .B(new_n984), .ZN(G69));
  AOI21_X1  g799(.A(new_n351), .B1(G227), .B2(G900), .ZN(new_n986));
  INV_X1    g800(.A(new_n865), .ZN(new_n987));
  NOR4_X1   g801(.A1(new_n608), .A2(new_n777), .A3(new_n987), .A4(new_n671), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n733), .A2(new_n851), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n683), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n779), .B1(new_n784), .B2(new_n786), .ZN(new_n994));
  AOI21_X1  g808(.A(G953), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n566), .A2(new_n573), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n473), .A2(new_n474), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT126), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(G900), .A2(G953), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n767), .A2(new_n670), .A3(new_n716), .A4(new_n842), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n882), .A2(new_n989), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n994), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n998), .B(new_n1000), .C1(new_n1003), .C2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n995), .A2(KEYINPUT126), .A3(new_n998), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n986), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1006), .ZN(new_n1008));
  INV_X1    g822(.A(new_n986), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1008), .A2(new_n999), .A3(new_n1009), .A4(new_n1004), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n1003), .B2(new_n977), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n568), .A2(new_n572), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n673), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n911), .A2(new_n1018), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n993), .A2(new_n994), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1013), .B1(new_n1021), .B2(new_n977), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n925), .B(new_n1020), .C1(new_n673), .C2(new_n1022), .ZN(G57));
endmodule


