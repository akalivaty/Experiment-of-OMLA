//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT89), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n203), .A2(new_n204), .B1(new_n205), .B2(new_n202), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n202), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n206), .A2(KEYINPUT90), .A3(G8gat), .A4(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT91), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(KEYINPUT91), .A3(new_n212), .ZN(new_n216));
  NOR2_X1   g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  XOR2_X1   g016(.A(new_n217), .B(KEYINPUT14), .Z(new_n218));
  XNOR2_X1  g017(.A(G43gat), .B(G50gat), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT88), .B(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G29gat), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n218), .A2(new_n220), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n222), .A2(G29gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n217), .B(KEYINPUT14), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT15), .B(new_n219), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n215), .A2(new_n216), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT17), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n213), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n229), .A2(KEYINPUT18), .A3(new_n230), .A4(new_n234), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n224), .A2(new_n227), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n211), .A2(KEYINPUT91), .A3(new_n212), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT91), .B1(new_n211), .B2(new_n212), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n229), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n230), .B(KEYINPUT13), .Z(new_n244));
  AOI21_X1  g043(.A(KEYINPUT92), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT92), .ZN(new_n246));
  INV_X1    g045(.A(new_n244), .ZN(new_n247));
  AOI211_X1 g046(.A(new_n246), .B(new_n247), .C1(new_n242), .C2(new_n229), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n237), .B(new_n238), .C1(new_n245), .C2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT11), .ZN(new_n251));
  INV_X1    g050(.A(G169gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G197gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(KEYINPUT12), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n244), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n246), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n243), .A2(KEYINPUT92), .A3(new_n244), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n237), .A2(new_n238), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n256), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT32), .ZN(new_n267));
  XNOR2_X1  g066(.A(G15gat), .B(G43gat), .ZN(new_n268));
  INV_X1    g067(.A(G71gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT74), .ZN(new_n271));
  INV_X1    g070(.A(G99gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n267), .B1(new_n273), .B2(KEYINPUT33), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G190gat), .ZN(new_n278));
  INV_X1    g077(.A(G183gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT27), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT27), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G183gat), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n276), .A2(new_n278), .A3(new_n280), .A4(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G176gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n252), .A2(new_n286), .A3(KEYINPUT26), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT26), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  AND2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n287), .B(new_n288), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  AND4_X1   g091(.A1(new_n276), .A2(new_n278), .A3(new_n280), .A4(new_n282), .ZN(new_n293));
  NOR2_X1   g092(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n252), .A2(new_n286), .ZN(new_n296));
  AND2_X1   g095(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n297));
  NOR2_X1   g096(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n296), .B(KEYINPUT66), .C1(new_n297), .C2(new_n298), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n252), .A2(new_n286), .A3(KEYINPUT23), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NOR3_X1   g108(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n288), .A2(KEYINPUT24), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n307), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n285), .A2(new_n295), .B1(new_n303), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n304), .A2(new_n306), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT25), .ZN(new_n322));
  NAND2_X1  g121(.A1(G113gat), .A2(G120gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(G113gat), .A2(G120gat), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT70), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G113gat), .ZN(new_n327));
  INV_X1    g126(.A(G120gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n323), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT71), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT1), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G127gat), .B(G134gat), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n326), .A2(new_n331), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G134gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(G127gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT69), .B(G134gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(G127gat), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT1), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n322), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT72), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n317), .A2(new_n322), .A3(new_n345), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n317), .A2(new_n322), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n344), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n353));
  NAND2_X1  g152(.A1(G227gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n352), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n274), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n267), .A2(KEYINPUT33), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n352), .A2(new_n355), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT73), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n273), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n358), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n347), .A2(new_n351), .A3(new_n354), .A4(new_n349), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n367), .B(KEYINPUT34), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n358), .B(new_n368), .C1(new_n364), .C2(new_n365), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT36), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(KEYINPUT36), .A3(new_n371), .ZN(new_n375));
  INV_X1    g174(.A(G141gat), .ZN(new_n376));
  INV_X1    g175(.A(G148gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT2), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT2), .ZN(new_n382));
  NAND2_X1  g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n378), .A2(new_n380), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G162gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G155gat), .ZN(new_n386));
  INV_X1    g185(.A(G155gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G162gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(KEYINPUT78), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G155gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n379), .B1(new_n394), .B2(G162gat), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n378), .A2(new_n386), .A3(new_n388), .A4(new_n383), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n344), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n339), .A2(KEYINPUT69), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT69), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(G134gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n401), .A3(G127gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(G127gat), .B2(new_n339), .ZN(new_n403));
  INV_X1    g202(.A(new_n343), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT78), .B(G155gat), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT2), .B1(new_n406), .B2(new_n385), .ZN(new_n407));
  INV_X1    g206(.A(new_n396), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n405), .A2(new_n409), .A3(new_n338), .A4(new_n390), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n344), .A2(KEYINPUT80), .A3(new_n397), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT4), .B1(new_n344), .B2(new_n397), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n407), .A2(new_n408), .B1(new_n389), .B2(new_n384), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n405), .A4(new_n338), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n422), .A3(KEYINPUT79), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n392), .A2(G155gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n387), .A2(KEYINPUT78), .ZN(new_n425));
  OAI21_X1  g224(.A(G162gat), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n396), .B1(new_n426), .B2(KEYINPUT2), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n384), .A2(new_n389), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT3), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n390), .B(new_n430), .C1(new_n395), .C2(new_n396), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n344), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n410), .A2(new_n433), .A3(KEYINPUT4), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n423), .A2(new_n413), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n412), .A2(KEYINPUT81), .A3(new_n414), .A4(new_n415), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n418), .A2(new_n435), .A3(KEYINPUT5), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n432), .A3(new_n439), .A4(new_n413), .ZN(new_n440));
  XOR2_X1   g239(.A(KEYINPUT82), .B(KEYINPUT0), .Z(new_n441));
  XNOR2_X1  g240(.A(G1gat), .B(G29gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G57gat), .B(G85gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n437), .A2(new_n440), .ZN(new_n449));
  INV_X1    g248(.A(new_n445), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(G211gat), .A2(G218gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(G211gat), .A2(G218gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(G197gat), .A2(G204gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(G197gat), .A2(G204gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G211gat), .B(G218gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(G197gat), .B(G204gat), .ZN(new_n464));
  INV_X1    g263(.A(new_n461), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT75), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n303), .A2(new_n316), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT67), .B(G190gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT27), .B(G183gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n294), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n296), .A2(new_n289), .A3(new_n306), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n287), .A2(new_n288), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n285), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n305), .B1(new_n303), .B2(new_n320), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n469), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT29), .B1(new_n317), .B2(new_n322), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n467), .B(new_n479), .C1(new_n480), .C2(new_n468), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n477), .B2(new_n478), .ZN(new_n483));
  INV_X1    g282(.A(new_n469), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n483), .A2(new_n484), .B1(new_n350), .B2(new_n468), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n481), .B1(new_n485), .B2(new_n467), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT76), .ZN(new_n488));
  XNOR2_X1  g287(.A(G8gat), .B(G36gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(G64gat), .ZN(new_n490));
  INV_X1    g289(.A(G92gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT30), .A4(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n481), .B(new_n492), .C1(new_n485), .C2(new_n467), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT76), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  INV_X1    g296(.A(new_n492), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n486), .A2(new_n498), .ZN(new_n499));
  AND4_X1   g298(.A1(new_n493), .A2(new_n496), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n437), .A2(KEYINPUT83), .A3(new_n440), .A4(new_n445), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n453), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n451), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n454), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G50gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G228gat), .ZN(new_n507));
  INV_X1    g306(.A(G233gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n467), .A2(new_n482), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT84), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT3), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT29), .B1(new_n462), .B2(new_n466), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT84), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n420), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n467), .B1(new_n431), .B2(new_n482), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n397), .A2(new_n514), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n429), .A3(new_n509), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT85), .B1(new_n520), .B2(new_n517), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n431), .A2(new_n482), .ZN(new_n522));
  INV_X1    g321(.A(new_n467), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT85), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n510), .B1(new_n397), .B2(KEYINPUT3), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n519), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G22gat), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n518), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n518), .B2(new_n528), .ZN(new_n531));
  XNOR2_X1  g330(.A(G78gat), .B(G106gat), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n532), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n521), .A2(new_n527), .ZN(new_n535));
  INV_X1    g334(.A(new_n515), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n430), .B1(new_n514), .B2(KEYINPUT84), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n397), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n509), .B1(new_n538), .B2(new_n524), .ZN(new_n539));
  OAI21_X1  g338(.A(G22gat), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n528), .A3(new_n529), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n534), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n506), .B1(new_n533), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n532), .B1(new_n530), .B2(new_n531), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n541), .A3(new_n534), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n505), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n374), .A2(new_n375), .B1(new_n504), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n500), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n413), .B1(new_n438), .B2(new_n432), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT39), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n412), .A2(new_n415), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(new_n414), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n450), .B1(new_n551), .B2(new_n552), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  NAND3_X1  g358(.A1(new_n550), .A2(new_n559), .A3(new_n451), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n486), .A2(KEYINPUT37), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n498), .B1(new_n486), .B2(KEYINPUT37), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT38), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n523), .B(new_n479), .C1(new_n480), .C2(new_n468), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(KEYINPUT37), .C1(new_n485), .C2(new_n523), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT38), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n563), .B(new_n494), .C1(new_n562), .C2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n503), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT6), .B1(new_n448), .B2(new_n451), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n560), .B(new_n547), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n547), .A2(new_n370), .A3(new_n371), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT35), .B1(new_n574), .B2(new_n504), .ZN(new_n575));
  INV_X1    g374(.A(new_n371), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n359), .B1(new_n356), .B2(new_n357), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n273), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n368), .B1(new_n578), .B2(new_n358), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n454), .A2(new_n500), .A3(KEYINPUT87), .A4(new_n503), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT35), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n547), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT87), .B1(new_n571), .B2(new_n500), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n575), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n266), .B1(new_n573), .B2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G57gat), .B(G64gat), .Z(new_n587));
  OR2_X1    g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n589), .B(new_n588), .C1(new_n594), .C2(new_n591), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n597));
  INV_X1    g396(.A(G231gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n508), .ZN(new_n599));
  OAI211_X1 g398(.A(G231gat), .B(G233gat), .C1(new_n596), .C2(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n605), .A3(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n240), .B2(new_n241), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G183gat), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n279), .B(new_n608), .C1(new_n240), .C2(new_n241), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G211gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n610), .A2(new_n607), .A3(new_n611), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n615), .ZN(new_n618));
  INV_X1    g417(.A(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(new_n612), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT7), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(G85gat), .A3(G92gat), .A4(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(G85gat), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n628), .B(new_n629), .C1(new_n633), .C2(new_n491), .ZN(new_n634));
  NAND2_X1  g433(.A1(G99gat), .A2(G106gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(KEYINPUT8), .A2(new_n635), .B1(new_n633), .B2(new_n491), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G99gat), .B(G106gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n632), .A2(new_n638), .A3(new_n634), .A4(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n627), .B1(new_n239), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT96), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n645), .B(new_n627), .C1(new_n239), .C2(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n233), .A2(new_n648), .A3(new_n231), .A4(new_n642), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n233), .A2(new_n231), .A3(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT95), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G134gat), .B(G162gat), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n644), .A2(new_n646), .B1(KEYINPUT95), .B2(new_n650), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(new_n649), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n626), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n655), .A3(new_n649), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n625), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n639), .A2(KEYINPUT97), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n596), .A2(new_n641), .A3(new_n640), .A4(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n593), .A2(new_n663), .A3(new_n595), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n642), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n641), .A4(new_n640), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G176gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(G204gat), .Z(new_n675));
  AND2_X1   g474(.A1(new_n664), .A2(new_n666), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n672), .B(new_n675), .C1(new_n676), .C2(new_n671), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  INV_X1    g477(.A(new_n671), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n668), .B2(new_n669), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n676), .A2(new_n671), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n621), .A2(new_n662), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n586), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n571), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT98), .B(G1gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1324gat));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n586), .A2(new_n550), .A3(new_n684), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT99), .Z(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n690), .A2(new_n689), .A3(new_n692), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n691), .B2(G8gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1325gat));
  NAND2_X1  g495(.A1(new_n374), .A2(new_n375), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n685), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n372), .A2(G15gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n685), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n547), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT100), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n701), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(new_n621), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n654), .A2(new_n657), .A3(new_n626), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n625), .B1(new_n659), .B2(new_n660), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n705), .A2(new_n708), .A3(new_n683), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n586), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(G29gat), .ZN(new_n711));
  INV_X1    g510(.A(new_n571), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n573), .A2(new_n585), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(KEYINPUT44), .A3(new_n662), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n266), .A2(new_n705), .A3(new_n683), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n706), .B2(new_n707), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n658), .A2(KEYINPUT102), .A3(new_n661), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n585), .A2(new_n722), .B1(new_n572), .B2(new_n549), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n575), .B(KEYINPUT101), .C1(new_n583), .C2(new_n584), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n716), .B(new_n717), .C1(new_n725), .C2(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n726), .B2(new_n571), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n714), .A2(new_n727), .ZN(G1328gat));
  NOR2_X1   g527(.A1(new_n500), .A2(new_n222), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n710), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n731));
  OR2_X1    g530(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n731), .B2(new_n730), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT104), .B1(new_n726), .B2(new_n500), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n222), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n726), .A2(KEYINPUT104), .A3(new_n500), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(G1329gat));
  OAI21_X1  g537(.A(G43gat), .B1(new_n726), .B2(new_n697), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n372), .A2(G43gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n710), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n739), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n739), .B2(new_n743), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1330gat));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n547), .A2(G50gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n710), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n748), .A2(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n585), .A2(new_n722), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n573), .A3(new_n724), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n719), .A2(new_n720), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n760), .A2(new_n548), .A3(new_n716), .A4(new_n717), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n750), .B(new_n754), .C1(G50gat), .C2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n750), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(G50gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n754), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n762), .A2(new_n766), .ZN(G1331gat));
  NAND4_X1  g566(.A1(new_n266), .A2(new_n705), .A3(new_n708), .A4(new_n683), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n723), .B2(new_n724), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n569), .B2(new_n570), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n454), .A2(KEYINPUT107), .A3(new_n503), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n550), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT49), .B(G64gat), .Z(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(G1333gat));
  INV_X1    g579(.A(new_n697), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n269), .B1(new_n769), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n372), .A2(G71gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n769), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n548), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n265), .A2(new_n705), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n662), .ZN(new_n790));
  AOI211_X1 g589(.A(new_n788), .B(new_n790), .C1(new_n723), .C2(new_n724), .ZN(new_n791));
  INV_X1    g590(.A(new_n790), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT51), .B1(new_n756), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n683), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n633), .A3(new_n712), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n789), .A2(new_n683), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n716), .B(new_n799), .C1(new_n725), .C2(KEYINPUT44), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800), .B2(new_n571), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(G1336gat));
  NAND3_X1  g601(.A1(new_n550), .A2(new_n491), .A3(new_n683), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT108), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n791), .B2(new_n793), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT109), .ZN(new_n806));
  OAI21_X1  g605(.A(G92gat), .B1(new_n800), .B2(new_n500), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n808), .B(new_n804), .C1(new_n791), .C2(new_n793), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT110), .B(new_n804), .C1(new_n791), .C2(new_n793), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n760), .A2(new_n550), .A3(new_n716), .A4(new_n799), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(new_n816), .B2(G92gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n811), .A2(new_n818), .ZN(G1337gat));
  NAND3_X1  g618(.A1(new_n796), .A2(new_n272), .A3(new_n580), .ZN(new_n820));
  OAI21_X1  g619(.A(G99gat), .B1(new_n800), .B2(new_n697), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1338gat));
  NOR2_X1   g621(.A1(new_n547), .A2(G106gat), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n683), .B(new_n823), .C1(new_n791), .C2(new_n793), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n800), .A2(new_n547), .ZN(new_n825));
  XNOR2_X1  g624(.A(KEYINPUT111), .B(G106gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1339gat));
  NAND3_X1  g630(.A1(new_n668), .A2(new_n669), .A3(new_n679), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n672), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n675), .B1(new_n680), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n677), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n835), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT113), .B(KEYINPUT55), .C1(new_n833), .C2(new_n835), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(new_n258), .B2(new_n264), .ZN(new_n844));
  INV_X1    g643(.A(new_n255), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n243), .A2(new_n244), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n230), .B1(new_n229), .B2(new_n234), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n264), .A2(new_n683), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n721), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n249), .B2(new_n257), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n843), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n264), .A2(KEYINPUT114), .A3(new_n848), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n853), .A2(new_n757), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n705), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n684), .A2(new_n266), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n708), .A2(new_n617), .A3(new_n620), .A4(new_n795), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT112), .B1(new_n860), .B2(new_n265), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n863), .A2(new_n550), .A3(new_n574), .A4(new_n773), .ZN(new_n864));
  AOI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n265), .ZN(new_n865));
  AND4_X1   g664(.A1(new_n757), .A2(new_n853), .A3(new_n854), .A4(new_n855), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n265), .A2(new_n854), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n264), .A2(new_n683), .A3(new_n848), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n757), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n621), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n862), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n571), .A2(new_n550), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n872), .A2(new_n547), .A3(new_n580), .A4(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n327), .A3(new_n266), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n865), .A2(new_n875), .ZN(G1340gat));
  AOI21_X1  g675(.A(G120gat), .B1(new_n864), .B2(new_n683), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n874), .A2(new_n328), .A3(new_n795), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1341gat));
  INV_X1    g678(.A(G127gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n880), .A3(new_n705), .ZN(new_n881));
  OAI21_X1  g680(.A(G127gat), .B1(new_n874), .B2(new_n621), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1342gat));
  NOR2_X1   g682(.A1(new_n863), .A2(new_n773), .ZN(new_n884));
  INV_X1    g683(.A(new_n574), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n500), .A2(new_n662), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT115), .Z(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n884), .A2(new_n341), .A3(new_n885), .A4(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  XOR2_X1   g689(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G134gat), .B1(new_n874), .B2(new_n708), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G1343gat));
  NAND2_X1  g694(.A1(new_n697), .A2(new_n873), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n863), .B2(new_n547), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n547), .A2(new_n897), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n839), .A2(new_n840), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n837), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n258), .B2(new_n264), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n708), .B1(new_n849), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n705), .B1(new_n903), .B2(new_n856), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n899), .B1(new_n904), .B2(new_n862), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n896), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n376), .B1(new_n906), .B2(new_n265), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n548), .A3(new_n697), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n550), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n376), .A3(new_n265), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n908), .A2(new_n911), .A3(new_n912), .A4(KEYINPUT58), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n912), .A2(KEYINPUT58), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(KEYINPUT58), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n909), .A2(G141gat), .A3(new_n550), .A4(new_n266), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n914), .B(new_n915), .C1(new_n916), .C2(new_n907), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n913), .A2(new_n917), .ZN(G1344gat));
  NAND3_X1  g717(.A1(new_n910), .A2(new_n377), .A3(new_n683), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n872), .A2(new_n899), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n903), .B1(new_n708), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n621), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n860), .A2(new_n265), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n547), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n921), .B1(new_n928), .B2(KEYINPUT57), .ZN(new_n929));
  INV_X1    g728(.A(new_n896), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n683), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n377), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n929), .A2(KEYINPUT119), .A3(new_n683), .A4(new_n930), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n920), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g734(.A(KEYINPUT59), .B(new_n377), .C1(new_n906), .C2(new_n683), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n919), .B1(new_n935), .B2(new_n936), .ZN(G1345gat));
  NAND2_X1  g736(.A1(new_n910), .A2(new_n705), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n910), .A2(KEYINPUT120), .A3(new_n705), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n621), .A2(new_n406), .ZN(new_n943));
  AOI22_X1  g742(.A1(new_n942), .A2(new_n406), .B1(new_n906), .B2(new_n943), .ZN(G1346gat));
  AND2_X1   g743(.A1(new_n906), .A2(new_n757), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n888), .A2(new_n385), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n945), .A2(new_n385), .B1(new_n909), .B2(new_n946), .ZN(G1347gat));
  NOR2_X1   g746(.A1(new_n863), .A2(new_n712), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n574), .A2(new_n500), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n252), .A3(new_n265), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT121), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n547), .B1(new_n857), .B2(new_n862), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n773), .A2(new_n955), .A3(new_n550), .A4(new_n580), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n771), .A2(new_n772), .A3(new_n550), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT122), .B1(new_n957), .B2(new_n372), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT123), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n956), .A2(new_n958), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n872), .A2(new_n961), .A3(new_n962), .A4(new_n547), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n266), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n953), .A2(new_n965), .ZN(G1348gat));
  OAI21_X1  g765(.A(G176gat), .B1(new_n964), .B2(new_n795), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n286), .A3(new_n683), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1349gat));
  NAND3_X1  g768(.A1(new_n960), .A2(new_n963), .A3(new_n705), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G183gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n705), .A2(new_n472), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  AND4_X1   g772(.A1(new_n571), .A2(new_n872), .A3(new_n949), .A4(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n971), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n977), .A2(KEYINPUT60), .A3(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT60), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n978), .B1(new_n971), .B2(new_n975), .ZN(new_n982));
  AOI211_X1 g781(.A(KEYINPUT124), .B(new_n974), .C1(new_n970), .C2(G183gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n980), .A2(new_n984), .ZN(G1350gat));
  NAND3_X1  g784(.A1(new_n960), .A2(new_n963), .A3(new_n662), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT125), .B1(new_n986), .B2(G190gat), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n986), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n951), .A2(new_n471), .A3(new_n757), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n987), .A2(new_n988), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(G1351gat));
  INV_X1    g793(.A(new_n929), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n781), .A2(new_n957), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n266), .A2(new_n254), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n781), .A2(new_n500), .A3(new_n547), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n948), .A2(new_n265), .A3(new_n1000), .ZN(new_n1001));
  AOI22_X1  g800(.A1(new_n998), .A2(new_n999), .B1(new_n254), .B2(new_n1001), .ZN(G1352gat));
  XOR2_X1   g801(.A(KEYINPUT126), .B(G204gat), .Z(new_n1003));
  NAND4_X1  g802(.A1(new_n948), .A2(new_n683), .A3(new_n1000), .A4(new_n1003), .ZN(new_n1004));
  XOR2_X1   g803(.A(new_n1004), .B(KEYINPUT62), .Z(new_n1005));
  NOR3_X1   g804(.A1(new_n995), .A2(new_n795), .A3(new_n997), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1005), .B1(new_n1006), .B2(new_n1003), .ZN(G1353gat));
  NAND3_X1  g806(.A1(new_n929), .A2(new_n705), .A3(new_n996), .ZN(new_n1008));
  OAI21_X1  g807(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1011), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n1012));
  NAND2_X1  g811(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1008), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n621), .A2(G211gat), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n948), .A2(new_n1000), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1012), .A2(new_n1014), .A3(new_n1016), .ZN(G1354gat));
  INV_X1    g816(.A(G218gat), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n708), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n948), .A2(new_n757), .A3(new_n1000), .ZN(new_n1020));
  AOI22_X1  g819(.A1(new_n998), .A2(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(G1355gat));
endmodule


