//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260;
  OR2_X1    g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0002(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT0), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n201), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n204), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n207), .B(new_n213), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G169), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT13), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(G1), .B(G13), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G97), .ZN(new_n252));
  INV_X1    g0052(.A(G232), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G226), .B2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n252), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n250), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n251), .A2(new_n260), .B1(G238), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n250), .A2(G274), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G45), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n271), .A3(new_n249), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n272), .A2(new_n273), .A3(new_n261), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n272), .B2(new_n261), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n267), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n247), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n265), .A2(new_n247), .A3(new_n276), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n246), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT14), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n278), .A2(G179), .A3(new_n279), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT76), .B1(new_n280), .B2(new_n281), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n280), .A2(KEYINPUT76), .A3(new_n281), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n282), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n215), .A2(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n211), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G50), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n211), .A2(new_n248), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n288), .B1(new_n289), .B2(new_n221), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n210), .B1(new_n204), .B2(new_n248), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT11), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT69), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT69), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(new_n261), .A3(G13), .A4(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n215), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT12), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n293), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n211), .A2(G1), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(G68), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT75), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(new_n308), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n295), .B(new_n303), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n287), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n311), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n278), .A2(new_n279), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G200), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n278), .A2(G190), .A3(new_n279), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n259), .A2(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G222), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT3), .B(G33), .ZN(new_n321));
  INV_X1    g0121(.A(G223), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(G1698), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n320), .B1(new_n221), .B2(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n251), .B1(G226), .B2(new_n264), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(G190), .A3(new_n276), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n304), .A2(G50), .A3(new_n306), .ZN(new_n327));
  OAI21_X1  g0127(.A(G20), .B1(new_n201), .B2(G50), .ZN(new_n328));
  INV_X1    g0128(.A(G150), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n328), .B1(new_n329), .B2(new_n291), .C1(new_n330), .C2(new_n289), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n293), .B1(new_n290), .B2(new_n301), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT9), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n326), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT10), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n325), .A2(new_n276), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G200), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n343), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n347));
  INV_X1    g0147(.A(new_n330), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n350), .B1(new_n211), .B2(new_n221), .C1(new_n289), .C2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n293), .B1(new_n221), .B2(new_n301), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n304), .A2(G77), .A3(new_n306), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n259), .A2(G107), .ZN(new_n356));
  INV_X1    g0156(.A(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n321), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n358), .B2(new_n253), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n259), .A2(new_n357), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(G238), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT68), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n276), .B1(new_n222), .B2(new_n263), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n355), .B1(G200), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT70), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(new_n368), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n364), .A2(new_n246), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n355), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT73), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n375), .A3(new_n355), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n364), .A2(KEYINPUT72), .A3(G179), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT72), .B1(new_n364), .B2(G179), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n374), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n334), .B1(new_n341), .B2(new_n246), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n325), .A2(new_n382), .A3(new_n276), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NOR4_X1   g0184(.A1(new_n318), .A2(new_n346), .A3(new_n380), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n293), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G58), .A2(G68), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n201), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G20), .ZN(new_n389));
  INV_X1    g0189(.A(new_n291), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G159), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(KEYINPUT77), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT77), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n211), .B1(new_n201), .B2(new_n387), .ZN(new_n394));
  INV_X1    g0194(.A(G159), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n291), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n393), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n321), .B2(G20), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n215), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n386), .B1(new_n403), .B2(KEYINPUT16), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT78), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n257), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n258), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n257), .A2(new_n406), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT7), .B(new_n211), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n215), .B1(new_n410), .B2(new_n400), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n405), .B1(new_n411), .B2(new_n398), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n330), .A2(new_n305), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n304), .A2(new_n414), .B1(new_n301), .B2(new_n330), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n322), .A2(G1698), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n257), .A3(new_n258), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT80), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n321), .A2(KEYINPUT80), .A3(new_n417), .ZN(new_n421));
  AND4_X1   g0221(.A1(G226), .A2(new_n257), .A3(new_n258), .A4(G1698), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n420), .A2(new_n421), .B1(new_n422), .B2(KEYINPUT79), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n321), .A2(G226), .A3(G1698), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT79), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n424), .A2(new_n425), .B1(G33), .B2(G87), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n363), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n263), .A2(new_n253), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n276), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G169), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n272), .A2(new_n261), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT67), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n272), .A2(new_n273), .A3(new_n261), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n428), .B1(new_n435), .B2(new_n267), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n321), .A2(KEYINPUT79), .A3(G226), .A4(G1698), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT80), .B1(new_n321), .B2(new_n417), .ZN(new_n438));
  AND4_X1   g0238(.A1(KEYINPUT80), .A2(new_n417), .A3(new_n257), .A4(new_n258), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n422), .A2(KEYINPUT79), .B1(new_n248), .B2(new_n217), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n251), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n436), .A2(new_n442), .A3(G179), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n431), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n416), .A2(KEYINPUT18), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT18), .B1(new_n416), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n415), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n404), .B2(new_n412), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT81), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n427), .A2(new_n430), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n366), .ZN(new_n452));
  INV_X1    g0252(.A(G200), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n427), .B2(new_n430), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n436), .A2(new_n442), .A3(new_n450), .A4(new_n366), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n449), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT82), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(KEYINPUT82), .B(new_n449), .C1(new_n452), .C2(new_n456), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(KEYINPUT17), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n457), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n447), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n385), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n268), .A2(G1), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(KEYINPUT5), .B2(new_n249), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT84), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n467), .B(new_n471), .C1(KEYINPUT5), .C2(new_n249), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n266), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n321), .A2(G257), .A3(G1698), .ZN(new_n475));
  INV_X1    g0275(.A(G294), .ZN(new_n476));
  OAI221_X1 g0276(.A(new_n475), .B1(new_n248), .B2(new_n476), .C1(new_n358), .C2(new_n218), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n477), .A2(new_n251), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(G264), .A3(new_n250), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT91), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT91), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n473), .A2(new_n481), .A3(G264), .A4(new_n250), .ZN(new_n482));
  AOI211_X1 g0282(.A(new_n474), .B(new_n478), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G179), .ZN(new_n484));
  INV_X1    g0284(.A(new_n474), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n477), .A2(new_n251), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n479), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G169), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n321), .A2(new_n211), .A3(G87), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT22), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n223), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n223), .A3(G20), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n494), .A2(KEYINPUT90), .B1(new_n495), .B2(G20), .ZN(new_n496));
  AOI211_X1 g0296(.A(new_n493), .B(new_n496), .C1(KEYINPUT90), .C2(new_n494), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n490), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n491), .B1(new_n497), .B2(new_n490), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n293), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n293), .B(new_n301), .C1(new_n261), .C2(G33), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT25), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n300), .B2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n223), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n501), .A2(G107), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n484), .A2(new_n488), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n487), .A2(G190), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n485), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n509), .B2(new_n453), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n500), .A2(new_n505), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n321), .A2(G257), .A3(new_n357), .ZN(new_n514));
  INV_X1    g0314(.A(G303), .ZN(new_n515));
  OAI221_X1 g0315(.A(new_n514), .B1(new_n515), .B2(new_n321), .C1(new_n323), .C2(new_n224), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n251), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n473), .A2(G270), .A3(new_n250), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n485), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n382), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n211), .C1(G33), .C2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n293), .C1(new_n211), .C2(G116), .ZN(new_n524));
  XOR2_X1   g0324(.A(new_n524), .B(KEYINPUT20), .Z(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n301), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n304), .B1(G1), .B2(new_n248), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n526), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n520), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n529), .A2(new_n519), .A3(KEYINPUT21), .A4(G169), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n529), .B1(new_n519), .B2(G200), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n366), .B2(new_n519), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n529), .A2(G169), .A3(new_n519), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT21), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n532), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n319), .A2(KEYINPUT4), .A3(G244), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n360), .A2(G250), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n521), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT4), .B1(new_n319), .B2(G244), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n251), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n473), .A2(G257), .A3(new_n250), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n543), .A2(new_n485), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n382), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n223), .A2(KEYINPUT6), .A3(G97), .ZN(new_n547));
  XOR2_X1   g0347(.A(G97), .B(G107), .Z(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(KEYINPUT6), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(G20), .B1(G77), .B2(new_n390), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n410), .A2(new_n400), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(new_n223), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n293), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n300), .A2(G97), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n501), .B2(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n543), .A2(new_n485), .A3(new_n544), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n246), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n546), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(G200), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n543), .A2(G190), .A3(new_n485), .A4(new_n544), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n560), .A2(new_n553), .A3(new_n555), .A4(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT86), .B1(new_n358), .B2(new_n216), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n360), .A2(G244), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G116), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n358), .A2(KEYINPUT86), .A3(new_n216), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n251), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n362), .A2(new_n218), .A3(new_n467), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n570), .A2(KEYINPUT85), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(KEYINPUT85), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n571), .A2(new_n572), .B1(new_n267), .B2(new_n467), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n382), .ZN(new_n575));
  NOR3_X1   g0375(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n576), .B(KEYINPUT87), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n211), .B1(new_n252), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n321), .A2(new_n211), .A3(G68), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n578), .B1(new_n289), .B2(new_n522), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT88), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(KEYINPUT88), .A3(new_n581), .A4(new_n582), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n293), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n351), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n501), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n301), .A2(new_n351), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n569), .A2(new_n573), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n246), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n575), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n386), .B1(new_n583), .B2(new_n584), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n586), .B1(new_n301), .B2(new_n351), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(G200), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT89), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n501), .A2(new_n598), .A3(G87), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT89), .B1(new_n528), .B2(new_n217), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n569), .A2(new_n573), .A3(G190), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n596), .A2(new_n597), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n513), .A2(new_n538), .A3(new_n563), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n466), .A2(new_n605), .ZN(G372));
  INV_X1    g0406(.A(new_n466), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n594), .A2(new_n603), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT92), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT26), .ZN(new_n610));
  INV_X1    g0410(.A(new_n559), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT92), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n594), .A2(new_n603), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT94), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n594), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n575), .A2(new_n591), .A3(KEYINPUT94), .A4(new_n593), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n611), .A2(new_n594), .A3(new_n603), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(KEYINPUT26), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n510), .A2(new_n511), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n609), .A2(new_n621), .A3(new_n563), .A4(new_n613), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT93), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n532), .A2(new_n623), .A3(new_n537), .ZN(new_n624));
  INV_X1    g0424(.A(new_n537), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n530), .A2(new_n531), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT93), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n506), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n614), .B(new_n620), .C1(new_n622), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n607), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n630), .B(KEYINPUT95), .Z(new_n631));
  INV_X1    g0431(.A(new_n447), .ZN(new_n632));
  INV_X1    g0432(.A(new_n312), .ZN(new_n633));
  INV_X1    g0433(.A(new_n379), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n317), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n461), .A2(new_n464), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n632), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n346), .B(KEYINPUT96), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n384), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n631), .A2(new_n640), .ZN(G369));
  NAND3_X1  g0441(.A1(new_n261), .A2(new_n211), .A3(G13), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n625), .B2(new_n626), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n500), .B2(new_n505), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT97), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n513), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n506), .A2(new_n648), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n529), .A2(new_n647), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n538), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n624), .A2(new_n627), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n658), .B2(new_n656), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n513), .A2(new_n652), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n506), .A2(new_n647), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n655), .B1(new_n660), .B2(new_n664), .ZN(G399));
  NOR2_X1   g0465(.A1(new_n577), .A2(G116), .ZN(new_n666));
  INV_X1    g0466(.A(new_n205), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(G1), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n208), .B2(new_n669), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT28), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT31), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n557), .A2(new_n592), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n520), .A3(new_n508), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT30), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT98), .B1(new_n483), .B2(new_n545), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT98), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n509), .A2(new_n678), .A3(new_n557), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n592), .A2(new_n519), .A3(new_n382), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT99), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT99), .ZN(new_n684));
  AOI211_X1 g0484(.A(new_n684), .B(new_n681), .C1(new_n677), .C2(new_n679), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n673), .B(new_n676), .C1(new_n683), .C2(new_n685), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n686), .A2(new_n647), .B1(new_n605), .B2(KEYINPUT31), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n680), .A2(new_n682), .ZN(new_n688));
  AOI211_X1 g0488(.A(new_n673), .B(new_n648), .C1(new_n676), .C2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n608), .A2(new_n559), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n618), .B1(new_n693), .B2(new_n610), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n506), .A2(new_n625), .A3(new_n626), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n622), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n609), .A2(new_n613), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n610), .B1(new_n697), .B2(new_n611), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n648), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n629), .A2(new_n648), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n692), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n672), .B1(new_n703), .B2(G1), .ZN(G364));
  INV_X1    g0504(.A(G13), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n261), .B1(new_n706), .B2(G45), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n668), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n210), .B1(G20), .B2(new_n246), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n211), .A2(new_n382), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n714), .A2(new_n366), .A3(new_n453), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n321), .B1(new_n716), .B2(new_n290), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n713), .B(KEYINPUT101), .Z(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(G190), .A3(G200), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n382), .A2(G200), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT102), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n722), .A2(new_n211), .A3(new_n366), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n720), .A2(new_n221), .B1(new_n217), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n714), .A2(new_n453), .A3(G190), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n717), .B(new_n725), .C1(G68), .C2(new_n726), .ZN(new_n727));
  NOR4_X1   g0527(.A1(new_n211), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G159), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT32), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n722), .A2(new_n211), .A3(G190), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n223), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n718), .A2(new_n366), .A3(G200), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n730), .B(new_n733), .C1(G58), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n366), .A2(G200), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n211), .B1(new_n736), .B2(new_n382), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT103), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(KEYINPUT103), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n727), .B(new_n735), .C1(new_n522), .C2(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(G311), .A2(new_n719), .B1(new_n734), .B2(G322), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n321), .B1(new_n728), .B2(G329), .ZN(new_n744));
  INV_X1    g0544(.A(G326), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n716), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT33), .B(G317), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n726), .B2(new_n747), .ZN(new_n748));
  AOI22_X1  g0548(.A1(G283), .A2(new_n731), .B1(new_n723), .B2(G303), .ZN(new_n749));
  INV_X1    g0549(.A(new_n741), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G294), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n743), .A2(new_n748), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n712), .B1(new_n742), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n711), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n321), .A2(new_n205), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT100), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(G355), .B1(new_n526), .B2(new_n667), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n244), .A2(G45), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n667), .A2(new_n321), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n269), .A2(new_n271), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n208), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n710), .B(new_n753), .C1(new_n757), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n756), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n659), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n709), .B1(new_n659), .B2(G330), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G330), .B2(new_n659), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(G396));
  AOI22_X1  g0572(.A1(new_n371), .A2(new_n379), .B1(new_n355), .B2(new_n647), .ZN(new_n773));
  AND3_X1   g0573(.A1(new_n379), .A2(new_n355), .A3(new_n647), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n701), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n629), .A2(new_n775), .A3(new_n648), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n692), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n709), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n692), .A2(new_n777), .A3(new_n778), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n711), .A2(new_n754), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n710), .B1(new_n221), .B2(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n726), .A2(G150), .B1(new_n715), .B2(G137), .ZN(new_n785));
  INV_X1    g0585(.A(new_n734), .ZN(new_n786));
  INV_X1    g0586(.A(G143), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n785), .B1(new_n786), .B2(new_n787), .C1(new_n395), .C2(new_n720), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT34), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n259), .B1(new_n728), .B2(G132), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n790), .B1(new_n724), .B2(new_n290), .C1(new_n215), .C2(new_n732), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G58), .B2(new_n750), .ZN(new_n792));
  INV_X1    g0592(.A(new_n726), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n728), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n259), .B1(new_n796), .B2(new_n797), .C1(new_n716), .C2(new_n515), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n795), .B(new_n798), .C1(G97), .C2(new_n750), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n526), .A2(new_n720), .B1(new_n786), .B2(new_n476), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n732), .A2(new_n217), .B1(new_n724), .B2(new_n223), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n789), .A2(new_n792), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n784), .B1(new_n712), .B2(new_n803), .C1(new_n775), .C2(new_n755), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n782), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G384));
  NOR2_X1   g0606(.A1(new_n706), .A2(new_n261), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT38), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n431), .A2(new_n443), .A3(new_n645), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n416), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(KEYINPUT37), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n811), .A2(new_n459), .A3(new_n460), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT37), .B1(new_n462), .B2(new_n810), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n465), .A2(new_n449), .A3(new_n645), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT106), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n465), .A2(KEYINPUT106), .A3(new_n449), .A4(new_n645), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n808), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n404), .B1(KEYINPUT16), .B2(new_n403), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n415), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n809), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n459), .A2(new_n460), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(KEYINPUT104), .B1(new_n824), .B2(KEYINPUT37), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n824), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(new_n813), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n636), .A2(new_n632), .ZN(new_n829));
  INV_X1    g0629(.A(new_n645), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n829), .A2(new_n830), .A3(new_n822), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n831), .A3(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT108), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT108), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n828), .A2(new_n831), .A3(new_n834), .A4(KEYINPUT38), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n820), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n317), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n311), .B(new_n647), .C1(new_n287), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n311), .A2(new_n647), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n282), .A2(new_n283), .ZN(new_n840));
  INV_X1    g0640(.A(new_n286), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n284), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n317), .B(new_n839), .C1(new_n842), .C2(new_n313), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n775), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n686), .A2(new_n647), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n605), .A2(KEYINPUT31), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n676), .B1(new_n683), .B2(new_n685), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n849), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n845), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n836), .A2(KEYINPUT40), .A3(new_n851), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n824), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n853), .A2(new_n825), .A3(new_n812), .ZN(new_n854));
  INV_X1    g0654(.A(new_n822), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n465), .A2(new_n645), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n808), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT105), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n832), .ZN(new_n859));
  OAI211_X1 g0659(.A(KEYINPUT105), .B(new_n808), .C1(new_n854), .C2(new_n856), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(new_n851), .A3(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT110), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT110), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n861), .A2(new_n865), .A3(new_n862), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n852), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n848), .A2(new_n850), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n607), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n867), .B1(new_n607), .B2(new_n868), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n870), .A2(new_n871), .A3(new_n691), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT111), .Z(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n634), .A2(new_n648), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n778), .A2(new_n875), .ZN(new_n876));
  AND4_X1   g0676(.A1(new_n860), .A2(new_n859), .A3(new_n844), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n447), .B2(new_n645), .ZN(new_n878));
  XNOR2_X1  g0678(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n820), .A2(new_n833), .A3(new_n835), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n859), .A2(KEYINPUT39), .A3(new_n860), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n312), .A2(new_n647), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n607), .B1(new_n700), .B2(new_n702), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n640), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n885), .B(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n807), .B1(new_n874), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n874), .B2(new_n888), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(G116), .A3(new_n212), .A4(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT36), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n209), .A2(G77), .A3(new_n387), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(G50), .B2(new_n215), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(G1), .A3(new_n705), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(new_n894), .A3(new_n897), .ZN(G367));
  NAND2_X1  g0698(.A1(new_n556), .A2(new_n647), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n563), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n611), .A2(new_n647), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n653), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT113), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n563), .A2(new_n506), .A3(new_n899), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n559), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT112), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n648), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n903), .B2(KEYINPUT42), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n596), .A2(new_n601), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n697), .B1(new_n912), .B2(new_n648), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n618), .A2(new_n911), .A3(new_n647), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n904), .A2(new_n910), .B1(KEYINPUT43), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n660), .A2(new_n664), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n900), .A2(new_n901), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n923), .A2(KEYINPUT114), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n668), .B(KEYINPUT41), .Z(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n655), .A2(new_n920), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT45), .Z(new_n928));
  NOR2_X1   g0728(.A1(new_n655), .A2(new_n920), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(new_n919), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n653), .B1(new_n663), .B2(new_n650), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(new_n660), .Z(new_n934));
  NAND2_X1  g0734(.A1(new_n703), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n703), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n926), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n707), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n918), .A2(KEYINPUT114), .A3(new_n922), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n918), .A2(new_n922), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n924), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n762), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n757), .B1(new_n205), .B2(new_n351), .C1(new_n236), .C2(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n944), .A2(new_n709), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n723), .A2(G116), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT46), .Z(new_n947));
  NOR2_X1   g0747(.A1(new_n732), .A2(new_n522), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n949), .B1(new_n786), .B2(new_n515), .C1(new_n794), .C2(new_n720), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n741), .A2(new_n223), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n321), .B1(new_n728), .B2(G317), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n793), .B2(new_n476), .C1(new_n797), .C2(new_n716), .ZN(new_n953));
  OR4_X1    g0753(.A1(new_n947), .A2(new_n950), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G50), .A2(new_n719), .B1(new_n734), .B2(G150), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G58), .A2(new_n723), .B1(new_n731), .B2(G77), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n750), .A2(G68), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n259), .B1(new_n728), .B2(G137), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n793), .B2(new_n395), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G143), .B2(new_n715), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n954), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  OAI221_X1 g0763(.A(new_n945), .B1(new_n712), .B2(new_n963), .C1(new_n915), .C2(new_n767), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n942), .A2(new_n964), .ZN(G387));
  OAI211_X1 g0765(.A(new_n666), .B(new_n268), .C1(new_n215), .C2(new_n221), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT50), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n330), .B2(G50), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n348), .A2(KEYINPUT50), .A3(new_n290), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n763), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n762), .B1(new_n233), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n759), .B1(G116), .B2(new_n577), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n205), .A2(G107), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n757), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n734), .A2(G50), .B1(G77), .B2(new_n723), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n949), .B(new_n977), .C1(new_n215), .C2(new_n720), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n741), .A2(new_n351), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n259), .B1(new_n728), .B2(G150), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n793), .B2(new_n330), .C1(new_n395), .C2(new_n716), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n734), .A2(G317), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n726), .A2(G311), .B1(new_n715), .B2(G322), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(new_n720), .C2(new_n515), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT48), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n750), .A2(G283), .B1(G294), .B2(new_n723), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT49), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n259), .B1(new_n745), .B2(new_n796), .C1(new_n732), .C2(new_n526), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n991), .B2(KEYINPUT49), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n982), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n709), .B(new_n976), .C1(new_n995), .C2(new_n712), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n664), .B2(new_n756), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n934), .B2(new_n708), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n668), .B(KEYINPUT115), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n935), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n703), .A2(new_n934), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(G393));
  INV_X1    g0802(.A(new_n999), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n932), .A2(new_n935), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT116), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT116), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n932), .A2(new_n1006), .A3(new_n935), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n936), .B(new_n1003), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n932), .A2(new_n707), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n241), .A2(new_n943), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n757), .B1(new_n522), .B2(new_n205), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n709), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n734), .A2(G159), .B1(G150), .B2(new_n715), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT51), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n321), .B1(new_n796), .B2(new_n787), .C1(new_n793), .C2(new_n290), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G87), .B2(new_n731), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n750), .A2(G77), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n719), .A2(new_n348), .B1(G68), .B2(new_n723), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n734), .A2(G311), .B1(G317), .B2(new_n715), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT52), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n321), .B1(new_n728), .B2(G322), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n793), .B2(new_n515), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n733), .A2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n719), .A2(G294), .B1(G283), .B2(new_n723), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n526), .C2(new_n741), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1014), .A2(new_n1019), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1012), .B1(new_n1027), .B2(new_n711), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n920), .B2(new_n767), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1009), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1008), .A2(new_n1030), .ZN(G390));
  NAND2_X1  g0831(.A1(new_n876), .A2(new_n844), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n883), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n880), .A2(new_n881), .A3(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n648), .B(new_n775), .C1(new_n696), .C2(new_n698), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n875), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n883), .B1(new_n1037), .B2(new_n844), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n836), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n691), .B1(new_n848), .B2(new_n850), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n845), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(G330), .B(new_n775), .C1(new_n687), .C2(new_n689), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n844), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n836), .B2(new_n1038), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT117), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1035), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1050), .B1(new_n1035), .B2(new_n1049), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1045), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n607), .A2(new_n1041), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n886), .A2(new_n640), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1048), .A2(new_n1037), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1041), .A2(new_n775), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n1047), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n876), .B1(new_n1044), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1055), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1053), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1045), .B(new_n1062), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n999), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n783), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n709), .B1(new_n348), .B2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n259), .B1(new_n796), .B2(new_n476), .C1(new_n716), .C2(new_n794), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G107), .B2(new_n726), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G68), .A2(new_n731), .B1(new_n723), .B2(G87), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G97), .A2(new_n719), .B1(new_n734), .B2(G116), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1071), .A2(new_n1017), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n715), .A2(G128), .ZN(new_n1075));
  INV_X1    g0875(.A(G125), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n321), .C1(new_n1076), .C2(new_n796), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n732), .A2(new_n290), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G132), .C2(new_n734), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n723), .A2(G150), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G159), .A2(new_n750), .B1(new_n1080), .B2(KEYINPUT53), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(KEYINPUT53), .C2(new_n1080), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT54), .B(G143), .Z(new_n1083));
  AOI22_X1  g0883(.A1(new_n719), .A2(new_n1083), .B1(G137), .B2(new_n726), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT118), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1074), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1069), .B1(new_n1086), .B2(new_n711), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n882), .B2(new_n755), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1053), .B2(new_n707), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1067), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G378));
  NOR2_X1   g0891(.A1(new_n321), .A2(G41), .ZN(new_n1092));
  AOI211_X1 g0892(.A(G50), .B(new_n1092), .C1(new_n248), .C2(new_n249), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1092), .B1(new_n794), .B2(new_n796), .C1(new_n716), .C2(new_n526), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G97), .B2(new_n726), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n734), .A2(G107), .B1(G77), .B2(new_n723), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n719), .A2(new_n588), .B1(G58), .B2(new_n731), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1095), .A2(new_n957), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT58), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1093), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G128), .A2(new_n734), .B1(new_n719), .B2(G137), .ZN(new_n1101));
  INV_X1    g0901(.A(G132), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n793), .A2(new_n1102), .B1(new_n716), .B2(new_n1076), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n723), .B2(new_n1083), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(new_n329), .C2(new_n741), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT59), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n731), .A2(G159), .ZN(new_n1107));
  AOI211_X1 g0907(.A(G33), .B(G41), .C1(new_n728), .C2(G124), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1105), .A2(KEYINPUT59), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1100), .B1(new_n1099), .B2(new_n1098), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n711), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n710), .B1(new_n290), .B2(new_n783), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n384), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n639), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n334), .A2(new_n645), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1115), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1121), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n1119), .A3(new_n1114), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1112), .B(new_n1113), .C1(new_n1125), .C2(new_n755), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n836), .A2(KEYINPUT40), .A3(new_n851), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n861), .A2(new_n865), .A3(new_n862), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n865), .B1(new_n861), .B2(new_n862), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n1128), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1125), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n864), .A2(new_n866), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(G330), .A3(new_n1128), .A4(new_n1125), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT119), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n878), .B2(new_n884), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1127), .B1(new_n1141), .B2(new_n708), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1055), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1065), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT120), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1065), .A2(new_n1143), .A3(KEYINPUT120), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT57), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1125), .B1(new_n867), .B2(G330), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n885), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1133), .A2(new_n1135), .A3(new_n884), .A4(new_n878), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1003), .B1(new_n1148), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT57), .B1(new_n1148), .B2(new_n1141), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT121), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(KEYINPUT121), .B(KEYINPUT57), .C1(new_n1148), .C2(new_n1141), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1142), .B1(new_n1158), .B2(new_n1159), .ZN(G375));
  NAND2_X1  g0960(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n708), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1162), .A2(KEYINPUT122), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1047), .A2(new_n754), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n709), .B1(G68), .B2(new_n1068), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n259), .B1(new_n796), .B2(new_n515), .C1(new_n716), .C2(new_n476), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G116), .B2(new_n726), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n979), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G77), .A2(new_n731), .B1(new_n723), .B2(G97), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G107), .A2(new_n719), .B1(new_n734), .B2(G283), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n716), .A2(new_n1102), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n259), .B(new_n1172), .C1(new_n726), .C2(new_n1083), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n719), .A2(G150), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n734), .A2(G137), .B1(G58), .B2(new_n731), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n750), .A2(G50), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n723), .A2(G159), .B1(G128), .B2(new_n728), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT123), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1171), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1165), .B1(new_n1180), .B2(new_n711), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1162), .A2(KEYINPUT122), .B1(new_n1164), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1163), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1161), .A2(new_n1143), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1063), .A2(new_n926), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(G381));
  AND3_X1   g0986(.A1(new_n1065), .A2(new_n1143), .A3(KEYINPUT120), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT120), .B1(new_n1065), .B2(new_n1143), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1140), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1138), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1149), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT121), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n1155), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n1090), .A3(new_n1142), .ZN(new_n1196));
  OR4_X1    g0996(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1197));
  OR4_X1    g0997(.A1(G387), .A2(new_n1196), .A3(G381), .A4(new_n1197), .ZN(G407));
  OAI211_X1 g0998(.A(G407), .B(G213), .C1(G343), .C2(new_n1196), .ZN(G409));
  NAND2_X1  g0999(.A1(new_n646), .A2(G213), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(G378), .B(new_n1142), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1189), .A2(new_n1191), .A3(new_n925), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1126), .B1(new_n1204), .B2(new_n707), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1090), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1201), .B1(new_n1202), .B2(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1184), .A2(KEYINPUT60), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1184), .A2(KEYINPUT60), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1208), .A2(new_n999), .A3(new_n1063), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1183), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(new_n805), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n805), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1207), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT63), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1201), .A2(G2897), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1215), .B(new_n1221), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1207), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1207), .A2(KEYINPUT63), .A3(new_n1216), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(G393), .B(new_n771), .ZN(new_n1225));
  OR3_X1    g1025(.A1(new_n1008), .A2(new_n1030), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1008), .B2(new_n1030), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n964), .A3(new_n942), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1226), .A2(new_n1227), .B1(new_n964), .B2(new_n942), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1229), .A2(KEYINPUT61), .A3(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1219), .A2(new_n1223), .A3(new_n1224), .A4(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT62), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1207), .A2(new_n1233), .A3(new_n1216), .ZN(new_n1234));
  XOR2_X1   g1034(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1207), .B2(new_n1222), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1207), .B2(new_n1216), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT125), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1230), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(KEYINPUT125), .A3(new_n1228), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1232), .B1(new_n1238), .B2(new_n1243), .ZN(G405));
  NAND2_X1  g1044(.A1(G375), .A2(new_n1090), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1245), .A2(new_n1202), .A3(new_n1215), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1215), .B1(new_n1245), .B2(new_n1202), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1243), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT127), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1243), .B(KEYINPUT127), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1202), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G378), .B1(new_n1195), .B2(new_n1142), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1216), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1245), .A2(new_n1202), .A3(new_n1215), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1254), .A2(new_n1255), .A3(KEYINPUT126), .A4(new_n1256), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1250), .A2(new_n1251), .B1(new_n1259), .B2(new_n1260), .ZN(G402));
endmodule


