//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  AND2_X1   g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n203), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n206), .B1(new_n209), .B2(new_n210), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G68), .B(G77), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XOR2_X1   g0035(.A(G50), .B(G58), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  XOR2_X1   g0041(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g0043(.A1(G226), .A2(G1698), .ZN(new_n244));
  AOI21_X1  g0044(.A(new_n244), .B1(new_n219), .B2(G1698), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n245), .A2(new_n250), .B1(G33), .B2(G97), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n207), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n256), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n253), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n251), .A2(new_n253), .B1(new_n213), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n207), .B2(new_n252), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n265), .A2(KEYINPUT71), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT71), .B1(new_n265), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n243), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n253), .A2(G274), .A3(new_n266), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT71), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n265), .A2(KEYINPUT71), .A3(new_n266), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G1), .A2(G13), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT66), .B(G1), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n256), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G238), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G97), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n219), .A2(G1698), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G226), .B2(G1698), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n282), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n278), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n275), .A2(new_n281), .A3(new_n289), .A4(new_n242), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n270), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT14), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT73), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(G238), .A2(new_n280), .B1(new_n288), .B2(new_n278), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n296), .A2(KEYINPUT73), .A3(new_n242), .A4(new_n275), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT13), .B1(new_n263), .B2(new_n269), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n295), .A2(new_n297), .A3(G179), .A4(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT14), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n291), .A2(new_n300), .A3(G169), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n293), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT12), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n258), .A2(new_n260), .A3(G13), .A4(G20), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n305), .B2(new_n212), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n304), .A2(KEYINPUT12), .A3(G68), .ZN(new_n307));
  NAND3_X1  g0107(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n277), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT68), .B1(new_n247), .B2(G20), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT68), .ZN(new_n312));
  INV_X1    g0112(.A(G20), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(G33), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n314), .A3(G77), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G20), .A2(G33), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(G50), .B1(G20), .B2(new_n212), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n310), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n306), .A2(new_n307), .B1(KEYINPUT11), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n304), .A2(new_n310), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n258), .A2(new_n260), .A3(G20), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(G68), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(KEYINPUT11), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n302), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n291), .A2(G200), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n295), .A2(new_n297), .A3(G190), .A4(new_n298), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n325), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT74), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT16), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n248), .A2(new_n313), .A3(new_n249), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n313), .A4(new_n249), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n212), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(G58), .A2(G68), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G58), .A2(G68), .ZN(new_n340));
  OAI21_X1  g0140(.A(G20), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n316), .A2(G159), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n333), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT76), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT76), .B(new_n333), .C1(new_n338), .C2(new_n343), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT7), .B1(new_n287), .B2(new_n313), .ZN(new_n348));
  INV_X1    g0148(.A(new_n337), .ZN(new_n349));
  OAI21_X1  g0149(.A(G68), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT75), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n341), .B2(new_n342), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n341), .A2(new_n351), .A3(new_n342), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n350), .B(KEYINPUT16), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n346), .A2(new_n347), .A3(new_n309), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n218), .A2(KEYINPUT8), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT8), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G58), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n305), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n321), .A2(KEYINPUT77), .A3(new_n359), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n310), .A3(new_n304), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT77), .B1(new_n321), .B2(new_n359), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT78), .B(new_n361), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n321), .A2(new_n359), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n320), .A3(new_n362), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT78), .B1(new_n370), .B2(new_n361), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n355), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n271), .ZN(new_n374));
  INV_X1    g0174(.A(G223), .ZN(new_n375));
  INV_X1    g0175(.A(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G226), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G1698), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n377), .B(new_n379), .C1(new_n285), .C2(new_n286), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n247), .A2(new_n214), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n253), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n261), .A2(G232), .A3(new_n253), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT80), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n261), .A2(KEYINPUT80), .A3(G232), .A4(new_n253), .ZN(new_n387));
  AOI211_X1 g0187(.A(new_n374), .B(new_n383), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n271), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT79), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G223), .A2(G1698), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n378), .B2(G1698), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n381), .B1(new_n393), .B2(new_n250), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n391), .B1(new_n394), .B2(new_n253), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n383), .A2(KEYINPUT79), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n388), .A2(G169), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n373), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT18), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n399), .B1(new_n355), .B2(new_n372), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G190), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n407), .A2(KEYINPUT81), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(KEYINPUT81), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n395), .A2(new_n396), .A3(new_n410), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n388), .A2(G200), .B1(new_n390), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n355), .A2(new_n412), .A3(new_n372), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n355), .A2(new_n412), .A3(KEYINPUT17), .A4(new_n372), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n406), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n250), .A2(G222), .A3(new_n376), .ZN(new_n419));
  INV_X1    g0219(.A(G77), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n250), .A2(G1698), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT67), .B(G223), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n419), .B1(new_n420), .B2(new_n250), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n278), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n374), .B1(new_n280), .B2(G226), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT9), .ZN(new_n428));
  NOR2_X1   g0228(.A1(G50), .A2(G58), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n313), .B1(new_n429), .B2(new_n212), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT69), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n311), .A2(new_n314), .ZN(new_n432));
  INV_X1    g0232(.A(G150), .ZN(new_n433));
  INV_X1    g0233(.A(new_n316), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n360), .A2(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n309), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G50), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n309), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n305), .A2(new_n437), .B1(new_n438), .B2(new_n321), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n427), .A2(G190), .B1(new_n428), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n440), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(KEYINPUT9), .B1(new_n426), .B2(G200), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT10), .ZN(new_n445));
  INV_X1    g0245(.A(G169), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n442), .B1(new_n426), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(G179), .B2(new_n426), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n360), .A2(new_n434), .B1(new_n313), .B2(new_n420), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT15), .B(G87), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n432), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n309), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n320), .A2(G77), .A3(new_n321), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n305), .A2(new_n420), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT70), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT70), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n452), .A2(new_n457), .A3(new_n453), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n250), .A2(G232), .A3(new_n376), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n287), .A2(G107), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(new_n421), .C2(new_n213), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n278), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n374), .B1(new_n280), .B2(G244), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n446), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n397), .A3(new_n464), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(G200), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n463), .A2(G190), .A3(new_n464), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n456), .A2(new_n469), .A3(new_n458), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n418), .A2(new_n445), .A3(new_n448), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n332), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n476), .A2(new_n220), .A3(G107), .ZN(new_n477));
  XNOR2_X1  g0277(.A(G97), .B(G107), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n479), .A2(new_n313), .B1(new_n420), .B2(new_n434), .ZN(new_n480));
  INV_X1    g0280(.A(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n336), .B2(new_n337), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n309), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n305), .A2(new_n220), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n279), .A2(G33), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n485), .A2(G97), .A3(new_n310), .A4(new_n304), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G250), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT82), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(new_n376), .C1(new_n285), .C2(new_n286), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n376), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n278), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g0296(.A(KEYINPUT5), .B(G41), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n279), .A2(new_n497), .A3(G45), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G257), .A3(new_n253), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n265), .A2(new_n279), .A3(new_n497), .A4(G45), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n502), .A3(new_n397), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n490), .A2(new_n491), .B1(G33), .B2(G283), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT82), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n488), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n488), .A2(new_n505), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n504), .B(new_n493), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n501), .B1(new_n508), .B2(new_n278), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n487), .B(new_n503), .C1(G169), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n486), .A2(new_n484), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n220), .A2(new_n481), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n476), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n477), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G20), .B1(G77), .B2(new_n316), .ZN(new_n517));
  OAI21_X1  g0317(.A(G107), .B1(new_n348), .B2(new_n349), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n511), .B1(new_n519), .B2(new_n309), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n496), .A2(new_n502), .A3(G190), .ZN(new_n521));
  INV_X1    g0321(.A(G200), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n521), .C1(new_n522), .C2(new_n509), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n510), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n258), .A2(new_n260), .A3(G45), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n525), .A2(new_n278), .A3(new_n264), .ZN(new_n526));
  OAI211_X1 g0326(.A(G238), .B(new_n376), .C1(new_n285), .C2(new_n286), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G116), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n526), .B1(new_n278), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT83), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n279), .A2(new_n533), .A3(G45), .ZN(new_n534));
  OAI21_X1  g0334(.A(G250), .B1(new_n276), .B2(new_n277), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(KEYINPUT84), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT84), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n535), .B1(KEYINPUT83), .B2(new_n525), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(new_n534), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n531), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n311), .A2(new_n314), .A3(G97), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n313), .B(G68), .C1(new_n285), .C2(new_n286), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n313), .B1(new_n282), .B2(new_n545), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n513), .A2(new_n214), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n309), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n305), .A2(new_n450), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n320), .A2(G87), .A3(new_n485), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n543), .A2(KEYINPUT85), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT85), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n537), .A2(KEYINPUT84), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n540), .A2(new_n539), .A3(new_n534), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n522), .B1(new_n561), .B2(new_n531), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n558), .B1(new_n562), .B2(new_n555), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(G190), .A3(new_n531), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT86), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n561), .A2(KEYINPUT86), .A3(G190), .A4(new_n531), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n557), .A2(new_n563), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n551), .A2(new_n309), .B1(new_n305), .B2(new_n450), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n320), .A2(new_n485), .ZN(new_n570));
  INV_X1    g0370(.A(new_n450), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n542), .A2(new_n446), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n561), .A2(new_n397), .A3(new_n531), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n524), .A2(new_n568), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n313), .B(G87), .C1(new_n285), .C2(new_n286), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT22), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n250), .A2(new_n579), .A3(new_n313), .A4(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT90), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n529), .B2(G20), .ZN(new_n584));
  OR3_X1    g0384(.A1(new_n313), .A2(KEYINPUT23), .A3(G107), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n313), .A2(KEYINPUT90), .A3(G33), .A4(G116), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT23), .B1(new_n313), .B2(G107), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n581), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n582), .B1(new_n581), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n309), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n481), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT25), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n304), .B2(G107), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n570), .A2(G107), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n215), .A2(new_n376), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n221), .A2(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n285), .C2(new_n286), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G294), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT91), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(KEYINPUT91), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(KEYINPUT5), .A2(G41), .ZN(new_n605));
  NOR2_X1   g0405(.A1(KEYINPUT5), .A2(G41), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(G264), .B(new_n253), .C1(new_n525), .C2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT92), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n498), .A2(KEYINPUT92), .A3(G264), .A4(new_n253), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n604), .A2(new_n278), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(G200), .B1(new_n612), .B2(new_n500), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n253), .B1(new_n602), .B2(new_n603), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(new_n500), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n614), .A2(G190), .A3(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n591), .B(new_n595), .C1(new_n613), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n591), .A2(new_n595), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n610), .A2(new_n611), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n598), .A2(KEYINPUT91), .A3(new_n599), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT91), .B1(new_n598), .B2(new_n599), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n278), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n619), .A2(new_n622), .A3(G179), .A4(new_n500), .ZN(new_n623));
  OAI21_X1  g0423(.A(G169), .B1(new_n614), .B2(new_n615), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n320), .A2(G116), .A3(new_n485), .ZN(new_n628));
  INV_X1    g0428(.A(G116), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n305), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n494), .B(new_n313), .C1(G33), .C2(new_n220), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(G20), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n309), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT20), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n628), .B(new_n630), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(G270), .B(new_n253), .C1(new_n525), .C2(new_n607), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n500), .ZN(new_n639));
  OAI211_X1 g0439(.A(G257), .B(new_n376), .C1(new_n285), .C2(new_n286), .ZN(new_n640));
  INV_X1    g0440(.A(G303), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n285), .A2(new_n286), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT87), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n250), .A2(KEYINPUT87), .A3(G257), .A4(new_n376), .ZN(new_n645));
  OAI211_X1 g0445(.A(G264), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT88), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT88), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n250), .A2(new_n648), .A3(G264), .A4(G1698), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n644), .A2(new_n645), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n639), .B1(new_n650), .B2(new_n278), .ZN(new_n651));
  NAND2_X1  g0451(.A1(KEYINPUT21), .A2(G169), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI211_X1 g0453(.A(new_n397), .B(new_n639), .C1(new_n650), .C2(new_n278), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n637), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n410), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n637), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n657), .B(new_n658), .C1(new_n522), .C2(new_n651), .ZN(new_n659));
  XOR2_X1   g0459(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n660));
  NAND2_X1  g0460(.A1(new_n637), .A2(G169), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n651), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n655), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NOR4_X1   g0463(.A1(new_n475), .A2(new_n576), .A3(new_n627), .A4(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n299), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n300), .B1(new_n291), .B2(G169), .ZN(new_n666));
  AOI211_X1 g0466(.A(KEYINPUT14), .B(new_n446), .C1(new_n270), .C2(new_n290), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n330), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n668), .A2(new_n325), .B1(new_n669), .B2(new_n468), .ZN(new_n670));
  INV_X1    g0470(.A(new_n417), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n406), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n445), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n448), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT94), .Z(new_n675));
  INV_X1    g0475(.A(new_n510), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n568), .A2(KEYINPUT26), .A3(new_n676), .A4(new_n575), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n555), .B1(new_n542), .B2(G200), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n564), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n575), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n655), .A2(new_n662), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT93), .B1(new_n618), .B2(new_n625), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n591), .A2(new_n595), .B1(new_n623), .B2(new_n624), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT93), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n684), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n678), .A2(new_n564), .B1(new_n573), .B2(new_n574), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n524), .A2(new_n617), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n575), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n474), .B1(new_n683), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n675), .A2(new_n693), .ZN(G369));
  AND2_X1   g0494(.A1(new_n313), .A2(G13), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n279), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  OAI21_X1  g0497(.A(G213), .B1(new_n696), .B2(KEYINPUT27), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n658), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n684), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n663), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n700), .B1(new_n591), .B2(new_n595), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n627), .A2(new_n706), .B1(new_n626), .B2(new_n700), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n618), .A2(new_n625), .A3(KEYINPUT93), .ZN(new_n709));
  INV_X1    g0509(.A(new_n700), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n709), .A2(new_n685), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n619), .A2(new_n622), .A3(new_n500), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n614), .A2(new_n615), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n522), .A2(new_n712), .B1(new_n713), .B2(new_n407), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n618), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n687), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n651), .A2(G179), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n651), .B2(new_n652), .ZN(new_n718));
  INV_X1    g0518(.A(new_n651), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(G169), .A3(new_n637), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n718), .A2(new_n637), .B1(new_n720), .B2(new_n660), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n710), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n711), .B1(new_n716), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n708), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n204), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n549), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n210), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT98), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n627), .A2(new_n663), .A3(new_n710), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n524), .A2(new_n568), .A3(new_n575), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n619), .A2(new_n622), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT96), .B1(new_n542), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT96), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n612), .A2(new_n737), .A3(new_n561), .A4(new_n531), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n736), .A2(new_n738), .A3(new_n509), .A4(new_n654), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n509), .A2(KEYINPUT30), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n736), .A3(new_n738), .A4(new_n654), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n509), .A2(new_n651), .A3(G179), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n542), .A2(KEYINPUT97), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n542), .A2(KEYINPUT97), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n744), .A2(new_n745), .A3(new_n712), .A4(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n741), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT95), .B(KEYINPUT31), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n700), .A2(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n733), .A2(new_n734), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n739), .A2(new_n740), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n747), .A2(new_n743), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n710), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT31), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n732), .B1(new_n757), .B2(G330), .ZN(new_n758));
  INV_X1    g0558(.A(G330), .ZN(new_n759));
  AOI211_X1 g0559(.A(KEYINPUT98), .B(new_n759), .C1(new_n751), .C2(new_n756), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n575), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n680), .B2(KEYINPUT26), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n626), .A2(new_n655), .A3(new_n662), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n524), .A2(new_n764), .A3(new_n617), .A4(new_n690), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n568), .A2(new_n681), .A3(new_n676), .A4(new_n575), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(KEYINPUT29), .A3(new_n700), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n679), .A2(new_n575), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n510), .A2(new_n523), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n769), .A2(new_n770), .A3(new_n715), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n721), .B1(new_n709), .B2(new_n685), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n762), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n677), .A2(new_n682), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n710), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n768), .B1(new_n775), .B2(KEYINPUT29), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n761), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n731), .B1(new_n777), .B2(G1), .ZN(G364));
  AOI21_X1  g0578(.A(new_n257), .B1(new_n695), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n726), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n703), .A2(G330), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n705), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT99), .Z(new_n784));
  INV_X1    g0584(.A(new_n781), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n277), .B1(G20), .B2(new_n446), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(G20), .A2(G179), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n522), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n410), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n407), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n313), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n792), .A2(new_n437), .B1(new_n220), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n313), .A2(G179), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G159), .ZN(new_n800));
  INV_X1    g0600(.A(new_n788), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n797), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n800), .A2(KEYINPUT32), .B1(new_n420), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n796), .A2(G190), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n214), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n287), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT101), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n656), .A2(new_n522), .A3(new_n801), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n790), .A2(G190), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n810), .A2(G58), .B1(G68), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n796), .A2(new_n407), .A3(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n481), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n800), .B2(KEYINPUT32), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n804), .A2(new_n808), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n794), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n810), .A2(G322), .B1(G294), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n813), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n791), .A2(G326), .B1(G283), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n802), .A2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n250), .B(new_n822), .C1(G329), .C2(new_n799), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT33), .B(G317), .ZN(new_n824));
  INV_X1    g0624(.A(new_n805), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n811), .A2(new_n824), .B1(new_n825), .B2(G303), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n818), .A2(new_n820), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n787), .B1(new_n816), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G13), .A2(G33), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(G20), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n786), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n237), .A2(G45), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n725), .A2(new_n250), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n833), .B(new_n834), .C1(G45), .C2(new_n210), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n725), .A2(new_n287), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n836), .A2(G355), .B1(new_n629), .B2(new_n725), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT100), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n785), .B(new_n828), .C1(new_n832), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n831), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n703), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n784), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT102), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  AOI21_X1  g0645(.A(new_n700), .B1(new_n456), .B2(new_n458), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n471), .B1(new_n846), .B2(KEYINPUT105), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT105), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n848), .B(new_n700), .C1(new_n456), .C2(new_n458), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n468), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n850), .A2(new_n468), .A3(new_n700), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n683), .B2(new_n692), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n468), .A2(new_n710), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n846), .A2(KEYINPUT105), .ZN(new_n855));
  INV_X1    g0655(.A(new_n849), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n471), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n854), .B1(new_n857), .B2(new_n468), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n853), .B1(new_n775), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n781), .B1(new_n761), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n761), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n786), .A2(new_n829), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n785), .B1(new_n420), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n287), .B1(new_n799), .B2(G132), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n212), .B2(new_n813), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n794), .A2(new_n218), .B1(new_n805), .B2(new_n437), .ZN(new_n866));
  INV_X1    g0666(.A(new_n802), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n811), .A2(G150), .B1(G159), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(G137), .ZN(new_n869));
  XNOR2_X1  g0669(.A(KEYINPUT103), .B(G143), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n868), .B1(new_n792), .B2(new_n869), .C1(new_n809), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT34), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n865), .B(new_n866), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n813), .A2(new_n214), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(G107), .B2(new_n825), .ZN(new_n876));
  INV_X1    g0676(.A(G283), .ZN(new_n877));
  INV_X1    g0677(.A(new_n811), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .C1(new_n641), .C2(new_n792), .ZN(new_n879));
  INV_X1    g0679(.A(G294), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n809), .A2(new_n880), .B1(new_n220), .B2(new_n794), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n287), .B1(new_n802), .B2(new_n629), .C1(new_n821), .C2(new_n798), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n874), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n885), .A2(KEYINPUT104), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n786), .B1(new_n885), .B2(KEYINPUT104), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n863), .B1(new_n858), .B2(new_n830), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n861), .A2(new_n888), .ZN(G384));
  NOR2_X1   g0689(.A1(new_n279), .A2(new_n695), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n326), .A2(new_n710), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n330), .B(new_n891), .C1(new_n668), .C2(new_n325), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n326), .B(new_n710), .C1(new_n302), .C2(new_n669), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n858), .ZN(new_n895));
  INV_X1    g0695(.A(new_n753), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n700), .B1(new_n896), .B2(new_n741), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n897), .A2(KEYINPUT31), .B1(new_n734), .B2(new_n733), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n754), .A2(new_n749), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n373), .A2(new_n699), .ZN(new_n901));
  XNOR2_X1  g0701(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n401), .A2(new_n901), .A3(new_n413), .A4(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n355), .A2(new_n412), .A3(new_n372), .ZN(new_n904));
  INV_X1    g0704(.A(new_n699), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n370), .A2(new_n361), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n353), .A2(new_n352), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n333), .B1(new_n907), .B2(new_n338), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n354), .A3(new_n309), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n399), .A2(new_n905), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT107), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n905), .B1(new_n909), .B2(new_n906), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n406), .B2(new_n417), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n911), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT107), .B1(new_n903), .B2(new_n911), .ZN(new_n921));
  OAI211_X1 g0721(.A(KEYINPUT38), .B(new_n918), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n900), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n854), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n850), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n892), .B2(new_n893), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n716), .A2(new_n721), .A3(new_n659), .A4(new_n700), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n754), .A2(new_n755), .B1(new_n930), .B2(new_n576), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n754), .A2(new_n749), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT110), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n902), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n401), .A2(new_n901), .A3(new_n413), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n904), .A2(new_n403), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n905), .B1(new_n355), .B2(new_n372), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n936), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n936), .A2(new_n937), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n417), .A2(new_n942), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n373), .A2(new_n400), .A3(new_n404), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n404), .B1(new_n373), .B2(new_n400), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n415), .A2(KEYINPUT109), .A3(new_n416), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n941), .B1(new_n948), .B2(new_n939), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n922), .B1(new_n949), .B2(KEYINPUT38), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n733), .A2(new_n734), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n899), .B(new_n951), .C1(new_n755), .C2(new_n754), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(KEYINPUT110), .A3(new_n929), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n935), .A2(KEYINPUT40), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n926), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT111), .ZN(new_n956));
  INV_X1    g0756(.A(new_n952), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n475), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n759), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT112), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n851), .B1(new_n773), .B2(new_n774), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n894), .B1(new_n962), .B2(new_n854), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT38), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n966), .B2(new_n922), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n946), .A2(new_n699), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT108), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n894), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n853), .B2(new_n927), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n919), .B2(new_n923), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT108), .ZN(new_n973));
  INV_X1    g0773(.A(new_n968), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT39), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n950), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n327), .A2(new_n710), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n966), .A2(KEYINPUT39), .A3(new_n922), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n969), .A2(new_n975), .A3(new_n980), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n474), .B(new_n768), .C1(new_n775), .C2(KEYINPUT29), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n675), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n981), .B(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n890), .B1(new_n961), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n961), .B2(new_n984), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n988));
  NOR4_X1   g0788(.A1(new_n987), .A2(new_n988), .A3(new_n629), .A4(new_n209), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT36), .ZN(new_n990));
  OAI21_X1  g0790(.A(G77), .B1(new_n218), .B2(new_n212), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n991), .A2(new_n210), .B1(G50), .B2(new_n212), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n279), .A2(G13), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n986), .A2(new_n994), .ZN(G367));
  INV_X1    g0795(.A(new_n834), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n832), .B1(new_n204), .B2(new_n450), .C1(new_n232), .C2(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n997), .A2(new_n781), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n556), .A2(new_n700), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n762), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n769), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n813), .A2(new_n420), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n810), .B2(G150), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n870), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n791), .A2(new_n1004), .B1(new_n817), .B2(G68), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n250), .B1(new_n798), .B2(new_n869), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G50), .B2(new_n867), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n811), .A2(G159), .B1(new_n825), .B2(G58), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(new_n1005), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n813), .A2(new_n220), .ZN(new_n1010));
  INV_X1    g0810(.A(G317), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n287), .B1(new_n802), .B2(new_n877), .C1(new_n1011), .C2(new_n798), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G294), .C2(new_n811), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n810), .A2(G303), .B1(G107), .B2(new_n817), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n821), .C2(new_n792), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n805), .A2(new_n629), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT46), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1009), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT47), .Z(new_n1019));
  OAI221_X1 g0819(.A(new_n998), .B1(new_n841), .B2(new_n1001), .C1(new_n1019), .C2(new_n787), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n524), .B1(new_n520), .B2(new_n700), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n676), .A2(new_n710), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n723), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT45), .Z(new_n1025));
  NOR2_X1   g0825(.A1(new_n723), .A2(new_n1023), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT44), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(new_n708), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n722), .A2(new_n716), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n707), .B2(new_n722), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(new_n704), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n777), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n777), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n726), .B(KEYINPUT41), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n780), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1021), .A2(new_n626), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n710), .B1(new_n1038), .B2(new_n510), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1023), .A2(new_n716), .A3(new_n722), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(KEYINPUT42), .B2(new_n1040), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(KEYINPUT42), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1041), .A2(new_n1042), .B1(KEYINPUT43), .B2(new_n1001), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n708), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1020), .B1(new_n1037), .B2(new_n1047), .ZN(G387));
  NAND2_X1  g0848(.A1(new_n1033), .A2(new_n780), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n809), .A2(new_n1011), .B1(new_n641), .B2(new_n802), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT115), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n791), .A2(G322), .B1(new_n811), .B2(G311), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT116), .Z(new_n1053));
  AND2_X1   g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT48), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(KEYINPUT48), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n817), .A2(G283), .B1(new_n825), .B2(G294), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT117), .Z(new_n1059));
  OR2_X1    g0859(.A1(new_n1059), .A2(KEYINPUT49), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(KEYINPUT49), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n813), .A2(new_n629), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n250), .B(new_n1062), .C1(G326), .C2(new_n799), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n805), .A2(new_n420), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n791), .B2(G159), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n360), .B2(new_n878), .C1(new_n437), .C2(new_n809), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n250), .B1(new_n802), .B2(new_n212), .C1(new_n433), .C2(new_n798), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n794), .A2(new_n450), .ZN(new_n1069));
  NOR4_X1   g0869(.A1(new_n1067), .A2(new_n1010), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT114), .Z(new_n1071));
  AOI21_X1  g0871(.A(new_n787), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n728), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1073), .A2(new_n836), .B1(new_n481), .B2(new_n725), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n229), .A2(new_n255), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n360), .B2(G50), .ZN(new_n1077));
  AOI21_X1  g0877(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n728), .A3(new_n1078), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n360), .A2(new_n1076), .A3(G50), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n834), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1074), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n785), .B1(new_n1082), .B2(new_n832), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n707), .B2(new_n841), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n777), .A2(new_n1033), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n726), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n777), .A2(new_n1033), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1049), .B1(new_n1072), .B2(new_n1084), .C1(new_n1086), .C2(new_n1087), .ZN(G393));
  INV_X1    g0888(.A(new_n1029), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1085), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n726), .A3(new_n1034), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1021), .A2(new_n831), .A3(new_n1022), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n832), .B1(new_n220), .B2(new_n204), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n240), .B2(new_n834), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n821), .A2(new_n809), .B1(new_n792), .B2(new_n1011), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n878), .A2(new_n641), .B1(new_n629), .B2(new_n794), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n814), .B(new_n1097), .C1(G283), .C2(new_n825), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n287), .B1(new_n802), .B2(new_n880), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G322), .B2(new_n799), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n287), .B(new_n875), .C1(new_n799), .C2(new_n1004), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n817), .A2(G77), .B1(new_n825), .B2(G68), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n810), .A2(G159), .B1(new_n791), .B2(G150), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1102), .B(new_n1103), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n878), .A2(new_n437), .B1(new_n802), .B2(new_n360), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT119), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1109), .A2(KEYINPUT119), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1101), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n785), .B(new_n1094), .C1(new_n1113), .C2(new_n786), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1029), .A2(new_n780), .B1(new_n1092), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1091), .A2(new_n1115), .ZN(G390));
  NAND2_X1  g0916(.A1(new_n977), .A2(new_n979), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n978), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n963), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n767), .A2(new_n700), .A3(new_n858), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n927), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n894), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n950), .A3(new_n1118), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n858), .B(new_n894), .C1(new_n758), .C2(new_n760), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n952), .A2(G330), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n895), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n977), .A2(new_n979), .B1(new_n963), .B2(new_n1118), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1124), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n830), .B1(new_n977), .B2(new_n979), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n791), .A2(G128), .B1(G50), .B2(new_n819), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n869), .B2(new_n878), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n810), .A2(G132), .B1(G159), .B2(new_n817), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n287), .B1(new_n799), .B2(G125), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n1138), .C1(new_n802), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT53), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n805), .B2(new_n433), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n825), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1136), .B(new_n1140), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n791), .A2(G283), .B1(new_n811), .B2(G107), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n420), .B2(new_n794), .C1(new_n629), .C2(new_n809), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n813), .A2(new_n212), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n287), .B1(new_n802), .B2(new_n220), .C1(new_n880), .C2(new_n798), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1146), .A2(new_n806), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n786), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n862), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n781), .C1(new_n359), .C2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1134), .A2(new_n1152), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(KEYINPUT121), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT121), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1133), .A2(new_n780), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT120), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n952), .A2(G330), .A3(new_n858), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1122), .B1(new_n1158), .B2(new_n970), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1125), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n858), .B1(new_n758), .B2(new_n760), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1128), .B1(new_n1161), .B2(new_n970), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n962), .A2(new_n854), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n474), .A2(G330), .A3(new_n952), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n675), .A2(new_n982), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1157), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n726), .B1(new_n1168), .B2(new_n1132), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1170), .A2(KEYINPUT120), .A3(new_n1132), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1156), .B1(new_n1169), .B2(new_n1171), .ZN(G378));
  NAND3_X1  g0972(.A1(new_n926), .A2(new_n954), .A3(G330), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n445), .A2(new_n448), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n440), .A2(new_n699), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT55), .Z(new_n1176));
  AND2_X1   g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OR3_X1    g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1173), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n759), .B1(new_n924), .B2(new_n925), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n954), .A3(new_n1183), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1185), .A2(new_n1188), .A3(new_n975), .A4(new_n1190), .ZN(new_n1191));
  AND4_X1   g0991(.A1(G330), .A2(new_n926), .A3(new_n954), .A4(new_n1183), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1183), .B1(new_n1189), .B2(new_n954), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n981), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1184), .A2(new_n829), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n781), .B1(G50), .B2(new_n1151), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n250), .A2(G41), .ZN(new_n1198));
  AOI211_X1 g0998(.A(G50), .B(new_n1198), .C1(new_n247), .C2(new_n254), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1198), .B1(new_n877), .B2(new_n798), .C1(new_n450), .C2(new_n802), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1065), .B(new_n1200), .C1(G68), .C2(new_n817), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n791), .A2(G116), .B1(G58), .B2(new_n819), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n810), .A2(G107), .B1(G97), .B2(new_n811), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT58), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n810), .A2(G128), .B1(G132), .B2(new_n811), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n817), .A2(G150), .B1(G137), .B2(new_n867), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1139), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n791), .A2(G125), .B1(new_n825), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n819), .A2(G159), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1206), .B1(new_n1205), .B2(new_n1204), .C1(new_n1212), .C2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1197), .B1(new_n1217), .B2(new_n786), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1195), .A2(new_n780), .B1(new_n1196), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1128), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n756), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n748), .A2(new_n750), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n930), .B2(new_n576), .ZN(new_n1223));
  OAI21_X1  g1023(.A(G330), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT98), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n757), .A2(new_n732), .A3(G330), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n928), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1220), .B1(new_n1227), .B2(new_n894), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1163), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1228), .A2(new_n1229), .B1(new_n1125), .B2(new_n1159), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1167), .B1(new_n1132), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1195), .A2(new_n1231), .A3(KEYINPUT57), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n726), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1231), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1219), .B1(new_n1233), .B2(new_n1234), .ZN(G375));
  OAI211_X1 g1035(.A(new_n1166), .B(new_n1160), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT123), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT123), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n1166), .A4(new_n1160), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n1036), .A3(new_n1170), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT124), .Z(new_n1243));
  NAND2_X1  g1043(.A1(new_n970), .A2(new_n829), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n781), .B1(G68), .B2(new_n1151), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n810), .A2(G137), .B1(G58), .B2(new_n819), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n791), .A2(G132), .B1(new_n811), .B2(new_n1209), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n817), .A2(G50), .B1(new_n825), .B2(G159), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n250), .B1(new_n802), .B2(new_n433), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G128), .B2(new_n799), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n810), .A2(G283), .B1(G116), .B2(new_n811), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n250), .B(new_n1002), .C1(G107), .C2(new_n867), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1069), .B1(G294), .B2(new_n791), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n805), .A2(new_n220), .B1(new_n798), .B2(new_n641), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT125), .Z(new_n1257));
  OAI21_X1  g1057(.A(new_n1251), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1245), .B1(new_n1258), .B2(new_n786), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1164), .A2(new_n780), .B1(new_n1244), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1243), .A2(new_n1260), .ZN(G381));
  INV_X1    g1061(.A(G390), .ZN(new_n1262));
  INV_X1    g1062(.A(G384), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OR2_X1    g1064(.A1(G393), .A2(G396), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1264), .A2(G387), .A3(G378), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G375), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1243), .A3(new_n1267), .A4(new_n1260), .ZN(G407));
  OR3_X1    g1068(.A1(G375), .A2(G343), .A3(G378), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(G407), .A2(G213), .A3(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  INV_X1    g1071(.A(G213), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1272), .A2(G343), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(G2897), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT60), .B1(new_n1230), .B2(new_n1166), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT60), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n726), .B1(new_n1236), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1281), .B2(new_n1260), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1260), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1263), .B(new_n1283), .C1(new_n1277), .C2(new_n1280), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1275), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1279), .B1(new_n1241), .B2(new_n1276), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1263), .B1(new_n1286), .B2(new_n1283), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1281), .A2(G384), .A3(new_n1260), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(new_n1274), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1285), .A2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G378), .B(new_n1219), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n779), .B2(new_n1132), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1170), .A2(KEYINPUT120), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n727), .B1(new_n1294), .B2(new_n1133), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1168), .A2(new_n1132), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1293), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1195), .A2(new_n1231), .A3(new_n1036), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1219), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1273), .B1(new_n1291), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1271), .B1(new_n1290), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1291), .A2(new_n1300), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1273), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1306));
  AND4_X1   g1106(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1303), .B1(new_n1301), .B2(new_n1306), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1302), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G387), .A2(new_n1262), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(G393), .B(new_n844), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G390), .B(new_n1020), .C1(new_n1037), .C2(new_n1047), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(new_n1289), .A3(new_n1285), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1317), .A2(new_n1320), .A3(new_n1271), .A4(new_n1315), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1304), .A2(KEYINPUT63), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT126), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT126), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1301), .A2(new_n1324), .A3(KEYINPUT63), .A4(new_n1306), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  OAI22_X1  g1126(.A1(new_n1309), .A2(new_n1315), .B1(new_n1321), .B2(new_n1326), .ZN(G405));
  OAI22_X1  g1127(.A1(new_n1267), .A2(G378), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1291), .A2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1306), .A2(new_n1297), .A3(G375), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1328), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1330), .B1(new_n1328), .B2(new_n1331), .ZN(new_n1334));
  OAI22_X1  g1134(.A1(new_n1333), .A2(new_n1334), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1334), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1336), .A2(new_n1315), .A3(new_n1332), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(G402));
endmodule


