//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g035(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n459), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  XNOR2_X1  g048(.A(new_n462), .B(KEYINPUT68), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n466), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  MUX2_X1   g054(.A(G100), .B(G112), .S(G2105), .Z(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G136), .B1(G2104), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n477), .A2(new_n481), .ZN(G162));
  NAND2_X1  g057(.A1(KEYINPUT4), .A2(G138), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n460), .B2(new_n461), .ZN(new_n484));
  AND2_X1   g059(.A1(G102), .A2(G2104), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n466), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n460), .B2(new_n461), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n468), .A2(new_n469), .A3(G138), .A4(new_n466), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n486), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  AND3_X1   g071(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(G126), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n489), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G2105), .B1(new_n493), .B2(new_n492), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(new_n486), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G88), .B1(new_n518), .B2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n514), .A2(new_n519), .A3(KEYINPUT72), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G166));
  AND2_X1   g099(.A1(new_n516), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n528), .C1(new_n529), .C2(new_n517), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n510), .A2(new_n515), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n517), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI221_X1 g112(.A(KEYINPUT73), .B1(new_n517), .B2(new_n534), .C1(new_n532), .C2(new_n533), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n508), .B2(new_n509), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  AND2_X1   g122(.A1(G68), .A2(G543), .ZN(new_n548));
  OR3_X1    g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n549), .A2(G651), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n516), .A2(G81), .B1(new_n518), .B2(G43), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT76), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G188));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n517), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n515), .A2(new_n565), .A3(G53), .A4(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n516), .A2(G91), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n508), .B2(new_n509), .ZN(new_n570));
  AND2_X1   g145(.A1(G78), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  INV_X1    g150(.A(new_n509), .ZN(new_n576));
  OR3_X1    g151(.A1(new_n576), .A2(G74), .A3(new_n507), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n516), .A2(G87), .B1(G651), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n515), .A2(G49), .A3(G543), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n510), .A2(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G48), .B2(new_n518), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n510), .A2(G86), .A3(new_n515), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n510), .A2(new_n589), .A3(G86), .A4(new_n515), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n586), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n511), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n541), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(new_n595), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n516), .A2(G85), .B1(new_n518), .B2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  XOR2_X1   g175(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n532), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n601), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n604), .A2(G92), .A3(new_n510), .A4(new_n515), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n603), .A2(new_n605), .B1(G54), .B2(new_n518), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(new_n508), .B2(new_n509), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT81), .ZN(new_n610));
  OR3_X1    g185(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT82), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT82), .B1(new_n608), .B2(new_n610), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n611), .A2(G651), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n614), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g190(.A(new_n614), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  XOR2_X1   g192(.A(G299), .B(KEYINPUT83), .Z(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G860), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n614), .B1(G559), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT84), .ZN(G148));
  NOR2_X1   g198(.A1(new_n553), .A2(G868), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n614), .A2(G559), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n479), .A2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n475), .A2(G123), .ZN(new_n629));
  AND2_X1   g204(.A1(G111), .A2(G2105), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G99), .B2(new_n466), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n628), .B(new_n629), .C1(new_n467), .C2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT13), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(G156));
  INV_X1    g214(.A(G14), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2427), .ZN(new_n644));
  INV_X1    g219(.A(G2430), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n640), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n647), .B2(new_n653), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT85), .Z(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n660), .B1(new_n666), .B2(new_n657), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n658), .B2(new_n665), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n658), .A2(new_n661), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n664), .B1(new_n669), .B2(KEYINPUT17), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n663), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G2096), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n678), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  AOI211_X1 g257(.A(new_n680), .B(new_n682), .C1(new_n675), .C2(new_n679), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(G229));
  NOR2_X1   g264(.A1(G16), .A2(G23), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT86), .Z(new_n691));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n692));
  NAND2_X1  g267(.A1(G288), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n578), .A2(new_n581), .A3(KEYINPUT87), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  MUX2_X1   g274(.A(G6), .B(G305), .S(G16), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(G22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT88), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n696), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1971), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n699), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(G25), .A2(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n479), .A2(G131), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n475), .A2(G119), .ZN(new_n713));
  MUX2_X1   g288(.A(G95), .B(G107), .S(G2105), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G2104), .ZN(new_n715));
  AND3_X1   g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n711), .B1(new_n716), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G24), .B(G290), .S(G16), .Z(new_n720));
  INV_X1    g295(.A(G1986), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n709), .A2(new_n710), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT36), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT31), .B(G11), .Z(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n632), .B2(new_n726), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n696), .A2(G21), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G168), .B2(new_n696), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1966), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n696), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n696), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n729), .B(new_n732), .C1(G1961), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n726), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n726), .ZN(new_n738));
  INV_X1    g313(.A(G2078), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(G32), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n475), .A2(G129), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT93), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT26), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n467), .A2(G2105), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(G105), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G141), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n478), .A2(KEYINPUT92), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n479), .B2(G141), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n743), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n741), .B1(new_n753), .B2(new_n726), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  OAI211_X1 g330(.A(new_n736), .B(new_n740), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G35), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G162), .B2(G29), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT29), .Z(new_n759));
  INV_X1    g334(.A(G2090), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT95), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n756), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  MUX2_X1   g338(.A(G104), .B(G116), .S(G2105), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n475), .A2(G128), .B1(G2104), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n479), .A2(G140), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT89), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n726), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n554), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G16), .B2(G19), .ZN(new_n775));
  INV_X1    g350(.A(G1341), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  INV_X1    g354(.A(new_n614), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G4), .B2(G16), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n777), .B(new_n778), .C1(new_n779), .C2(new_n782), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n746), .A2(G103), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT25), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(KEYINPUT25), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n468), .A2(new_n469), .A3(G127), .ZN(new_n787));
  INV_X1    g362(.A(G115), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n467), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n785), .A2(new_n786), .B1(G2105), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G139), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n478), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT91), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G29), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G33), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT90), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G2072), .ZN(new_n798));
  OR2_X1    g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  NAND2_X1  g374(.A1(KEYINPUT24), .A2(G34), .ZN(new_n800));
  AOI21_X1  g375(.A(G29), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G160), .B2(G29), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G2084), .Z(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n782), .B2(new_n779), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n696), .A2(G20), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT23), .Z(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G299), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1956), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n734), .B2(G1961), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n754), .A2(new_n755), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n783), .A2(new_n798), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI211_X1 g387(.A(new_n773), .B(new_n812), .C1(new_n759), .C2(new_n760), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT95), .B1(new_n759), .B2(new_n760), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n724), .A2(new_n763), .A3(new_n813), .A4(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NAND2_X1  g391(.A1(new_n780), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n541), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n532), .A2(new_n821), .B1(new_n822), .B2(new_n517), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n551), .A2(KEYINPUT96), .A3(new_n552), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT96), .B1(new_n551), .B2(new_n552), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n553), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n824), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n551), .A2(KEYINPUT96), .A3(new_n552), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n818), .B(new_n833), .Z(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n621), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n824), .A2(new_n621), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n632), .B(G160), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G162), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n716), .A2(new_n636), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n479), .A2(G142), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n475), .A2(G130), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(KEYINPUT99), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(KEYINPUT99), .ZN(new_n850));
  OR3_X1    g425(.A1(new_n466), .A2(KEYINPUT98), .A3(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT98), .B1(new_n466), .B2(G118), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n846), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AND4_X1   g430(.A1(new_n636), .A2(new_n712), .A3(new_n713), .A4(new_n715), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n845), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n845), .B2(new_n856), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n844), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n767), .A2(new_n495), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n767), .A2(new_n495), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n753), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n862), .B(new_n863), .C1(new_n752), .C2(new_n743), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n793), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n793), .A2(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n865), .A2(new_n868), .A3(new_n866), .A4(new_n793), .ZN(new_n872));
  AOI211_X1 g447(.A(new_n859), .B(new_n861), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  AND4_X1   g448(.A1(KEYINPUT100), .A2(new_n871), .A3(new_n872), .A4(new_n860), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n843), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g452(.A(KEYINPUT101), .B(new_n843), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n873), .A2(new_n874), .ZN(new_n880));
  AOI21_X1  g455(.A(G37), .B1(new_n880), .B2(new_n842), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g458(.A1(new_n830), .A2(G868), .ZN(new_n884));
  XNOR2_X1  g459(.A(G166), .B(G305), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n695), .B(G290), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n885), .B(new_n886), .Z(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT42), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n833), .B(new_n625), .ZN(new_n890));
  AOI21_X1  g465(.A(G299), .B1(new_n613), .B2(new_n606), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n606), .A2(G299), .A3(new_n613), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n891), .B2(KEYINPUT102), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT103), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n896), .B2(KEYINPUT41), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  OAI211_X1 g476(.A(KEYINPUT104), .B(new_n901), .C1(new_n893), .C2(new_n895), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n780), .B2(G299), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n905));
  NAND4_X1  g480(.A1(new_n904), .A2(new_n892), .A3(new_n894), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n890), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n889), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n884), .B1(new_n910), .B2(G868), .ZN(G295));
  AOI21_X1  g486(.A(new_n884), .B1(new_n910), .B2(G868), .ZN(G331));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  AOI21_X1  g488(.A(G168), .B1(new_n539), .B2(new_n542), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n539), .A2(G168), .A3(new_n542), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n827), .A2(new_n832), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n827), .A2(new_n832), .B1(new_n915), .B2(new_n916), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n918), .A2(new_n896), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n916), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n833), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(KEYINPUT107), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n917), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n920), .B1(new_n926), .B2(new_n907), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT108), .B1(new_n927), .B2(new_n887), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n917), .B1(new_n919), .B2(KEYINPUT107), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n833), .A2(KEYINPUT107), .A3(new_n921), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n902), .A2(new_n906), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n904), .A2(new_n892), .A3(new_n894), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT104), .B1(new_n932), .B2(new_n901), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n929), .A2(new_n930), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n920), .ZN(new_n935));
  AND4_X1   g510(.A1(KEYINPUT108), .A2(new_n934), .A3(new_n887), .A4(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n913), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n927), .A2(new_n887), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n922), .A2(new_n917), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n932), .A2(new_n905), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n943), .A2(KEYINPUT41), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n918), .B2(new_n919), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n930), .B2(new_n929), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n947), .B2(new_n932), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n942), .B1(new_n948), .B2(new_n887), .ZN(new_n949));
  INV_X1    g524(.A(new_n887), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n896), .B1(new_n926), .B2(new_n946), .ZN(new_n951));
  OAI211_X1 g526(.A(KEYINPUT109), .B(new_n950), .C1(new_n951), .C2(new_n945), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n941), .B1(new_n953), .B2(new_n937), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n940), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n953), .B2(new_n937), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n934), .A2(new_n887), .A3(new_n935), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n927), .A2(KEYINPUT108), .A3(new_n887), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n952), .A4(new_n949), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n939), .A2(new_n941), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n955), .B1(new_n967), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n495), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(G160), .A2(G40), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G2067), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n767), .B(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n977), .B2(new_n753), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT46), .Z(new_n981));
  NOR2_X1   g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT47), .Z(new_n983));
  NOR3_X1   g558(.A1(new_n975), .A2(G1986), .A3(G290), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT48), .Z(new_n985));
  NAND2_X1  g560(.A1(new_n753), .A2(new_n979), .ZN(new_n986));
  OAI21_X1  g561(.A(G1996), .B1(new_n743), .B2(new_n752), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n977), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n716), .B(new_n718), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n985), .B1(new_n990), .B2(new_n975), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n716), .A2(new_n718), .ZN(new_n992));
  OAI22_X1  g567(.A1(new_n988), .A2(new_n992), .B1(G2067), .B2(new_n767), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n974), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n983), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n522), .A2(G8), .A3(new_n523), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT55), .Z(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n501), .B2(new_n486), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n973), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n496), .B2(new_n503), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT112), .B1(new_n1003), .B2(new_n1000), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n502), .B1(new_n501), .B2(new_n486), .ZN(new_n1005));
  AND4_X1   g580(.A1(new_n502), .A2(new_n486), .A3(new_n491), .A4(new_n494), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n969), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT50), .ZN(new_n1009));
  AOI211_X1 g584(.A(G2090), .B(new_n1002), .C1(new_n1004), .C2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n504), .B2(new_n969), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n973), .B1(new_n1011), .B2(KEYINPUT111), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT111), .B1(new_n970), .B2(new_n971), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1971), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(G8), .B(new_n998), .C1(new_n1010), .C2(new_n1015), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n693), .A2(G1976), .A3(new_n694), .ZN(new_n1017));
  INV_X1    g592(.A(G40), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n465), .A2(new_n472), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n999), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G8), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1021), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n693), .A2(G1976), .A3(new_n694), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n515), .A2(G48), .A3(G543), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1030), .B(new_n587), .C1(new_n1031), .C2(new_n541), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G1981), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(KEYINPUT113), .A3(G1981), .ZN(new_n1036));
  INV_X1    g611(.A(G1981), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n586), .A2(new_n591), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1029), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1036), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT113), .B1(new_n1032), .B2(G1981), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1029), .B(new_n1040), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1021), .B1(new_n1047), .B2(KEYINPUT49), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1028), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1016), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n998), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1007), .A2(KEYINPUT111), .A3(new_n971), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1014), .A2(new_n1052), .A3(new_n1019), .ZN(new_n1053));
  INV_X1    g628(.A(G1971), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(new_n760), .A3(new_n1019), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1055), .A2(KEYINPUT115), .A3(new_n1058), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(G8), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1050), .B1(new_n1051), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n972), .A2(new_n1019), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(KEYINPUT45), .B2(new_n1003), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n739), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT126), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1012), .A2(new_n739), .A3(new_n1014), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1001), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT127), .B(G1961), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1065), .A2(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(G301), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1074), .A2(G2084), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1067), .A2(G1966), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(G168), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT51), .ZN(new_n1082));
  AOI21_X1  g657(.A(G168), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  OAI211_X1 g659(.A(G8), .B(new_n1080), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1082), .A2(new_n1085), .A3(KEYINPUT62), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT62), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1064), .B(new_n1077), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1057), .A2(new_n1019), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1014), .A2(new_n1052), .A3(new_n1019), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n1092));
  OAI22_X1  g667(.A1(G1956), .A2(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(KEYINPUT118), .ZN(new_n1097));
  MUX2_X1   g672(.A(new_n1095), .B(new_n1097), .S(G299), .Z(new_n1098));
  NOR3_X1   g673(.A1(new_n1093), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1020), .A2(G2067), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1074), .B2(new_n779), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n780), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1098), .B(KEYINPUT120), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1099), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1101), .A2(KEYINPUT124), .A3(KEYINPUT60), .A4(new_n614), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1100), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1002), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT60), .B(new_n1109), .C1(new_n1110), .C2(G1348), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1108), .B1(new_n1111), .B2(new_n780), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n780), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(KEYINPUT125), .A3(new_n1115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT121), .B(G1996), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n973), .A2(new_n970), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT58), .B(G1341), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n1053), .A2(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n553), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1098), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT123), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT61), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n1098), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1099), .A2(KEYINPUT61), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1128), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1106), .B1(new_n1120), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT53), .B(new_n739), .C1(new_n970), .C2(new_n971), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1076), .B1(new_n1066), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(G171), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1143), .B2(new_n1077), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(G171), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1071), .A2(G301), .A3(new_n1076), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(KEYINPUT54), .A3(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1139), .A2(new_n1144), .A3(new_n1064), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1088), .B1(new_n1138), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1045), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1048), .B1(new_n1150), .B2(new_n1041), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT52), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1016), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1151), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n578), .A2(new_n581), .A3(new_n1025), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1038), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1157), .B1(new_n1023), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1062), .A2(G8), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT115), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1051), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G8), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1110), .A2(new_n760), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(new_n1055), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1156), .B1(new_n998), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(G168), .A2(G8), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1165), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT116), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT116), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1165), .A2(new_n1175), .A3(new_n1169), .A4(new_n1171), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1168), .A2(new_n998), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1178), .A2(new_n1169), .A3(KEYINPUT63), .A4(new_n1171), .ZN(new_n1179));
  AOI211_X1 g754(.A(KEYINPUT117), .B(new_n1162), .C1(new_n1177), .C2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT117), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1175), .B1(new_n1064), .B2(new_n1171), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1176), .A2(new_n1174), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1181), .B1(new_n1184), .B2(new_n1161), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1149), .A2(new_n1180), .A3(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(G290), .B(new_n721), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n975), .B1(new_n990), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n996), .B1(new_n1186), .B2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g764(.A(G319), .ZN(new_n1191));
  OR4_X1    g765(.A1(new_n1191), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1192), .B1(new_n879), .B2(new_n881), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n1193), .A2(new_n954), .A3(new_n940), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


