//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT83), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  OAI21_X1  g005(.A(G113), .B1(new_n191), .B2(KEYINPUT5), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT79), .ZN(new_n193));
  XNOR2_X1  g007(.A(G116), .B(G119), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n192), .A2(new_n193), .B1(new_n194), .B2(KEYINPUT5), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT5), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT79), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT2), .B(G113), .Z(new_n202));
  AOI22_X1  g016(.A1(new_n195), .A2(new_n201), .B1(new_n194), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G107), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n204), .A2(G107), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n203), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G110), .B(G122), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n220), .A2(new_n200), .B1(new_n202), .B2(new_n194), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT64), .B1(new_n223), .B2(G146), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G143), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G125), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n226), .A2(G143), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n228), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n234), .A2(KEYINPUT67), .A3(new_n239), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G125), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n238), .A2(KEYINPUT68), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n229), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n245), .A2(new_n246), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n237), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G224), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT7), .B1(new_n256), .B2(G953), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n216), .A2(new_n222), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT80), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n237), .A2(new_n254), .A3(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n245), .A2(KEYINPUT80), .A3(new_n253), .A4(new_n246), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n257), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n261), .A2(KEYINPUT81), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT81), .ZN(new_n265));
  INV_X1    g079(.A(new_n263), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n237), .A2(new_n254), .A3(new_n260), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n259), .B(KEYINPUT82), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n215), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n221), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n205), .A2(new_n208), .A3(new_n210), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(G101), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n274), .A2(new_n211), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n202), .A2(new_n194), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT2), .B(G113), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n190), .A2(G116), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n198), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n272), .A3(G101), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n217), .B(new_n271), .C1(new_n275), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n269), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n222), .B1(new_n215), .B2(new_n203), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n237), .A2(new_n254), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n257), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT81), .B1(new_n261), .B2(new_n263), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n266), .A2(new_n265), .A3(new_n267), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT82), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n189), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n271), .B1(new_n275), .B2(new_n282), .ZN(new_n293));
  INV_X1    g107(.A(new_n217), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT6), .A3(new_n283), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n256), .A2(G953), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n286), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT6), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n299), .A3(new_n294), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT78), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n296), .A2(new_n298), .A3(new_n303), .A4(new_n300), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n188), .B1(new_n292), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n288), .A2(new_n289), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n259), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n283), .A3(new_n269), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n302), .A2(new_n304), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n311), .A2(new_n189), .A3(new_n187), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G214), .B1(G237), .B2(G902), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT9), .B(G234), .ZN(new_n316));
  OAI21_X1  g130(.A(G221), .B1(new_n316), .B2(G902), .ZN(new_n317));
  INV_X1    g131(.A(G469), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n229), .A2(new_n232), .B1(new_n234), .B2(new_n230), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n281), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n275), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n238), .B1(new_n240), .B2(KEYINPUT1), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n322), .A2(new_n234), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n245), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n270), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT75), .B(KEYINPUT10), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT11), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G137), .ZN(new_n330));
  INV_X1    g144(.A(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT11), .A3(G134), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G131), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n336));
  INV_X1    g150(.A(G131), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n330), .A2(new_n332), .A3(new_n337), .A4(new_n333), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(KEYINPUT66), .A3(G131), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n245), .A2(new_n253), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT10), .A3(new_n270), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n321), .A2(new_n327), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G110), .B(G140), .ZN(new_n345));
  INV_X1    g159(.A(G953), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n346), .A2(G227), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n341), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n342), .A2(new_n270), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n215), .B1(new_n245), .B2(new_n323), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT12), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n243), .A2(new_n244), .B1(new_n252), .B2(new_n229), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n215), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n341), .B1(new_n325), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT77), .B1(new_n360), .B2(KEYINPUT12), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n351), .B(KEYINPUT12), .C1(new_n352), .C2(new_n353), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT76), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n365), .A3(KEYINPUT12), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n350), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n321), .A2(new_n327), .A3(new_n343), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n351), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n349), .B1(new_n370), .B2(new_n344), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n318), .B(new_n189), .C1(new_n368), .C2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n349), .A3(new_n344), .ZN(new_n373));
  INV_X1    g187(.A(new_n344), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(new_n362), .B2(new_n367), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n373), .B(G469), .C1(new_n375), .C2(new_n349), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n318), .A2(new_n189), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n372), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n314), .A2(new_n315), .A3(new_n317), .A4(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n381));
  NOR2_X1   g195(.A1(G475), .A2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n204), .ZN(new_n385));
  INV_X1    g199(.A(G140), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G125), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n246), .A2(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT84), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(G146), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n389), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n226), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G237), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n346), .A3(G214), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n223), .ZN(new_n399));
  NOR2_X1   g213(.A1(G237), .A2(G953), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(G143), .A3(G214), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n401), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT18), .A3(G131), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n396), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT16), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n386), .A3(G125), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n389), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n226), .ZN(new_n411));
  OAI211_X1 g225(.A(G146), .B(new_n409), .C1(new_n389), .C2(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND4_X1   g227(.A1(G143), .A2(new_n397), .A3(new_n346), .A4(G214), .ZN(new_n414));
  AOI21_X1  g228(.A(G143), .B1(new_n400), .B2(G214), .ZN(new_n415));
  OAI21_X1  g229(.A(G131), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT85), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n404), .A2(new_n418), .A3(G131), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n413), .B1(new_n420), .B2(KEYINPUT17), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT17), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n399), .A2(new_n337), .A3(new_n401), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n417), .A2(new_n419), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n407), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n417), .A2(new_n419), .A3(new_n423), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n390), .A2(KEYINPUT19), .A3(new_n392), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n389), .A2(KEYINPUT19), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n226), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n412), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n385), .B1(new_n430), .B2(new_n406), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n385), .A2(new_n425), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n431), .A2(new_n432), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n383), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n381), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n431), .A2(new_n432), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n421), .A2(new_n424), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n385), .A3(new_n406), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n431), .A2(new_n432), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n382), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(new_n436), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n437), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n425), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n385), .A2(KEYINPUT88), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n189), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G475), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n223), .A2(G128), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT13), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n247), .A2(new_n249), .A3(G143), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G134), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n329), .A3(new_n453), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n197), .A2(G122), .ZN(new_n460));
  INV_X1    g274(.A(G122), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G116), .ZN(new_n462));
  OR3_X1    g276(.A1(new_n460), .A2(new_n462), .A3(G107), .ZN(new_n463));
  OAI21_X1  g277(.A(G107), .B1(new_n460), .B2(new_n462), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT14), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n197), .A3(G122), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT14), .B1(new_n461), .B2(G116), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT89), .B(new_n468), .C1(new_n469), .C2(new_n462), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT89), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n197), .A2(G122), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n471), .B(new_n472), .C1(new_n460), .C2(KEYINPUT14), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n470), .A2(new_n473), .A3(new_n474), .A4(G107), .ZN(new_n475));
  INV_X1    g289(.A(new_n459), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n329), .B1(new_n456), .B2(new_n453), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n475), .B(new_n463), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n473), .A2(G107), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n474), .B1(new_n479), .B2(new_n470), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n466), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G217), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n316), .A2(new_n482), .A3(G953), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n483), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n466), .B(new_n485), .C1(new_n478), .C2(new_n480), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n189), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G478), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n484), .A2(KEYINPUT91), .A3(new_n189), .A4(new_n486), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n487), .A2(new_n495), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(G234), .A2(G237), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n501), .A2(G952), .A3(new_n346), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT21), .B(G898), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT93), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n501), .A2(G902), .A3(G953), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n446), .A2(new_n452), .A3(new_n500), .A4(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT94), .B1(new_n380), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT24), .B(G110), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT73), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n238), .A2(G119), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT68), .B(G128), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(G119), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(KEYINPUT23), .A3(G119), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT23), .B1(new_n238), .B2(G119), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(new_n513), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n512), .A2(new_n515), .B1(new_n519), .B2(G110), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n412), .A3(new_n395), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n512), .A2(new_n515), .B1(new_n519), .B2(G110), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n413), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT22), .B(G137), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n346), .A2(G221), .A3(G234), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT74), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n521), .A2(new_n523), .A3(new_n527), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n482), .B1(G234), .B2(new_n189), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(G902), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n532), .B2(G902), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n530), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n531), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n534), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT65), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n236), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n319), .A2(KEYINPUT65), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(new_n340), .A3(new_n339), .A4(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n547));
  INV_X1    g361(.A(new_n333), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n329), .A2(G137), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n342), .A2(new_n338), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n339), .A2(new_n340), .A3(new_n319), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n338), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n358), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT30), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n280), .ZN(new_n558));
  INV_X1    g372(.A(new_n280), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n358), .B2(new_n554), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT69), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n339), .A2(new_n340), .A3(new_n319), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n551), .A2(new_n562), .A3(new_n563), .A4(new_n559), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT26), .B(G101), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n400), .A2(G210), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n561), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT31), .B1(new_n558), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n559), .B1(new_n552), .B2(new_n556), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n561), .A2(new_n564), .A3(new_n570), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT31), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT28), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n553), .B2(new_n560), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n233), .A2(KEYINPUT65), .A3(new_n235), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT65), .B1(new_n233), .B2(new_n235), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n555), .B1(new_n582), .B2(new_n351), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n561), .B(new_n564), .C1(new_n583), .C2(new_n559), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n579), .B1(new_n584), .B2(KEYINPUT28), .ZN(new_n585));
  OAI22_X1  g399(.A1(new_n572), .A2(new_n576), .B1(new_n585), .B2(new_n570), .ZN(new_n586));
  NOR2_X1   g400(.A1(G472), .A2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT71), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n591), .B(KEYINPUT32), .C1(new_n586), .C2(new_n587), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT29), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n569), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n561), .A2(new_n564), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n551), .A2(new_n562), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n280), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT72), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n559), .B1(new_n551), .B2(new_n562), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT72), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n578), .B(new_n595), .C1(new_n603), .C2(new_n577), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n569), .B(new_n579), .C1(new_n584), .C2(KEYINPUT28), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n569), .B1(new_n573), .B2(new_n596), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n594), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n604), .B(new_n189), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G472), .ZN(new_n609));
  INV_X1    g423(.A(new_n587), .ZN(new_n610));
  INV_X1    g424(.A(new_n596), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n546), .A2(new_n551), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n280), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n577), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n569), .B1(new_n614), .B2(new_n579), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n558), .A2(KEYINPUT31), .A3(new_n571), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n575), .B1(new_n573), .B2(new_n574), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n610), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT32), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n542), .B1(new_n593), .B2(new_n621), .ZN(new_n622));
  AND4_X1   g436(.A1(new_n446), .A2(new_n452), .A3(new_n500), .A4(new_n508), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n379), .A2(new_n317), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT94), .ZN(new_n626));
  INV_X1    g440(.A(new_n315), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n306), .B2(new_n313), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n623), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n510), .A2(new_n622), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT95), .B(G101), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G3));
  INV_X1    g446(.A(new_n187), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n292), .B2(new_n305), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n507), .B(new_n627), .C1(new_n634), .C2(new_n313), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n489), .A2(new_n490), .A3(new_n496), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT98), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n489), .A2(new_n638), .A3(new_n490), .A4(new_n496), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n484), .A2(new_n640), .A3(new_n486), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n484), .A2(KEYINPUT96), .A3(new_n640), .A4(new_n486), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n485), .A2(KEYINPUT97), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n640), .B1(new_n481), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n481), .B2(new_n645), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n490), .A2(G902), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n637), .A2(new_n639), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n446), .B2(new_n452), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n635), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n542), .ZN(new_n653));
  INV_X1    g467(.A(G472), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n586), .B2(new_n189), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n619), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n625), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT34), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n437), .A2(new_n661), .A3(new_n444), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n437), .B2(new_n444), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n445), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n635), .A2(new_n665), .A3(new_n452), .A4(new_n499), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n657), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT35), .B(G107), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(new_n656), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n541), .B1(new_n538), .B2(new_n539), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT36), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n528), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n524), .B(new_n673), .Z(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(new_n535), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n510), .A2(new_n629), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  AOI21_X1  g494(.A(new_n676), .B1(new_n593), .B2(new_n621), .ZN(new_n681));
  INV_X1    g495(.A(new_n445), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n435), .A2(new_n381), .A3(new_n436), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT87), .B1(new_n443), .B2(KEYINPUT20), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT99), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n682), .B1(new_n685), .B2(new_n662), .ZN(new_n686));
  INV_X1    g500(.A(new_n502), .ZN(new_n687));
  INV_X1    g501(.A(new_n506), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n687), .B1(new_n688), .B2(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n452), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n686), .A2(new_n500), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n627), .B1(new_n634), .B2(new_n313), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n625), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n681), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  XNOR2_X1  g509(.A(new_n689), .B(KEYINPUT39), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n625), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT40), .Z(new_n698));
  NOR2_X1   g512(.A1(new_n573), .A2(new_n574), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT101), .B1(new_n603), .B2(new_n570), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n600), .B(KEYINPUT72), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n701), .B(new_n569), .C1(new_n702), .C2(new_n596), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n699), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n189), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI211_X1 g520(.A(KEYINPUT102), .B(new_n699), .C1(new_n700), .C2(new_n703), .ZN(new_n707));
  OAI21_X1  g521(.A(G472), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n593), .A2(new_n620), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n314), .B(new_n710), .Z(new_n711));
  AOI21_X1  g525(.A(new_n500), .B1(new_n446), .B2(new_n452), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n315), .A3(new_n676), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n698), .A2(new_n709), .A3(new_n711), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n651), .A2(new_n716), .A3(new_n689), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n446), .A2(new_n452), .ZN(new_n718));
  INV_X1    g532(.A(new_n650), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n689), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT103), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n681), .A2(new_n693), .A3(new_n717), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  OAI21_X1  g537(.A(new_n591), .B1(new_n619), .B2(KEYINPUT32), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n588), .A2(KEYINPUT71), .A3(new_n589), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n620), .A4(new_n609), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n189), .B1(new_n368), .B2(new_n371), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n317), .A3(new_n372), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n726), .A2(new_n653), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n652), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT41), .B(G113), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NOR2_X1   g548(.A1(new_n666), .A2(new_n731), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT104), .B(G116), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G18));
  INV_X1    g551(.A(new_n676), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n726), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n623), .A2(new_n692), .A3(new_n730), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n190), .ZN(G21));
  OAI21_X1  g556(.A(new_n578), .B1(new_n603), .B2(new_n577), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n569), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n610), .B1(new_n744), .B2(new_n618), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n655), .A3(new_n542), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n729), .A2(new_n507), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n692), .A4(new_n712), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  AND2_X1   g563(.A1(new_n692), .A2(new_n730), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n745), .A2(new_n655), .A3(new_n676), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n721), .A2(new_n750), .A3(new_n717), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n721), .A2(new_n717), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n306), .A2(new_n315), .A3(new_n313), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n624), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n726), .A3(new_n653), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n588), .A2(new_n589), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n542), .B1(new_n621), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n756), .A2(new_n624), .A3(new_n754), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n721), .A3(new_n717), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n665), .A2(new_n452), .A3(new_n499), .A4(new_n689), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT105), .B1(new_n758), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT105), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n622), .A2(new_n691), .A3(new_n768), .A4(new_n757), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  OAI21_X1  g585(.A(new_n373), .B1(new_n375), .B2(new_n349), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n318), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n377), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n777), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT106), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n778), .A2(new_n372), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n781), .A2(new_n317), .A3(new_n696), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n719), .A2(new_n446), .A3(new_n452), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT43), .Z(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n670), .A3(new_n738), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n756), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(KEYINPUT107), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(KEYINPUT107), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n782), .B(new_n787), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  XOR2_X1   g605(.A(KEYINPUT108), .B(G137), .Z(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(G39));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n781), .A2(KEYINPUT109), .A3(new_n317), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT109), .B1(new_n781), .B2(new_n317), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n794), .B(KEYINPUT47), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n797), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n794), .A2(KEYINPUT47), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n794), .A2(KEYINPUT47), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n799), .A2(new_n800), .A3(new_n795), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n726), .A2(new_n653), .A3(new_n756), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n755), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT111), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n807));
  INV_X1    g621(.A(new_n805), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n807), .B(new_n808), .C1(new_n798), .C2(new_n802), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n386), .ZN(G42));
  INV_X1    g625(.A(new_n709), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n756), .A2(new_n729), .A3(new_n542), .A4(new_n687), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n651), .ZN(new_n815));
  OAI211_X1 g629(.A(G952), .B(new_n346), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n784), .A2(new_n502), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n746), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n816), .B1(new_n821), .B2(new_n750), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n819), .A2(new_n729), .A3(new_n756), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT48), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n761), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n824), .B1(new_n823), .B2(new_n761), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n814), .A2(new_n718), .A3(new_n719), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n823), .B2(new_n751), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n711), .A2(new_n315), .A3(new_n729), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n821), .A2(KEYINPUT50), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT50), .B1(new_n821), .B2(new_n830), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n829), .B(KEYINPUT51), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n819), .A2(new_n820), .A3(new_n756), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n728), .A2(new_n372), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n317), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n835), .B1(new_n803), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n827), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n837), .B1(new_n803), .B2(KEYINPUT119), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n798), .A2(new_n802), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n840), .B1(new_n844), .B2(new_n835), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n839), .B1(new_n845), .B2(KEYINPUT51), .ZN(new_n846));
  XNOR2_X1  g660(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n692), .A2(new_n712), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n689), .B(KEYINPUT113), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT114), .B1(new_n738), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n676), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n624), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n709), .A2(new_n848), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n722), .A2(new_n694), .A3(new_n752), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n726), .A2(new_n625), .A3(new_n692), .A4(new_n738), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n651), .A2(new_n716), .A3(new_n689), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n716), .B1(new_n651), .B2(new_n689), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n859), .B1(new_n862), .B2(new_n691), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(KEYINPUT52), .A3(new_n752), .A4(new_n855), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n759), .A2(new_n763), .B1(new_n767), .B2(new_n769), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n510), .B(new_n629), .C1(new_n622), .C2(new_n677), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n628), .A2(new_n508), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n446), .A2(new_n452), .A3(new_n499), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT112), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n869), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT112), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n508), .A4(new_n628), .ZN(new_n873));
  INV_X1    g687(.A(new_n657), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n731), .B1(new_n666), .B2(new_n652), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n748), .B1(new_n739), .B2(new_n740), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n657), .A2(new_n868), .A3(new_n815), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n721), .A2(new_n717), .A3(new_n751), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n690), .A2(new_n499), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n726), .A2(new_n665), .A3(new_n738), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n757), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n866), .A2(new_n876), .A3(new_n880), .A4(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(KEYINPUT117), .B(new_n847), .C1(new_n865), .C2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n764), .A2(new_n770), .A3(new_n885), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n878), .A2(new_n879), .ZN(new_n889));
  INV_X1    g703(.A(new_n877), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n875), .A4(new_n867), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n858), .A2(new_n864), .A3(new_n893), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n856), .A2(new_n893), .A3(new_n857), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT53), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n887), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n858), .A2(new_n864), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT117), .B1(new_n899), .B2(new_n847), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n899), .A2(new_n847), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n903), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  OAI22_X1  g722(.A1(new_n846), .A2(new_n908), .B1(G952), .B2(G953), .ZN(new_n909));
  INV_X1    g723(.A(new_n711), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n653), .A2(new_n315), .A3(new_n317), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n783), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n914), .A3(new_n812), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n909), .A2(new_n915), .ZN(G75));
  NAND2_X1  g730(.A1(new_n296), .A2(new_n300), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n298), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n901), .A2(new_n189), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(G210), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n346), .A2(G952), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n923), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n921), .B2(new_n188), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(G51));
  XNOR2_X1  g742(.A(new_n901), .B(KEYINPUT54), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n377), .B(KEYINPUT57), .Z(new_n930));
  OAI22_X1  g744(.A1(new_n929), .A2(new_n930), .B1(new_n371), .B2(new_n368), .ZN(new_n931));
  OAI211_X1 g745(.A(G902), .B(new_n776), .C1(new_n897), .C2(new_n900), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT121), .Z(new_n933));
  AOI21_X1  g747(.A(new_n925), .B1(new_n931), .B2(new_n933), .ZN(G54));
  NAND3_X1  g748(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n441), .A2(new_n442), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n925), .ZN(G60));
  INV_X1    g753(.A(new_n925), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n648), .B(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT59), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n940), .B1(new_n929), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n908), .B2(new_n943), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n897), .B2(new_n900), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n532), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n674), .B(new_n950), .C1(new_n897), .C2(new_n900), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(KEYINPUT61), .A3(new_n940), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n951), .B2(new_n532), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n954), .A2(new_n940), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n951), .A2(new_n532), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT61), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT124), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  INV_X1    g776(.A(new_n959), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n954), .A2(new_n940), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  INV_X1    g780(.A(new_n956), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n951), .A2(new_n952), .A3(new_n532), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n965), .B(new_n966), .C1(new_n969), .C2(new_n955), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n961), .A2(new_n970), .ZN(G66));
  OAI21_X1  g785(.A(G953), .B1(new_n505), .B2(new_n256), .ZN(new_n972));
  INV_X1    g786(.A(new_n891), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(G953), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n917), .B1(G898), .B2(new_n346), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G69));
  NAND2_X1  g790(.A1(new_n427), .A2(new_n428), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n557), .B(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n714), .A2(new_n752), .A3(new_n863), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n697), .A2(new_n756), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n982), .B(new_n622), .C1(new_n651), .C2(new_n871), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n791), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n803), .A2(new_n805), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n807), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n803), .A2(KEYINPUT111), .A3(new_n805), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n978), .B1(new_n988), .B2(G953), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n863), .A2(new_n752), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n761), .A2(new_n848), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n782), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n791), .A2(new_n866), .A3(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n994), .B(new_n346), .C1(new_n806), .C2(new_n809), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n978), .B1(G900), .B2(G953), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n990), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n989), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n346), .B1(G227), .B2(G900), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n999), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n989), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(G72));
  NOR2_X1   g817(.A1(new_n573), .A2(new_n596), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT126), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n570), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n988), .A2(new_n973), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  AOI21_X1  g823(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n994), .B(new_n973), .C1(new_n806), .C2(new_n809), .ZN(new_n1011));
  AOI211_X1 g825(.A(new_n570), .B(new_n1005), .C1(new_n1011), .C2(new_n1009), .ZN(new_n1012));
  INV_X1    g826(.A(new_n606), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1009), .B1(new_n1013), .B2(new_n699), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT127), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n940), .B1(new_n907), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1010), .A2(new_n1012), .A3(new_n1016), .ZN(G57));
endmodule


