//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n461), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n461), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n472), .B2(G101), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  AOI211_X1 g049(.A(KEYINPUT69), .B(new_n474), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n466), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g053(.A(KEYINPUT70), .B(new_n466), .C1(new_n473), .C2(new_n475), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n465), .B1(new_n478), .B2(new_n479), .ZN(G160));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n461), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n461), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n483), .B2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n462), .A2(KEYINPUT71), .A3(new_n461), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT72), .A3(G136), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  INV_X1    g070(.A(G136), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n488), .B1(new_n494), .B2(new_n497), .ZN(G162));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n481), .C2(new_n482), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n461), .C1(new_n481), .C2(new_n482), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n462), .A2(new_n506), .A3(G138), .A4(new_n461), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(new_n509), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n512), .B1(new_n513), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n516), .A2(new_n518), .B1(new_n515), .B2(G543), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n522), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n509), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n521), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n528), .B(new_n531), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n525), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT76), .B(G52), .Z(new_n543));
  OAI22_X1  g118(.A1(new_n521), .A2(new_n542), .B1(new_n529), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n519), .A2(new_n520), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(KEYINPUT77), .A3(G651), .ZN(new_n553));
  INV_X1    g128(.A(new_n521), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G81), .B1(G43), .B2(new_n530), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g134(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n560));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n529), .B2(new_n564), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n529), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n547), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n565), .A2(new_n566), .B1(new_n569), .B2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n521), .A2(KEYINPUT79), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n523), .A2(new_n572), .A3(new_n509), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(G91), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n547), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G49), .B2(new_n530), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n571), .A2(G87), .A3(new_n573), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n519), .A2(G61), .A3(new_n520), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G48), .B2(new_n530), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n571), .A2(G86), .A3(new_n573), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n525), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(KEYINPUT80), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n554), .A2(G85), .B1(G47), .B2(new_n530), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n592), .A2(KEYINPUT81), .A3(new_n593), .A4(new_n594), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G290));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G301), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n571), .A2(G92), .A3(new_n573), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT82), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n571), .A2(new_n604), .A3(G92), .A4(new_n573), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n547), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n613), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n606), .B2(new_n607), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n609), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n601), .B1(new_n622), .B2(new_n600), .ZN(G284));
  AOI21_X1  g198(.A(new_n601), .B1(new_n622), .B2(new_n600), .ZN(G321));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT85), .B1(new_n625), .B2(G868), .ZN(new_n626));
  NOR2_X1   g201(.A1(G168), .A2(new_n600), .ZN(new_n627));
  MUX2_X1   g202(.A(new_n626), .B(KEYINPUT85), .S(new_n627), .Z(G297));
  MUX2_X1   g203(.A(new_n626), .B(KEYINPUT85), .S(new_n627), .Z(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n622), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n556), .A2(new_n600), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n620), .B(KEYINPUT84), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n633), .A2(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n634), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n472), .A2(new_n462), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n493), .A2(G135), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(KEYINPUT86), .ZN(new_n645));
  INV_X1    g220(.A(G111), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n644), .A2(KEYINPUT86), .B1(new_n646), .B2(G2105), .ZN(new_n647));
  AOI22_X1  g222(.A1(new_n484), .A2(G123), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n641), .A2(new_n642), .A3(new_n650), .ZN(G156));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n655), .B(new_n661), .Z(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT87), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n668), .B2(new_n670), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(new_n687), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT20), .Z(new_n691));
  AOI211_X1 g266(.A(new_n689), .B(new_n691), .C1(new_n684), .C2(new_n688), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  XOR2_X1   g268(.A(G1981), .B(G1986), .Z(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n693), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT95), .Z(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n701), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(G1971), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G23), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT94), .Z(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G288), .B2(new_n701), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n704), .A2(G1971), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n705), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G6), .B(G305), .S(G16), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT32), .B(G1981), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT93), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  OR3_X1    g292(.A1(new_n713), .A2(KEYINPUT92), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT92), .B1(new_n713), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n718), .A2(KEYINPUT34), .A3(new_n719), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G24), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n597), .A2(new_n598), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G16), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n726), .A2(G1986), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(G1986), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(KEYINPUT90), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(KEYINPUT90), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT91), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n493), .A2(G131), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n737));
  INV_X1    g312(.A(G107), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G2105), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n484), .B2(G119), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n732), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n727), .A2(new_n728), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n722), .A2(new_n723), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT96), .B(KEYINPUT36), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n747), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n722), .A2(new_n745), .A3(new_n723), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n633), .A2(G16), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n701), .A2(G4), .ZN(new_n754));
  AND3_X1   g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n753), .B1(new_n752), .B2(new_n754), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n701), .A2(G5), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G301), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g336(.A1(G115), .A2(G2104), .ZN(new_n762));
  INV_X1    g337(.A(G127), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n483), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n461), .B1(new_n764), .B2(KEYINPUT99), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(KEYINPUT99), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n493), .A2(G139), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  NAND3_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G33), .B(new_n770), .S(G29), .Z(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(G2072), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT101), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(KEYINPUT101), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n761), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n732), .A2(G35), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n732), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT29), .ZN(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT24), .B(G34), .ZN(new_n781));
  AOI22_X1  g356(.A1(G160), .A2(G29), .B1(new_n733), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G2084), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT106), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n701), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT107), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G2084), .B2(new_n782), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n775), .A2(new_n780), .A3(new_n784), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n729), .A2(G32), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n493), .A2(KEYINPUT102), .A3(G141), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT102), .ZN(new_n795));
  INV_X1    g370(.A(G141), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n492), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n472), .A2(G105), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT103), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n484), .A2(G129), .ZN(new_n801));
  NAND3_X1  g376(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT26), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n798), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n793), .B1(new_n807), .B2(new_n729), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT27), .B(G1996), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n733), .A2(G26), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT28), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n484), .A2(G128), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT97), .ZN(new_n814));
  OR2_X1    g389(.A1(G104), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT98), .Z(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n493), .A2(G140), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n812), .B1(new_n820), .B2(G29), .ZN(new_n821));
  INV_X1    g396(.A(G2067), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n810), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n649), .A2(new_n732), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT30), .B(G28), .ZN(new_n826));
  OR2_X1    g401(.A1(KEYINPUT31), .A2(G11), .ZN(new_n827));
  NAND2_X1  g402(.A1(KEYINPUT31), .A2(G11), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n826), .A2(new_n729), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n758), .A2(new_n759), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n733), .A2(G27), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G164), .B2(new_n733), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G2078), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(G2078), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n830), .A2(new_n831), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n771), .A2(KEYINPUT100), .A3(G2072), .ZN(new_n837));
  OAI21_X1  g412(.A(KEYINPUT100), .B1(new_n771), .B2(G2072), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G16), .A2(G19), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n557), .B2(G16), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(G1341), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n701), .A2(G21), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G168), .B2(new_n701), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT104), .B(G1966), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n824), .A2(new_n839), .A3(new_n842), .A4(new_n846), .ZN(new_n847));
  NOR4_X1   g422(.A1(new_n755), .A2(new_n756), .A3(new_n792), .A4(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n751), .A2(new_n848), .ZN(G311));
  AND3_X1   g424(.A1(new_n751), .A2(KEYINPUT108), .A3(new_n848), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT108), .B1(new_n751), .B2(new_n848), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(G150));
  AOI22_X1  g427(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n525), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  INV_X1    g430(.A(G55), .ZN(new_n856));
  OAI22_X1  g431(.A1(new_n521), .A2(new_n855), .B1(new_n856), .B2(new_n529), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G860), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT37), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n622), .A2(G559), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n858), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n556), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n556), .A2(new_n867), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(new_n864), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n866), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n862), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n859), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n873), .A2(new_n874), .A3(new_n862), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n861), .B1(new_n876), .B2(new_n877), .ZN(G145));
  XNOR2_X1  g453(.A(new_n649), .B(KEYINPUT110), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(G160), .ZN(new_n880));
  INV_X1    g455(.A(G162), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n505), .A2(new_n507), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n499), .A2(new_n502), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT111), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n770), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n806), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n807), .A2(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n820), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n820), .B1(new_n896), .B2(new_n891), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n461), .A2(G118), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n898), .A2(KEYINPUT112), .ZN(new_n899));
  OAI21_X1  g474(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n898), .B2(KEYINPUT112), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n899), .A2(new_n901), .B1(new_n484), .B2(G130), .ZN(new_n902));
  INV_X1    g477(.A(G142), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n492), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n638), .ZN(new_n905));
  INV_X1    g480(.A(new_n741), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n895), .A2(new_n897), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT113), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n907), .B1(new_n895), .B2(new_n897), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI211_X1 g488(.A(KEYINPUT113), .B(new_n907), .C1(new_n895), .C2(new_n897), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n882), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n882), .A2(new_n908), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(new_n911), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT114), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n882), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n911), .B1(new_n909), .B2(new_n908), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n914), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT114), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n882), .A2(new_n908), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n925), .B2(new_n912), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT115), .B(KEYINPUT40), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n920), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n920), .B2(new_n927), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(G395));
  NAND2_X1  g506(.A1(new_n725), .A2(G303), .ZN(new_n932));
  XNOR2_X1  g507(.A(G305), .B(G288), .ZN(new_n933));
  NAND2_X1  g508(.A1(G290), .A2(G166), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n622), .B(new_n630), .C1(new_n869), .C2(new_n870), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n871), .B1(new_n633), .B2(G559), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n614), .A2(new_n625), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n618), .A2(G299), .A3(new_n609), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT116), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(KEYINPUT116), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n939), .A2(new_n940), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n939), .A2(new_n940), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(KEYINPUT41), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n943), .A2(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n938), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n938), .B1(new_n952), .B2(new_n948), .ZN(new_n954));
  OAI21_X1  g529(.A(G868), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n867), .A2(new_n600), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(G295));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n956), .ZN(G331));
  INV_X1    g533(.A(new_n870), .ZN(new_n959));
  AOI21_X1  g534(.A(G301), .B1(new_n959), .B2(new_n868), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n869), .A2(G171), .A3(new_n870), .ZN(new_n961));
  OAI21_X1  g536(.A(G286), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(G171), .B1(new_n869), .B2(new_n870), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(G301), .A3(new_n868), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(G168), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n950), .B2(new_n951), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n962), .A2(new_n965), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n947), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n935), .A2(new_n936), .ZN(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n937), .B1(new_n967), .B2(new_n969), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT43), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n973), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n968), .A2(KEYINPUT41), .A3(new_n943), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n971), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n947), .B1(new_n968), .B2(KEYINPUT41), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n917), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n975), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n972), .B2(new_n973), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n975), .A2(new_n979), .A3(KEYINPUT43), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(G397));
  INV_X1    g562(.A(KEYINPUT121), .ZN(new_n988));
  INV_X1    g563(.A(G1971), .ZN(new_n989));
  INV_X1    g564(.A(new_n465), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n461), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT68), .B1(new_n461), .B2(G2104), .ZN(new_n992));
  OAI21_X1  g567(.A(G101), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT69), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n472), .A2(new_n467), .A3(G101), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT70), .B1(new_n996), .B2(new_n466), .ZN(new_n997));
  INV_X1    g572(.A(new_n479), .ZN(new_n998));
  OAI211_X1 g573(.A(G40), .B(new_n990), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G164), .B2(G1384), .ZN(new_n1001));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n989), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n885), .A2(new_n1007), .A3(new_n1002), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(G40), .A3(new_n779), .A4(G160), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(G166), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT55), .B(G8), .C1(new_n522), .C2(new_n526), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AND4_X1   g591(.A1(KEYINPUT118), .A2(new_n1011), .A3(G8), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1013), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT118), .B1(new_n1018), .B2(new_n1016), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n478), .A2(new_n479), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n885), .A2(new_n1002), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1020), .A2(new_n1022), .A3(G40), .A4(new_n990), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n581), .A2(new_n582), .A3(G1976), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1023), .A2(G8), .A3(new_n1024), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n587), .A2(new_n1030), .A3(new_n588), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n523), .A2(G86), .A3(new_n509), .ZN(new_n1033));
  INV_X1    g608(.A(new_n585), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n523), .B2(G61), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1032), .B(new_n1033), .C1(new_n1035), .C2(new_n525), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G1981), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(KEYINPUT119), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(G8), .A3(new_n1023), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1038), .B2(KEYINPUT119), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1026), .B(new_n1029), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1017), .A2(new_n1019), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1023), .A2(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G288), .A2(G1976), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1031), .B(KEYINPUT120), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n988), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1050), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1011), .A2(G8), .A3(new_n1016), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1018), .A2(KEYINPUT118), .A3(new_n1016), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1052), .B(KEYINPUT121), .C1(new_n1057), .C2(new_n1043), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1051), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1016), .B1(new_n1011), .B2(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1043), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n845), .B1(new_n999), .B2(new_n1004), .ZN(new_n1062));
  INV_X1    g637(.A(G2084), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1009), .A2(G40), .A3(new_n1063), .A4(G160), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1013), .B(G286), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1057), .A2(new_n1061), .A3(KEYINPUT63), .A4(new_n1065), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1011), .A2(G8), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1016), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1076), .B(KEYINPUT49), .C1(new_n1031), .C2(new_n1037), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1045), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1042), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1078), .A2(new_n1079), .B1(KEYINPUT52), .B2(new_n1025), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(new_n1080), .A3(new_n1029), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1071), .B1(new_n1072), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n999), .A2(G2078), .A3(new_n1004), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT124), .B1(new_n1084), .B2(KEYINPUT53), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT45), .B1(new_n885), .B2(new_n1002), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1000), .B(G1384), .C1(new_n883), .C2(new_n884), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G2078), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(G40), .A3(new_n1089), .A4(G160), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(G160), .A2(G40), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n759), .ZN(new_n1096));
  INV_X1    g671(.A(G40), .ZN(new_n1097));
  AOI211_X1 g672(.A(new_n1097), .B(new_n465), .C1(new_n478), .C2(new_n479), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1092), .A2(G2078), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1088), .A3(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1096), .A2(G301), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1083), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1003), .A2(new_n1099), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n999), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT45), .B1(new_n1021), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1105), .B2(new_n1021), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1104), .A2(new_n1107), .B1(new_n1095), .B2(new_n759), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1091), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G171), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1062), .A2(new_n1064), .A3(G168), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  AOI21_X1  g689(.A(G168), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1117), .A3(G8), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1102), .A2(new_n1112), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1057), .A2(KEYINPUT125), .A3(new_n1061), .ZN(new_n1120));
  OAI211_X1 g695(.A(G301), .B(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1123), .B2(G301), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1083), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1082), .A2(new_n1119), .A3(new_n1120), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1023), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1127), .A2(new_n822), .B1(new_n1095), .B2(new_n753), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1095), .A2(new_n789), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n570), .B2(new_n574), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1098), .A2(new_n1088), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1130), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1129), .A2(new_n620), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1134), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1128), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n616), .A2(new_n619), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1098), .A2(new_n822), .A3(new_n1022), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n753), .B1(new_n999), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1147), .A3(KEYINPUT60), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1143), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n620), .B1(new_n1149), .B2(new_n1148), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1151), .A2(new_n1152), .B1(KEYINPUT60), .B2(new_n1128), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1130), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1134), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT61), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1141), .A2(new_n1157), .A3(new_n1137), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT58), .B(G1341), .Z(new_n1162));
  AND2_X1   g737(.A1(new_n1023), .A2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n999), .A2(G1996), .A3(new_n1004), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n557), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1161), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n557), .B(new_n1166), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1156), .A2(new_n1158), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1142), .B1(new_n1153), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1059), .B(new_n1070), .C1(new_n1126), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1142), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1128), .A2(KEYINPUT60), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1150), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n620), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1176), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1175), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1057), .A2(KEYINPUT125), .A3(new_n1061), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT125), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1185), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1051), .A2(new_n1058), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1190), .A2(new_n1191), .A3(KEYINPUT126), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n1195));
  AOI211_X1 g770(.A(G301), .B(new_n1123), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1196), .B(new_n1189), .C1(new_n1195), .C2(new_n1194), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1174), .A2(new_n1192), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1107), .A2(new_n999), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n820), .B(new_n822), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n806), .B(G1996), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n906), .A2(new_n743), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n906), .A2(new_n743), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(G290), .A2(G1986), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AND2_X1   g783(.A1(G290), .A2(G1986), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1199), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1198), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1204), .B(KEYINPUT127), .ZN(new_n1212));
  AOI22_X1  g787(.A1(new_n1203), .A2(new_n1212), .B1(new_n822), .B2(new_n893), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1199), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1199), .B1(new_n1201), .B2(new_n806), .ZN(new_n1216));
  OR2_X1    g791(.A1(new_n1214), .A2(G1996), .ZN(new_n1217));
  AND2_X1   g792(.A1(new_n1217), .A2(KEYINPUT46), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1217), .A2(KEYINPUT46), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1216), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT47), .Z(new_n1221));
  NOR3_X1   g796(.A1(G290), .A2(new_n1214), .A3(G1986), .ZN(new_n1222));
  OR2_X1    g797(.A1(new_n1222), .A2(KEYINPUT48), .ZN(new_n1223));
  AOI22_X1  g798(.A1(new_n1206), .A2(new_n1199), .B1(KEYINPUT48), .B2(new_n1222), .ZN(new_n1224));
  AOI211_X1 g799(.A(new_n1215), .B(new_n1221), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1211), .A2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g801(.A(G319), .ZN(new_n1228));
  NOR4_X1   g802(.A1(G229), .A2(new_n1228), .A3(G401), .A4(G227), .ZN(new_n1229));
  NOR3_X1   g803(.A1(new_n916), .A2(KEYINPUT114), .A3(new_n919), .ZN(new_n1230));
  AOI21_X1  g804(.A(new_n924), .B1(new_n923), .B2(new_n926), .ZN(new_n1231));
  OAI21_X1  g805(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g806(.A1(new_n984), .A2(new_n985), .ZN(new_n1233));
  NOR2_X1   g807(.A1(new_n1232), .A2(new_n1233), .ZN(G308));
  OAI221_X1 g808(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .C1(new_n984), .C2(new_n985), .ZN(G225));
endmodule


