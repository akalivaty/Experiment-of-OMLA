//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT2), .B(G113), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT2), .A2(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT2), .A2(G113), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n194), .A2(new_n188), .A3(new_n190), .A4(new_n195), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n193), .A2(KEYINPUT66), .A3(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT66), .B1(new_n193), .B2(new_n196), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  AOI21_X1  g017(.A(G128), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(KEYINPUT1), .A3(G146), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT65), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n208), .B(new_n205), .C1(new_n209), .C2(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n201), .A2(new_n203), .A3(new_n212), .A4(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n215), .B2(G134), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(G134), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n215), .A2(G134), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT11), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(G134), .B2(new_n215), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n218), .A2(KEYINPUT11), .A3(G137), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n223), .B(new_n225), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n214), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n201), .A2(new_n203), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n209), .A2(KEYINPUT0), .A3(G128), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n220), .A2(KEYINPUT11), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n226), .A2(new_n215), .A3(G134), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n223), .B1(new_n241), .B2(new_n225), .ZN(new_n242));
  INV_X1    g056(.A(new_n229), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n199), .B1(new_n232), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n230), .B1(new_n211), .B2(new_n213), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n236), .A2(new_n237), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G131), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n249), .B2(new_n229), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n193), .A2(new_n196), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n193), .A2(KEYINPUT66), .A3(new_n196), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n246), .A2(new_n250), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT28), .B1(new_n245), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT67), .B1(new_n256), .B2(KEYINPUT28), .ZN(new_n258));
  INV_X1    g072(.A(new_n213), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n207), .B2(new_n210), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n244), .B(new_n199), .C1(new_n260), .C2(new_n230), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G237), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G210), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(G101), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n257), .A2(new_n258), .A3(new_n264), .A4(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n251), .B1(new_n246), .B2(new_n250), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n261), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT28), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n279), .A2(new_n258), .A3(new_n264), .A4(new_n270), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(new_n246), .B2(new_n250), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n244), .B(KEYINPUT30), .C1(new_n260), .C2(new_n230), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n251), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n261), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n271), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n280), .A2(new_n286), .A3(new_n287), .A4(new_n272), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n276), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT29), .B1(new_n285), .B2(new_n271), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n290), .B2(new_n280), .ZN(new_n291));
  OAI21_X1  g105(.A(G472), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G472), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n284), .A2(new_n261), .A3(new_n270), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT31), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n284), .A2(new_n296), .A3(new_n261), .A4(new_n270), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n262), .B1(new_n261), .B2(new_n263), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n270), .B1(new_n301), .B2(new_n279), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n293), .B(new_n275), .C1(new_n298), .C2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n279), .A2(new_n264), .A3(new_n258), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n295), .B(new_n297), .C1(new_n306), .C2(new_n270), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(KEYINPUT32), .A3(new_n293), .A4(new_n275), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n292), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G140), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n313), .A3(new_n200), .ZN(new_n314));
  INV_X1    g128(.A(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G119), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n315), .A2(G119), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n318), .A2(G110), .A3(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT24), .B(G110), .Z(new_n321));
  XNOR2_X1  g135(.A(G119), .B(G128), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n310), .A3(G125), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT69), .B1(new_n312), .B2(G140), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n312), .A2(G140), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT16), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n328), .A2(KEYINPUT16), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n200), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n314), .B(new_n324), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  AOI211_X1 g151(.A(G146), .B(new_n331), .C1(new_n329), .C2(KEYINPUT16), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n321), .A2(new_n322), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n318), .A2(new_n319), .ZN(new_n341));
  INV_X1    g155(.A(G110), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n346), .B(new_n347), .Z(new_n348));
  NAND3_X1  g162(.A1(new_n337), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n314), .B1(new_n320), .B2(new_n323), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT16), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n310), .A2(G125), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n311), .B1(new_n353), .B2(KEYINPUT69), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n354), .B2(new_n326), .ZN(new_n355));
  OAI21_X1  g169(.A(G146), .B1(new_n355), .B2(new_n331), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT70), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n351), .B1(new_n358), .B2(new_n334), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n350), .B1(new_n359), .B2(new_n344), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n349), .A2(new_n360), .A3(new_n275), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n349), .A2(new_n360), .A3(KEYINPUT25), .A4(new_n275), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G217), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(G234), .B2(new_n275), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT71), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n369));
  INV_X1    g183(.A(new_n367), .ZN(new_n370));
  AOI211_X1 g184(.A(new_n369), .B(new_n370), .C1(new_n363), .C2(new_n364), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n349), .A2(new_n360), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n367), .A2(G902), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n368), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n309), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT72), .ZN(new_n379));
  INV_X1    g193(.A(G221), .ZN(new_n380));
  XOR2_X1   g194(.A(KEYINPUT9), .B(G234), .Z(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(new_n275), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G107), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n387), .A2(KEYINPUT3), .A3(G104), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT3), .B1(new_n387), .B2(G104), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n384), .B(new_n386), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT73), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(G104), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n393), .B2(G101), .ZN(new_n394));
  AOI211_X1 g208(.A(KEYINPUT73), .B(new_n384), .C1(new_n386), .C2(new_n392), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n260), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G104), .B(G107), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT73), .B1(new_n398), .B2(new_n384), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n391), .A3(G101), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n213), .B(new_n205), .C1(G128), .C2(new_n209), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(new_n390), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n249), .A2(new_n229), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT76), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT12), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n211), .B2(new_n213), .ZN(new_n411));
  OAI211_X1 g225(.A(KEYINPUT74), .B(new_n390), .C1(new_n394), .C2(new_n395), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT74), .B1(new_n401), .B2(new_n390), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G101), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n419), .A3(G101), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n238), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n403), .A2(new_n410), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n405), .A2(KEYINPUT75), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT75), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n249), .A2(new_n424), .A3(new_n229), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n415), .A2(new_n421), .A3(new_n422), .A4(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G140), .ZN(new_n428));
  INV_X1    g242(.A(G227), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(G953), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n428), .B(new_n430), .Z(new_n431));
  INV_X1    g245(.A(KEYINPUT12), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n404), .A2(new_n432), .A3(new_n407), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n409), .A2(new_n427), .A3(new_n431), .A4(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT74), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n396), .A2(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(new_n410), .B(new_n260), .C1(new_n437), .C2(new_n412), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n421), .A2(new_n422), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n405), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n431), .B1(new_n440), .B2(new_n427), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n383), .B(new_n275), .C1(new_n435), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n431), .ZN(new_n445));
  AND4_X1   g259(.A1(new_n415), .A2(new_n421), .A3(new_n422), .A4(new_n426), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n421), .A2(new_n422), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n406), .B1(new_n447), .B2(new_n415), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n445), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(G902), .B1(new_n449), .B2(new_n434), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT78), .A3(new_n383), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n383), .A2(new_n275), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n427), .A2(new_n431), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n448), .B1(new_n454), .B2(KEYINPUT77), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT77), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n427), .A2(new_n456), .A3(new_n431), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n409), .A2(new_n427), .A3(new_n433), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n455), .A2(new_n457), .B1(new_n445), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n453), .B1(new_n459), .B2(G469), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n382), .B1(new_n452), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT79), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n188), .A2(KEYINPUT5), .ZN(new_n463));
  INV_X1    g277(.A(G113), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n196), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n437), .B2(new_n412), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n418), .A2(new_n420), .A3(new_n251), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n468), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n413), .B2(new_n414), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n418), .A2(new_n420), .A3(new_n251), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(KEYINPUT79), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G110), .B(G122), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n471), .A2(new_n475), .A3(KEYINPUT6), .A4(new_n477), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n469), .A2(new_n470), .A3(new_n477), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n260), .A2(new_n312), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n247), .A2(G125), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n266), .A2(G224), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G210), .B1(G237), .B2(G902), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT80), .Z(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(KEYINPUT7), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n487), .A2(new_n494), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n472), .A2(new_n396), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n472), .A2(new_n396), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n476), .B(KEYINPUT8), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n275), .B1(new_n501), .B2(new_n482), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n491), .A2(new_n493), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n493), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n482), .B1(new_n478), .B2(new_n479), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n489), .B1(new_n506), .B2(new_n481), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n507), .B2(new_n502), .ZN(new_n508));
  OAI21_X1  g322(.A(G214), .B1(G237), .B2(G902), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n461), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(KEYINPUT82), .A2(KEYINPUT18), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n265), .A2(new_n266), .A3(G214), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT81), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(G143), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT81), .B(G143), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n516), .B(new_n223), .C1(new_n514), .C2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n517), .A2(new_n514), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n223), .B1(new_n520), .B2(new_n516), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n513), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n512), .A3(new_n516), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n312), .A2(KEYINPUT69), .A3(G140), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n313), .A2(new_n325), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n311), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n314), .B1(new_n526), .B2(new_n200), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G113), .B(G122), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n385), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT83), .Z(new_n531));
  INV_X1    g345(.A(KEYINPUT84), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n517), .A2(new_n514), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n265), .A2(new_n266), .A3(G214), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(KEYINPUT81), .B2(new_n202), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT17), .B(G131), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n339), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n200), .B(new_n332), .C1(new_n526), .C2(new_n352), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n356), .A2(new_n532), .A3(new_n538), .A4(new_n536), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n516), .B1(new_n514), .B2(new_n517), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G131), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n518), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n528), .B(new_n531), .C1(new_n537), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT85), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n356), .A2(new_n538), .A3(new_n536), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n543), .A3(new_n539), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(KEYINPUT85), .A3(new_n528), .A4(new_n531), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n541), .A2(new_n518), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n329), .A2(KEYINPUT19), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n311), .A2(new_n313), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(KEYINPUT19), .B2(new_n555), .ZN(new_n556));
  OAI221_X1 g370(.A(new_n553), .B1(G146), .B2(new_n556), .C1(new_n335), .C2(new_n336), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n528), .ZN(new_n558));
  INV_X1    g372(.A(new_n530), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n562));
  NOR2_X1   g376(.A1(G475), .A2(G902), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n547), .A2(new_n551), .B1(new_n559), .B2(new_n558), .ZN(new_n565));
  INV_X1    g379(.A(new_n563), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT20), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n550), .A2(new_n528), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n559), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n552), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n275), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n564), .A2(new_n567), .B1(new_n571), .B2(G475), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT13), .B1(new_n202), .B2(G128), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n202), .A2(G128), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT87), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n315), .A2(G143), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n575), .A2(new_n576), .B1(KEYINPUT13), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT87), .B1(new_n573), .B2(new_n574), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n218), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g394(.A1(KEYINPUT86), .A2(G122), .ZN(new_n581));
  NAND2_X1  g395(.A1(KEYINPUT86), .A2(G122), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n189), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n189), .A2(G122), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n387), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n582), .ZN(new_n587));
  NOR2_X1   g401(.A1(KEYINPUT86), .A2(G122), .ZN(new_n588));
  OAI21_X1  g402(.A(G116), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(G107), .A3(new_n584), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n202), .A2(G128), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n315), .A2(G143), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n218), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT88), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT88), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n591), .A2(new_n592), .A3(new_n595), .A4(new_n218), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n586), .A2(new_n590), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT89), .B1(new_n580), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n586), .A2(new_n590), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n576), .B(new_n592), .C1(new_n577), .C2(KEYINPUT13), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n577), .A2(KEYINPUT13), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n579), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G134), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT89), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n594), .A2(new_n596), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n599), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n589), .A2(KEYINPUT14), .A3(G107), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n586), .A2(new_n590), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G134), .B1(new_n577), .B2(new_n574), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n593), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n589), .A2(KEYINPUT14), .A3(G107), .A4(new_n584), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT90), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n609), .A2(new_n611), .A3(KEYINPUT90), .A4(new_n612), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n607), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n381), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n619), .A2(new_n366), .A3(G953), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n607), .A2(new_n617), .A3(new_n620), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n275), .ZN(new_n625));
  INV_X1    g439(.A(G478), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(KEYINPUT15), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n625), .B(new_n627), .Z(new_n628));
  NAND2_X1  g442(.A1(G234), .A2(G237), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(G952), .A3(new_n266), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT91), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT21), .B(G898), .Z(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(G902), .A3(G953), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n572), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT92), .B1(new_n511), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n547), .A2(new_n551), .B1(new_n568), .B2(new_n559), .ZN(new_n637));
  OAI21_X1  g451(.A(G475), .B1(new_n637), .B2(G902), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n565), .A2(KEYINPUT20), .A3(new_n566), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n634), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n625), .B(new_n627), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT92), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n461), .A4(new_n510), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT72), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n377), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n379), .A2(new_n636), .A3(new_n646), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G101), .ZN(G3));
  NOR2_X1   g464(.A1(new_n442), .A2(new_n443), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT78), .B1(new_n450), .B2(new_n383), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n460), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n382), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n365), .A2(new_n367), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n369), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n365), .A2(KEYINPUT71), .A3(new_n367), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n374), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n504), .A2(new_n508), .A3(new_n634), .A4(new_n509), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n307), .A2(new_n275), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G472), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n303), .ZN(new_n663));
  NOR4_X1   g477(.A1(new_n655), .A2(new_n659), .A3(new_n660), .A4(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(G478), .B1(new_n624), .B2(new_n275), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT93), .B(KEYINPUT33), .Z(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n622), .B2(new_n623), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT94), .B1(new_n607), .B2(new_n617), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT33), .B1(new_n669), .B2(new_n621), .ZN(new_n670));
  AOI211_X1 g484(.A(KEYINPUT94), .B(new_n620), .C1(new_n607), .C2(new_n617), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT95), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n598), .A2(new_n606), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n615), .B2(new_n616), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n620), .B1(new_n674), .B2(KEYINPUT94), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n669), .A2(new_n621), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT95), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(KEYINPUT33), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n668), .B1(new_n672), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n626), .A2(G902), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n665), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT96), .B1(new_n681), .B2(new_n572), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT96), .ZN(new_n683));
  INV_X1    g497(.A(new_n680), .ZN(new_n684));
  AOI211_X1 g498(.A(new_n668), .B(new_n684), .C1(new_n672), .C2(new_n678), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n641), .B(new_n683), .C1(new_n685), .C2(new_n665), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n664), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT34), .B(G104), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G6));
  NAND2_X1  g504(.A1(new_n572), .A2(new_n643), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n664), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT35), .B(G107), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  NAND2_X1  g509(.A1(new_n337), .A2(new_n345), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n350), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n373), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n657), .A2(new_n658), .A3(new_n699), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n700), .A2(new_n303), .A3(new_n662), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n636), .A2(new_n646), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT37), .B(G110), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G12));
  NAND4_X1  g518(.A1(new_n461), .A2(new_n309), .A3(new_n510), .A4(new_n700), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n631), .B(KEYINPUT97), .Z(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(G900), .B2(new_n633), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n572), .A2(new_n643), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT98), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n655), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n309), .A2(new_n700), .ZN(new_n713));
  INV_X1    g527(.A(new_n709), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT98), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n713), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  XOR2_X1   g532(.A(new_n708), .B(KEYINPUT39), .Z(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n461), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT40), .Z(new_n722));
  AND2_X1   g536(.A1(new_n305), .A2(new_n308), .ZN(new_n723));
  INV_X1    g537(.A(new_n285), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n271), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n245), .A2(new_n256), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n275), .B1(new_n726), .B2(new_n270), .ZN(new_n727));
  OAI21_X1  g541(.A(G472), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n509), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n700), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n504), .A2(new_n508), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n572), .A2(new_n628), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n722), .A2(new_n729), .A3(new_n731), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G143), .ZN(G45));
  AND4_X1   g552(.A1(new_n461), .A2(new_n309), .A3(new_n510), .A4(new_n700), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n641), .B(new_n708), .C1(new_n685), .C2(new_n665), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G146), .ZN(G48));
  INV_X1    g557(.A(new_n450), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(G469), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n654), .B(new_n745), .C1(new_n651), .C2(new_n652), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT100), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n444), .A2(new_n451), .B1(G469), .B2(new_n744), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT100), .A3(new_n654), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n377), .A2(new_n660), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n687), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n751), .A3(new_n692), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  AND3_X1   g571(.A1(new_n748), .A2(new_n750), .A3(new_n510), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n309), .A2(new_n700), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n635), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G119), .ZN(G21));
  AOI21_X1  g576(.A(new_n270), .B1(new_n301), .B2(new_n257), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n298), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(G472), .A2(G902), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT101), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT102), .B(G472), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n661), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n764), .A2(KEYINPUT101), .A3(new_n765), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n659), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n641), .A2(new_n643), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n774), .A2(new_n642), .A3(new_n711), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n751), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G122), .ZN(G24));
  NAND4_X1  g591(.A1(new_n700), .A2(new_n770), .A3(new_n768), .A4(new_n771), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n740), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n758), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G125), .ZN(G27));
  INV_X1    g595(.A(KEYINPUT103), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n653), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n452), .A2(KEYINPUT103), .A3(new_n460), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n783), .A2(new_n654), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT104), .B1(new_n732), .B2(new_n509), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT104), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n787), .B(new_n730), .C1(new_n504), .C2(new_n508), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n785), .A2(new_n789), .A3(new_n378), .A4(new_n741), .ZN(new_n790));
  AND2_X1   g604(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n493), .B1(new_n491), .B2(new_n503), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n507), .A2(new_n505), .A3(new_n502), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n509), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n787), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n382), .B1(new_n653), .B2(new_n782), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n732), .A2(KEYINPUT104), .A3(new_n509), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n784), .ZN(new_n799));
  NOR2_X1   g613(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n791), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n799), .A2(new_n378), .A3(new_n741), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(new_n223), .ZN(G33));
  NAND4_X1  g618(.A1(new_n785), .A2(new_n789), .A3(new_n378), .A4(new_n714), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  NOR2_X1   g620(.A1(new_n681), .A2(new_n641), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT43), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n700), .A2(new_n663), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT44), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n796), .A2(new_n798), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(KEYINPUT44), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n459), .A2(G469), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT106), .ZN(new_n818));
  AND2_X1   g632(.A1(KEYINPUT45), .A2(G469), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n818), .B1(new_n817), .B2(new_n819), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n459), .A2(KEYINPUT45), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n453), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(KEYINPUT46), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n452), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT46), .B1(new_n823), .B2(new_n824), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n654), .A3(new_n720), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n812), .A2(KEYINPUT107), .A3(new_n813), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n816), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G137), .ZN(G39));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n828), .B2(new_n654), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n828), .A2(new_n834), .A3(new_n654), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n811), .A2(new_n309), .A3(new_n376), .A4(new_n740), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G140), .ZN(G42));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n748), .A2(new_n796), .A3(new_n750), .A4(new_n798), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n808), .A2(new_n706), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n841), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g662(.A(KEYINPUT116), .B(new_n846), .C1(new_n843), .C2(new_n844), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n378), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT48), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n729), .A2(new_n631), .A3(new_n659), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT117), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n687), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n850), .A2(new_n851), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n266), .A2(G952), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n706), .A2(new_n808), .A3(new_n751), .A4(new_n773), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n858), .B1(new_n859), .B2(new_n510), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n852), .A2(new_n856), .A3(new_n857), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n855), .A2(new_n572), .A3(new_n681), .ZN(new_n862));
  INV_X1    g676(.A(new_n778), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n848), .B2(new_n849), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n734), .A2(new_n509), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n867));
  XOR2_X1   g681(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n868));
  AOI21_X1  g682(.A(new_n867), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n862), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n749), .A2(new_n382), .ZN(new_n873));
  INV_X1    g687(.A(new_n837), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n835), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n846), .A2(new_n659), .A3(new_n772), .A4(new_n811), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n861), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n876), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT112), .B1(new_n836), .B2(new_n837), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n873), .B(KEYINPUT113), .Z(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n836), .A2(KEYINPUT112), .A3(new_n837), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n872), .B1(new_n884), .B2(new_n870), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n710), .A2(new_n716), .B1(new_n758), .B2(new_n779), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  INV_X1    g702(.A(new_n708), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n700), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n797), .A3(new_n784), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT110), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n729), .A2(new_n510), .A3(new_n735), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n890), .A2(new_n797), .A3(KEYINPUT110), .A4(new_n784), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n887), .A2(new_n888), .A3(new_n896), .A4(new_n742), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n715), .B1(new_n739), .B2(new_n714), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n705), .A2(KEYINPUT98), .A3(new_n709), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n780), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT109), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT109), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n717), .A2(new_n903), .A3(new_n780), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n902), .A2(new_n742), .A3(new_n896), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n898), .B1(new_n905), .B2(KEYINPUT52), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n753), .A2(new_n756), .A3(new_n776), .A4(new_n761), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n803), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n681), .A2(new_n572), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n664), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n649), .A2(new_n911), .ZN(new_n912));
  NOR4_X1   g726(.A1(new_n655), .A2(new_n643), .A3(new_n641), .A4(new_n889), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n713), .A3(new_n789), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n779), .A2(new_n785), .A3(new_n789), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n914), .A2(new_n805), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n702), .A2(new_n693), .A3(KEYINPUT108), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT108), .B1(new_n702), .B2(new_n693), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n912), .B(new_n916), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n906), .A2(new_n907), .A3(new_n909), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n702), .A2(new_n693), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT108), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n702), .A2(new_n693), .A3(KEYINPUT108), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n909), .A2(new_n926), .A3(new_n912), .A4(new_n916), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n896), .A2(new_n742), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT52), .B1(new_n928), .B2(new_n901), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n897), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT53), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n921), .A2(KEYINPUT54), .A3(new_n931), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n753), .A2(new_n756), .A3(new_n761), .A4(new_n776), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT111), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n933), .A2(new_n934), .A3(new_n792), .A4(new_n802), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT111), .B1(new_n803), .B2(new_n908), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT53), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n906), .A2(new_n937), .A3(new_n920), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT54), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n907), .B1(new_n927), .B2(new_n930), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n932), .A2(new_n941), .ZN(new_n942));
  OAI22_X1  g756(.A1(new_n886), .A2(new_n942), .B1(G952), .B2(G953), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n734), .A2(new_n729), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n376), .A2(new_n654), .A3(new_n509), .ZN(new_n945));
  INV_X1    g759(.A(new_n749), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(KEYINPUT49), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n946), .A2(KEYINPUT49), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n944), .A2(new_n947), .A3(new_n807), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n943), .A2(new_n949), .ZN(G75));
  NOR2_X1   g764(.A1(new_n484), .A2(new_n490), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n507), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT55), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n920), .A2(KEYINPUT53), .A3(new_n936), .A4(new_n935), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n742), .B1(new_n887), .B2(new_n903), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n717), .A2(new_n903), .A3(new_n780), .ZN(new_n956));
  INV_X1    g770(.A(new_n896), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n897), .B1(new_n958), .B2(new_n888), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n940), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(G902), .A3(new_n493), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT56), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n953), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT118), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI211_X1 g779(.A(KEYINPUT118), .B(new_n953), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n961), .A2(KEYINPUT119), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n275), .B1(new_n938), .B2(new_n940), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT119), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n970), .A3(new_n493), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n968), .A2(new_n962), .A3(new_n953), .A4(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n266), .A2(G952), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n967), .A2(new_n975), .ZN(G51));
  INV_X1    g790(.A(KEYINPUT120), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n275), .B(new_n823), .C1(new_n938), .C2(new_n940), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n453), .B(KEYINPUT57), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n939), .B1(new_n938), .B2(new_n940), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n449), .A2(new_n434), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n977), .B1(new_n984), .B2(new_n973), .ZN(new_n985));
  INV_X1    g799(.A(new_n983), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n960), .A2(KEYINPUT54), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n941), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(new_n979), .ZN(new_n989));
  OAI211_X1 g803(.A(KEYINPUT120), .B(new_n974), .C1(new_n989), .C2(new_n978), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n985), .A2(new_n990), .ZN(G54));
  AND3_X1   g805(.A1(new_n969), .A2(KEYINPUT58), .A3(G475), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n561), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n974), .ZN(new_n994));
  OR3_X1    g808(.A1(new_n992), .A2(KEYINPUT121), .A3(new_n561), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT121), .B1(new_n992), .B2(new_n561), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(G60));
  INV_X1    g811(.A(new_n679), .ZN(new_n998));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT59), .Z(new_n1000));
  NOR2_X1   g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n987), .B2(new_n941), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(KEYINPUT122), .B1(new_n1004), .B2(new_n974), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT122), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1003), .A2(new_n1006), .A3(new_n973), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1000), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n679), .B1(new_n942), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1005), .A2(new_n1007), .A3(new_n1009), .ZN(G63));
  NAND2_X1  g824(.A1(G217), .A2(G902), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT123), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT60), .Z(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n938), .B2(new_n940), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n973), .B1(new_n1014), .B2(new_n698), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n372), .B2(new_n1014), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT61), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(G66));
  AOI21_X1  g832(.A(new_n266), .B1(new_n632), .B2(G224), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n926), .A2(new_n933), .A3(new_n912), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1019), .B1(new_n1020), .B2(new_n266), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n506), .B(new_n481), .C1(G898), .C2(new_n266), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1021), .B(new_n1022), .Z(G69));
  NAND2_X1  g837(.A1(new_n379), .A2(new_n648), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n692), .A2(new_n910), .ZN(new_n1025));
  NOR4_X1   g839(.A1(new_n1024), .A2(new_n721), .A3(new_n811), .A4(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT125), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n832), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT126), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n955), .A2(new_n956), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n737), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT62), .Z(new_n1033));
  AND4_X1   g847(.A1(new_n266), .A2(new_n1030), .A3(new_n839), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n282), .A2(new_n283), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT124), .Z(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(new_n556), .Z(new_n1037));
  AND3_X1   g851(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n816), .A2(new_n831), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n378), .A2(new_n510), .A3(new_n735), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n829), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AND3_X1   g856(.A1(new_n792), .A2(new_n802), .A3(new_n805), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n839), .A2(new_n1031), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT127), .ZN(new_n1045));
  OR3_X1    g859(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1045), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1047));
  AOI21_X1  g861(.A(G953), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n429), .A2(G900), .A3(G953), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1037), .A2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g864(.A1(new_n1034), .A2(new_n1039), .B1(new_n1048), .B2(new_n1050), .ZN(G72));
  INV_X1    g865(.A(new_n725), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1020), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1030), .A2(new_n839), .A3(new_n1053), .A4(new_n1033), .ZN(new_n1054));
  NAND2_X1  g868(.A1(G472), .A2(G902), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT63), .Z(new_n1056));
  AOI21_X1  g870(.A(new_n1052), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n724), .A2(new_n271), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1046), .A2(new_n1053), .A3(new_n1047), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1058), .B1(new_n1059), .B2(new_n1056), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n286), .A2(new_n294), .ZN(new_n1061));
  NAND4_X1  g875(.A1(new_n921), .A2(new_n931), .A3(new_n1056), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1062), .A2(new_n974), .ZN(new_n1063));
  NOR3_X1   g877(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .ZN(G57));
endmodule


