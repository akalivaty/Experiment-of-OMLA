//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(KEYINPUT68), .ZN(new_n205));
  XOR2_X1   g004(.A(G127gat), .B(G134gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n203), .B(new_n202), .C1(new_n206), .C2(KEYINPUT68), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT69), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT28), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n216), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n217), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(G183gat), .B(G190gat), .Z(new_n228));
  AOI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(KEYINPUT24), .ZN(new_n229));
  INV_X1    g028(.A(new_n216), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n221), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(new_n216), .B2(KEYINPUT23), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n229), .A2(KEYINPUT66), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n234), .ZN(new_n237));
  XNOR2_X1  g036(.A(G183gat), .B(G190gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n226), .B1(new_n238), .B2(new_n225), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n231), .A2(G176gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G169gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(G169gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(new_n242), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n229), .A2(new_n232), .A3(new_n247), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n233), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n241), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n253), .B1(new_n241), .B2(new_n252), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n211), .B(new_n224), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n252), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n252), .A3(new_n253), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n223), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n210), .A2(KEYINPUT69), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G227gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT70), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n268), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT32), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT33), .B1(new_n267), .B2(new_n269), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n224), .B1(new_n254), .B2(new_n255), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n261), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n264), .A3(new_n256), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT34), .B1(new_n265), .B2(KEYINPUT71), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G15gat), .B(G43gat), .Z(new_n278));
  XNOR2_X1  g077(.A(G71gat), .B(G99gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n272), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n276), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n275), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT33), .ZN(new_n285));
  AOI211_X1 g084(.A(KEYINPUT70), .B(new_n264), .C1(new_n274), .C2(new_n256), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n268), .B1(new_n263), .B2(new_n265), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n288), .B2(new_n280), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n271), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n277), .B1(new_n272), .B2(new_n281), .ZN(new_n291));
  INV_X1    g090(.A(new_n271), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n284), .A3(new_n280), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT31), .B(G50gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G22gat), .ZN(new_n298));
  AND2_X1   g097(.A1(G228gat), .A2(G233gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(G155gat), .B(G162gat), .ZN(new_n300));
  XOR2_X1   g099(.A(G141gat), .B(G148gat), .Z(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  INV_X1    g101(.A(G162gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT2), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(new_n300), .A3(new_n304), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G197gat), .B(G204gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT22), .ZN(new_n313));
  INV_X1    g112(.A(G211gat), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT3), .B1(new_n321), .B2(new_n310), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n306), .A2(new_n308), .ZN(new_n323));
  OAI221_X1 g122(.A(new_n299), .B1(new_n311), .B2(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n311), .A2(new_n321), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n317), .A2(new_n326), .A3(new_n320), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n320), .A2(new_n326), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(new_n316), .A3(new_n312), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n332));
  OR3_X1    g131(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT29), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n331), .B2(KEYINPUT29), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n307), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n306), .A2(new_n308), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n325), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n298), .B(new_n324), .C1(new_n337), .C2(new_n299), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n297), .B1(new_n339), .B2(KEYINPUT79), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n324), .B1(new_n337), .B2(new_n299), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G22gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n342), .A2(KEYINPUT79), .A3(new_n338), .A4(new_n297), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n223), .B1(new_n252), .B2(new_n241), .ZN(new_n347));
  AND2_X1   g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(KEYINPUT29), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n260), .B2(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n352), .A2(new_n321), .ZN(new_n353));
  INV_X1    g152(.A(new_n321), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n260), .A2(new_n348), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n347), .A2(new_n351), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359));
  XOR2_X1   g158(.A(G8gat), .B(G36gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT74), .ZN(new_n361));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  NAND4_X1  g162(.A1(new_n353), .A2(new_n358), .A3(new_n359), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n353), .A2(new_n358), .A3(new_n363), .ZN(new_n365));
  INV_X1    g164(.A(new_n363), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n352), .A2(new_n321), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(new_n357), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT30), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n208), .A2(new_n209), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n336), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n323), .A2(new_n210), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT5), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(new_n370), .A3(new_n309), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n323), .A2(new_n210), .A3(KEYINPUT4), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n377), .A2(new_n379), .A3(new_n374), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT0), .ZN(new_n386));
  XNOR2_X1  g185(.A(G57gat), .B(G85gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n382), .A2(new_n384), .A3(KEYINPUT6), .A4(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n384), .A3(new_n389), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n382), .A2(new_n384), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n388), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT75), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n384), .A3(new_n398), .A4(new_n389), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n394), .A2(new_n396), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n364), .A2(new_n369), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n290), .A2(new_n294), .A3(new_n346), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT35), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n369), .A2(new_n364), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n396), .A2(new_n397), .A3(new_n393), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n392), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT83), .B(KEYINPUT35), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n408), .A2(new_n290), .A3(new_n294), .A4(new_n346), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n400), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n346), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT40), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT39), .ZN(new_n416));
  INV_X1    g215(.A(new_n374), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n388), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT39), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n417), .B2(new_n415), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n413), .B(new_n414), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n393), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n415), .A2(new_n417), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n388), .B(new_n418), .C1(new_n425), .C2(new_n421), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n414), .B1(new_n426), .B2(new_n413), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n369), .A2(new_n428), .A3(new_n364), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n429), .A2(new_n346), .ZN(new_n430));
  XOR2_X1   g229(.A(KEYINPUT82), .B(KEYINPUT37), .Z(new_n431));
  NAND3_X1  g230(.A1(new_n353), .A2(new_n358), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n366), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT37), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n353), .B2(new_n358), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT38), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n438));
  AND4_X1   g237(.A1(new_n437), .A2(new_n405), .A3(new_n438), .A4(new_n365), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n355), .A2(new_n354), .A3(new_n356), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n355), .A2(new_n442), .A3(new_n354), .A4(new_n356), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n352), .A2(new_n321), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n366), .A4(new_n432), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n436), .A2(new_n439), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n412), .B1(new_n430), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT36), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT72), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n451), .A2(KEYINPUT72), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT72), .A4(new_n451), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n410), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT15), .ZN(new_n460));
  NOR2_X1   g259(.A1(G43gat), .A2(G50gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G43gat), .A2(G50gat), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G36gat), .ZN(new_n465));
  AND2_X1   g264(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G29gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n472));
  INV_X1    g271(.A(G50gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G43gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(KEYINPUT85), .A2(G50gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n464), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n463), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT15), .B1(new_n481), .B2(new_n461), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n468), .B2(new_n470), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT17), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT17), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n471), .A2(new_n464), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n468), .A2(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n464), .ZN(new_n488));
  INV_X1    g287(.A(G1gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT16), .ZN(new_n490));
  INV_X1    g289(.A(G15gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G22gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n298), .A2(G15gat), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(G1gat), .B1(new_n492), .B2(new_n493), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n494), .A2(new_n495), .A3(G8gat), .ZN(new_n496));
  INV_X1    g295(.A(G8gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n298), .A2(G15gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n491), .A2(G22gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n489), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT86), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(G8gat), .B1(new_n494), .B2(new_n495), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n497), .A3(new_n501), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n484), .A2(new_n488), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n486), .B1(new_n487), .B2(new_n464), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n496), .A2(new_n502), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n508), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n508), .A2(new_n514), .A3(KEYINPUT18), .A4(new_n509), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n510), .B(new_n512), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n509), .B(KEYINPUT13), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G169gat), .B(G197gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n525), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n525), .B(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT12), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n522), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n521), .A4(new_n533), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(KEYINPUT87), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(KEYINPUT87), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n515), .A2(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n533), .B1(new_n539), .B2(new_n518), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n547));
  INV_X1    g346(.A(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G64gat), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G57gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n547), .B1(new_n552), .B2(KEYINPUT88), .ZN(new_n553));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n546), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(KEYINPUT89), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(new_n550), .A3(G57gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n560), .A3(new_n549), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n547), .B1(new_n544), .B2(new_n545), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n513), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n565));
  OAI211_X1 g364(.A(G231gat), .B(G233gat), .C1(new_n564), .C2(KEYINPUT21), .ZN(new_n566));
  INV_X1    g365(.A(G127gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n568), .B(new_n569), .C1(new_n557), .C2(new_n563), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n567), .B1(new_n566), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n565), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  INV_X1    g374(.A(new_n565), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT90), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G155gat), .ZN(new_n581));
  XOR2_X1   g380(.A(G183gat), .B(G211gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n574), .A2(new_n577), .A3(new_n583), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(KEYINPUT92), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT93), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT7), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(G85gat), .A3(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n596), .B2(new_n600), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n484), .A2(new_n606), .A3(new_n488), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT91), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n484), .A2(new_n606), .A3(KEYINPUT91), .A4(new_n488), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n588), .A2(KEYINPUT92), .ZN(new_n612));
  AND2_X1   g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n606), .B2(new_n510), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n591), .B1(new_n611), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n620));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n611), .A2(new_n591), .A3(new_n617), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  AOI211_X1 g424(.A(new_n590), .B(new_n616), .C1(new_n609), .C2(new_n610), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(new_n618), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT94), .B1(new_n587), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n585), .A2(new_n586), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI22_X1  g435(.A1(new_n557), .A2(new_n563), .B1(new_n603), .B2(new_n604), .ZN(new_n637));
  INV_X1    g436(.A(new_n546), .ZN(new_n638));
  INV_X1    g437(.A(new_n547), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n554), .B2(new_n555), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n549), .A2(new_n551), .A3(new_n555), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n561), .A2(new_n562), .ZN(new_n643));
  INV_X1    g442(.A(new_n604), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n602), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n637), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n564), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n636), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n637), .A2(new_n645), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n650), .B2(new_n636), .ZN(new_n651));
  XOR2_X1   g450(.A(G120gat), .B(G148gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT95), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n634), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n459), .A2(new_n543), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n459), .A2(KEYINPUT96), .A3(new_n543), .A4(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n411), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n404), .B1(new_n662), .B2(new_n663), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(new_n497), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  AOI21_X1  g470(.A(KEYINPUT97), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n671), .ZN(new_n675));
  AOI211_X1 g474(.A(new_n404), .B(new_n675), .C1(new_n662), .C2(new_n663), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n676), .A2(KEYINPUT97), .A3(KEYINPUT42), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n668), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(new_n673), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT42), .B1(new_n676), .B2(KEYINPUT97), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT98), .A4(new_n670), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(G1325gat));
  NOR2_X1   g481(.A1(new_n454), .A2(new_n455), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n491), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n456), .A2(new_n457), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n456), .A2(KEYINPUT99), .A3(new_n457), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n662), .B2(new_n663), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n684), .B1(new_n691), .B2(new_n491), .ZN(G1326gat));
  INV_X1    g491(.A(new_n346), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n664), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  NAND2_X1  g495(.A1(new_n459), .A2(new_n543), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n632), .A2(new_n658), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n628), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n469), .A3(new_n665), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n459), .B2(new_n628), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n450), .A3(new_n688), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n403), .A2(KEYINPUT101), .A3(new_n409), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT101), .B1(new_n403), .B2(new_n409), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n630), .A2(KEYINPUT44), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n705), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n538), .A2(new_n540), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n714));
  AOI211_X1 g513(.A(KEYINPUT87), .B(new_n533), .C1(new_n539), .C2(new_n518), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT100), .B1(new_n537), .B2(new_n541), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n698), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n703), .B1(new_n712), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n711), .ZN(new_n723));
  INV_X1    g522(.A(new_n707), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n708), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n723), .B1(new_n725), .B2(new_n706), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT102), .B(new_n720), .C1(new_n726), .C2(new_n705), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n722), .A2(new_n665), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n702), .B1(new_n728), .B2(new_n469), .ZN(G1328gat));
  INV_X1    g528(.A(new_n404), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n700), .A2(new_n465), .A3(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT46), .Z(new_n732));
  AND3_X1   g531(.A1(new_n722), .A2(new_n730), .A3(new_n727), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n465), .ZN(G1329gat));
  NAND2_X1  g533(.A1(new_n683), .A2(new_n475), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n697), .A2(new_n699), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n722), .A2(new_n727), .A3(new_n689), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n689), .B(new_n720), .C1(new_n726), .C2(new_n705), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G43gat), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n740), .A2(KEYINPUT103), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT103), .B1(new_n740), .B2(new_n743), .ZN(new_n745));
  OAI22_X1  g544(.A1(new_n738), .A2(KEYINPUT47), .B1(new_n744), .B2(new_n745), .ZN(G1330gat));
  AND2_X1   g545(.A1(new_n474), .A2(new_n476), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n346), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n700), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n722), .A2(new_n727), .A3(new_n693), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(KEYINPUT48), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n693), .B(new_n720), .C1(new_n726), .C2(new_n705), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(new_n748), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n758), .B(new_n754), .C1(new_n755), .C2(new_n748), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n753), .A2(KEYINPUT48), .B1(new_n757), .B2(new_n759), .ZN(G1331gat));
  NAND2_X1  g559(.A1(new_n718), .A2(new_n658), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n634), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n710), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n665), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n730), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT49), .B(G64gat), .Z(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(G1333gat));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n689), .ZN(new_n770));
  INV_X1    g569(.A(new_n683), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(G71gat), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n770), .A2(G71gat), .B1(new_n763), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n763), .A2(new_n693), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g576(.A1(new_n712), .A2(new_n632), .A3(new_n761), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n665), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G85gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n537), .A2(new_n541), .A3(KEYINPUT100), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n783), .A2(new_n632), .A3(new_n630), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n710), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n710), .B2(new_n784), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n665), .A2(new_n598), .A3(new_n658), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n780), .B1(new_n789), .B2(new_n790), .ZN(G1336gat));
  INV_X1    g590(.A(new_n784), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n725), .B2(new_n706), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n785), .A2(KEYINPUT106), .A3(KEYINPUT51), .ZN(new_n796));
  INV_X1    g595(.A(new_n658), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n404), .A2(G92gat), .A3(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n761), .A2(new_n632), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n730), .B(new_n800), .C1(new_n726), .C2(new_n705), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  INV_X1    g603(.A(new_n798), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n789), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n803), .B1(new_n802), .B2(new_n806), .ZN(G1337gat));
  NAND2_X1  g606(.A1(new_n778), .A2(new_n689), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G99gat), .ZN(new_n809));
  OR3_X1    g608(.A1(new_n771), .A2(G99gat), .A3(new_n797), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n789), .B2(new_n810), .ZN(G1338gat));
  OAI21_X1  g610(.A(new_n800), .B1(new_n726), .B2(new_n705), .ZN(new_n812));
  OAI21_X1  g611(.A(G106gat), .B1(new_n812), .B2(new_n346), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n346), .A2(G106gat), .A3(new_n797), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n787), .B2(new_n788), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT107), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n795), .A2(new_n796), .A3(new_n814), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT107), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n813), .A2(new_n815), .A3(new_n822), .A4(new_n816), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n821), .A3(new_n823), .ZN(G1339gat));
  NOR3_X1   g623(.A1(new_n634), .A2(new_n658), .A3(new_n783), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n647), .A2(new_n648), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n635), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n647), .A2(new_n648), .A3(new_n636), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n655), .B1(new_n649), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n657), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT55), .B1(new_n829), .B2(new_n831), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT108), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n519), .A2(new_n520), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n509), .B1(new_n508), .B2(new_n514), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n531), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n536), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n624), .B2(new_n627), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n829), .A2(new_n831), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT108), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n843), .A2(new_n844), .A3(new_n657), .A4(new_n832), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n835), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT109), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT109), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n835), .A2(new_n840), .A3(new_n845), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n658), .A2(new_n536), .A3(new_n838), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n835), .A2(new_n845), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n783), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n630), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n835), .A2(new_n845), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n855), .B(new_n851), .C1(new_n718), .C2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n850), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n825), .B1(new_n860), .B2(new_n587), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n411), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n771), .A2(new_n693), .A3(new_n730), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865), .B2(new_n783), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n861), .A2(new_n693), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT111), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n861), .B2(new_n693), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n730), .A2(new_n411), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n683), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n543), .A2(G113gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n866), .B1(new_n875), .B2(new_n876), .ZN(G1340gat));
  AOI21_X1  g676(.A(G120gat), .B1(new_n865), .B2(new_n658), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n658), .A2(G120gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n875), .B2(new_n879), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n874), .B2(new_n587), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n567), .A3(new_n632), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1342gat));
  NAND3_X1  g682(.A1(new_n871), .A2(new_n628), .A3(new_n873), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G134gat), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n630), .A2(G134gat), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT56), .B1(new_n864), .B2(new_n886), .ZN(new_n887));
  OR3_X1    g686(.A1(new_n864), .A2(KEYINPUT56), .A3(new_n886), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT112), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n885), .A2(KEYINPUT112), .A3(new_n887), .A4(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1343gat));
  NOR3_X1   g692(.A1(new_n689), .A2(new_n346), .A3(new_n730), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n542), .A2(G141gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n862), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT116), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n894), .A2(new_n862), .A3(new_n898), .A4(new_n895), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT58), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n687), .A2(new_n688), .A3(new_n872), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n825), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n851), .B1(new_n718), .B2(new_n857), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n628), .B1(new_n905), .B2(KEYINPUT110), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n906), .A2(new_n858), .B1(new_n847), .B2(new_n849), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n904), .B1(new_n907), .B2(new_n632), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT57), .B1(new_n908), .B2(new_n693), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n346), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n832), .A2(new_n657), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n834), .A2(KEYINPUT113), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT113), .ZN(new_n914));
  AOI211_X1 g713(.A(new_n914), .B(KEYINPUT55), .C1(new_n829), .C2(new_n831), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n851), .B1(new_n916), .B2(new_n542), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n630), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n632), .B1(new_n850), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n911), .B1(new_n919), .B2(new_n825), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT114), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g721(.A(KEYINPUT114), .B(new_n911), .C1(new_n919), .C2(new_n825), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n903), .B1(new_n909), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G141gat), .B1(new_n925), .B2(new_n542), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n900), .A2(new_n901), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n901), .B1(new_n900), .B2(new_n926), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n857), .B1(new_n782), .B2(new_n781), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT110), .B1(new_n929), .B2(new_n852), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n630), .A3(new_n858), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n632), .B1(new_n931), .B2(new_n850), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n693), .B1(new_n932), .B2(new_n825), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n924), .B1(new_n933), .B2(new_n910), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT115), .B1(new_n934), .B2(new_n902), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n936), .B(new_n903), .C1(new_n909), .C2(new_n924), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n783), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n894), .A2(new_n862), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n938), .A2(G141gat), .B1(new_n939), .B2(new_n895), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT58), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n927), .A2(new_n928), .B1(new_n940), .B2(new_n941), .ZN(G1344gat));
  NAND3_X1  g741(.A1(new_n935), .A2(new_n658), .A3(new_n937), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT118), .ZN(new_n944));
  INV_X1    g743(.A(G148gat), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(KEYINPUT59), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n943), .B2(new_n946), .ZN(new_n948));
  INV_X1    g747(.A(new_n911), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT119), .B1(new_n861), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n951), .B(new_n911), .C1(new_n932), .C2(new_n825), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n840), .A2(new_n912), .A3(new_n843), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n632), .B1(new_n918), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n542), .B2(new_n659), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n910), .B1(new_n955), .B2(new_n346), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n950), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n658), .A3(new_n903), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G148gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT120), .B1(new_n959), .B2(KEYINPUT59), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT59), .ZN(new_n962));
  AOI211_X1 g761(.A(new_n961), .B(new_n962), .C1(new_n958), .C2(G148gat), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n947), .A2(new_n948), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n939), .A2(new_n945), .A3(new_n658), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1345gat));
  NAND3_X1  g765(.A1(new_n939), .A2(KEYINPUT121), .A3(new_n632), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n967), .A2(new_n302), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n939), .A2(new_n632), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(KEYINPUT121), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n632), .A2(G155gat), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT122), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n935), .A2(new_n937), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n970), .A2(new_n973), .ZN(G1346gat));
  NAND3_X1  g773(.A1(new_n939), .A2(new_n303), .A3(new_n628), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n935), .A2(new_n628), .A3(new_n937), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n303), .ZN(G1347gat));
  NOR2_X1   g776(.A1(new_n665), .A2(new_n404), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n683), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n871), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(G169gat), .B1(new_n980), .B2(new_n542), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n867), .A2(new_n979), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n982), .A2(new_n248), .A3(new_n783), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1348gat));
  OAI21_X1  g783(.A(G176gat), .B1(new_n980), .B2(new_n797), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n982), .A2(new_n220), .A3(new_n658), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1349gat));
  NAND4_X1  g786(.A1(new_n868), .A2(new_n632), .A3(new_n870), .A4(new_n979), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G183gat), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n982), .A2(new_n212), .A3(new_n632), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(KEYINPUT123), .A3(new_n990), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g791(.A1(new_n982), .A2(new_n213), .A3(new_n628), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n871), .A2(new_n628), .A3(new_n979), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n994), .A2(new_n995), .A3(G190gat), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(new_n994), .B2(G190gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(G1351gat));
  NAND3_X1  g797(.A1(new_n687), .A2(new_n688), .A3(new_n978), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n933), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g799(.A(KEYINPUT124), .B(G197gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1000), .A2(new_n783), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n687), .A2(KEYINPUT125), .A3(new_n688), .A4(new_n978), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(new_n957), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1007), .A2(new_n542), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1002), .B1(new_n1008), .B2(new_n1001), .ZN(G1352gat));
  NAND3_X1  g808(.A1(new_n1006), .A2(new_n957), .A3(new_n658), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n1012));
  NAND4_X1  g811(.A1(new_n1006), .A2(new_n957), .A3(new_n1012), .A4(new_n658), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1011), .A2(G204gat), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n797), .A2(G204gat), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g815(.A(new_n1016), .B(KEYINPUT62), .Z(new_n1017));
  NAND2_X1  g816(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1014), .A2(new_n1017), .A3(KEYINPUT127), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1020), .A2(new_n1021), .ZN(G1353gat));
  NAND3_X1  g821(.A1(new_n1000), .A2(new_n314), .A3(new_n632), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1006), .A2(new_n957), .A3(new_n632), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1024), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(KEYINPUT63), .B1(new_n1024), .B2(G211gat), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(G1354gat));
  OAI21_X1  g826(.A(G218gat), .B1(new_n1007), .B2(new_n630), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1000), .A2(new_n315), .A3(new_n628), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1028), .A2(new_n1029), .ZN(G1355gat));
endmodule


