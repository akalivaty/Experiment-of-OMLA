//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  OAI21_X1  g000(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n202));
  NOR4_X1   g001(.A1(KEYINPUT85), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT85), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(KEYINPUT86), .B(new_n202), .C1(new_n203), .C2(new_n207), .ZN(new_n211));
  NAND2_X1  g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n202), .ZN(new_n218));
  NOR3_X1   g017(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n219));
  OAI22_X1  g018(.A1(new_n214), .A2(KEYINPUT15), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n212), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n216), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT89), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(G1gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT16), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT87), .B1(new_n226), .B2(G1gat), .ZN(new_n231));
  OAI21_X1  g030(.A(G8gat), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n226), .A2(G1gat), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n233), .A2(KEYINPUT87), .A3(new_n234), .A4(new_n229), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n224), .A2(new_n225), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n222), .B1(new_n213), .B2(new_n216), .ZN(new_n238));
  INV_X1    g037(.A(new_n236), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT89), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT90), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(new_n238), .B2(new_n239), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n221), .B1(new_n208), .B2(new_n209), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n215), .B1(new_n243), .B2(new_n211), .ZN(new_n244));
  NOR4_X1   g043(.A1(new_n244), .A2(new_n236), .A3(KEYINPUT90), .A4(new_n222), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n237), .B(new_n240), .C1(new_n242), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT88), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT13), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n224), .A2(new_n236), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n239), .B1(new_n238), .B2(KEYINPUT17), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n244), .A2(new_n253), .A3(new_n222), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n248), .B(new_n251), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT18), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n238), .A2(KEYINPUT17), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n253), .B1(new_n244), .B2(new_n222), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n239), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(KEYINPUT18), .A3(new_n248), .A4(new_n251), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n250), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G113gat), .B(G141gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G169gat), .B(G197gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n246), .A2(new_n249), .B1(new_n255), .B2(new_n256), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(new_n261), .A3(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G57gat), .B(G64gat), .Z(new_n275));
  INV_X1    g074(.A(KEYINPUT9), .ZN(new_n276));
  INV_X1    g075(.A(G71gat), .ZN(new_n277));
  INV_X1    g076(.A(G78gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G71gat), .B(G78gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n275), .A2(new_n281), .A3(new_n279), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT21), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n239), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT21), .ZN(new_n289));
  INV_X1    g088(.A(G231gat), .ZN(new_n290));
  INV_X1    g089(.A(G233gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n285), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n285), .B2(new_n289), .ZN(new_n296));
  OAI21_X1  g095(.A(G127gat), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n296), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n294), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n288), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n300), .A3(new_n288), .ZN(new_n303));
  XNOR2_X1  g102(.A(G183gat), .B(G211gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT91), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n306));
  INV_X1    g105(.A(G155gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n305), .B(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n302), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n302), .B2(new_n303), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(G232gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT41), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n313), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G99gat), .B(G106gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G85gat), .A2(G92gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT92), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT7), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT7), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT92), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(KEYINPUT92), .A3(new_n325), .ZN(new_n328));
  NAND2_X1  g127(.A1(G99gat), .A2(G106gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT8), .ZN(new_n330));
  OR2_X1    g129(.A1(G85gat), .A2(G92gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n320), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT93), .ZN(new_n334));
  NOR2_X1   g133(.A1(G85gat), .A2(G92gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n323), .A2(KEYINPUT7), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(new_n321), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n319), .A4(new_n330), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n333), .A2(new_n334), .A3(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n327), .A2(new_n332), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(KEYINPUT93), .A3(new_n319), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n258), .A2(new_n259), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G190gat), .B(G218gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT94), .ZN(new_n348));
  OAI22_X1  g147(.A1(new_n347), .A2(KEYINPUT94), .B1(new_n315), .B2(new_n314), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n224), .B2(new_n343), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n345), .B2(new_n350), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n318), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n345), .A2(new_n350), .ZN(new_n355));
  INV_X1    g154(.A(new_n348), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n317), .A3(new_n351), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G120gat), .B(G148gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G176gat), .B(G204gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n285), .A3(new_n342), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n333), .A2(new_n283), .A3(new_n284), .A4(new_n339), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n343), .A2(KEYINPUT10), .A3(new_n286), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G230gat), .A2(G233gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n365), .ZN(new_n371));
  INV_X1    g170(.A(new_n369), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n362), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n368), .B2(KEYINPUT95), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT95), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n366), .A2(new_n376), .A3(new_n367), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n362), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n374), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n312), .A2(new_n359), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT34), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(G183gat), .A2(G190gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT66), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT25), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT23), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n390), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT23), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(G169gat), .B2(G176gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n388), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n387), .A2(KEYINPUT64), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT64), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n400), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n386), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT65), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(KEYINPUT65), .A3(new_n386), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n393), .A2(new_n389), .A3(new_n396), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT25), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n398), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT26), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n389), .B1(new_n392), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT68), .ZN(new_n414));
  INV_X1    g213(.A(new_n392), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(KEYINPUT26), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n392), .A2(KEYINPUT68), .A3(new_n412), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n419));
  AND2_X1   g218(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT27), .B(G183gat), .ZN(new_n421));
  INV_X1    g220(.A(G190gat), .ZN(new_n422));
  AOI211_X1 g221(.A(new_n419), .B(new_n420), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n419), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n385), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n418), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT70), .B1(new_n411), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G127gat), .B(G134gat), .ZN(new_n428));
  INV_X1    g227(.A(G113gat), .ZN(new_n429));
  INV_X1    g228(.A(G120gat), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT1), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G113gat), .A2(G120gat), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n428), .A2(KEYINPUT69), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G127gat), .B(G134gat), .Z(new_n434));
  INV_X1    g233(.A(KEYINPUT69), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n434), .A2(new_n435), .A3(new_n432), .A4(new_n431), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OR3_X1    g238(.A1(new_n418), .A2(new_n423), .A3(new_n425), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT25), .B1(new_n442), .B2(new_n406), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n440), .B(new_n441), .C1(new_n443), .C2(new_n398), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n409), .A2(new_n410), .ZN(new_n446));
  INV_X1    g245(.A(new_n398), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n426), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n439), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G227gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(new_n291), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n383), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  AOI211_X1 g254(.A(KEYINPUT34), .B(new_n453), .C1(new_n445), .C2(new_n450), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n445), .A2(new_n453), .A3(new_n450), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  XNOR2_X1  g258(.A(G15gat), .B(G43gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(G71gat), .B(G99gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n458), .B(KEYINPUT32), .C1(new_n459), .C2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n458), .B2(KEYINPUT32), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n458), .A2(new_n459), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(KEYINPUT71), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT71), .B1(new_n464), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n457), .B(new_n463), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n464), .A2(new_n465), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n464), .A2(KEYINPUT71), .A3(new_n465), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(KEYINPUT73), .A3(new_n457), .A4(new_n463), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n477));
  INV_X1    g276(.A(new_n457), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n470), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(G141gat), .B(G148gat), .Z(new_n484));
  INV_X1    g283(.A(G162gat), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT2), .B1(new_n307), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G155gat), .B(G162gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n488), .A3(new_n486), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(G197gat), .A2(G204gat), .ZN(new_n493));
  AND2_X1   g292(.A1(G197gat), .A2(G204gat), .ZN(new_n494));
  AND2_X1   g293(.A1(G211gat), .A2(G218gat), .ZN(new_n495));
  OAI22_X1  g294(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(KEYINPUT22), .ZN(new_n496));
  XNOR2_X1  g295(.A(G211gat), .B(G218gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT29), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n492), .B1(new_n499), .B2(KEYINPUT3), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n490), .A2(new_n501), .A3(new_n491), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n498), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n483), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT78), .B1(G228gat), .B2(G233gat), .ZN(new_n507));
  INV_X1    g306(.A(G22gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT77), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n506), .A2(new_n509), .ZN(new_n511));
  XNOR2_X1  g310(.A(G78gat), .B(G106gat), .ZN(new_n512));
  OR3_X1    g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n511), .B2(new_n510), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT31), .B(G50gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n515), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G226gat), .A2(G233gat), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(KEYINPUT74), .Z(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n448), .B2(KEYINPUT29), .ZN(new_n521));
  INV_X1    g320(.A(new_n520), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n411), .B2(new_n426), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n498), .ZN(new_n525));
  XNOR2_X1  g324(.A(G8gat), .B(G36gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G64gat), .B(G92gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  XOR2_X1   g327(.A(new_n496), .B(new_n497), .Z(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n529), .A3(new_n523), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT30), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(KEYINPUT30), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n525), .A2(new_n530), .ZN(new_n534));
  INV_X1    g333(.A(new_n528), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT75), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT75), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n538), .A3(new_n535), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n532), .A2(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n439), .B(new_n492), .ZN(new_n541));
  NAND2_X1  g340(.A1(G225gat), .A2(G233gat), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT5), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n492), .A2(KEYINPUT3), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(new_n449), .A3(new_n502), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT76), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n544), .A2(new_n449), .A3(KEYINPUT76), .A4(new_n502), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n490), .A2(new_n491), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n439), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT4), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n542), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n543), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n549), .A2(new_n552), .A3(KEYINPUT5), .A4(new_n542), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G1gat), .B(G29gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT0), .ZN(new_n559));
  XNOR2_X1  g358(.A(G57gat), .B(G85gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n563));
  INV_X1    g362(.A(new_n561), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n555), .A2(new_n564), .A3(new_n556), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n555), .A2(new_n564), .A3(new_n556), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n564), .B1(new_n555), .B2(new_n556), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n568), .B2(KEYINPUT6), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n540), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT83), .B(KEYINPUT35), .Z(new_n572));
  NOR4_X1   g371(.A1(new_n480), .A2(new_n518), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n468), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(new_n518), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n477), .A2(KEYINPUT72), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n475), .A2(new_n578), .A3(new_n463), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n579), .A3(new_n478), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT35), .B1(new_n581), .B2(new_n571), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT79), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n553), .B2(new_n554), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n553), .A2(new_n584), .A3(new_n554), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(new_n541), .B2(new_n542), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT80), .B(KEYINPUT39), .ZN(new_n591));
  AOI211_X1 g390(.A(KEYINPUT79), .B(new_n542), .C1(new_n549), .C2(new_n552), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n593), .A3(new_n561), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT40), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n590), .A2(new_n593), .A3(KEYINPUT40), .A4(new_n561), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n596), .A2(new_n565), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n540), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n518), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n534), .A2(KEYINPUT37), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(KEYINPUT82), .A3(new_n535), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT82), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n525), .B2(new_n530), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n605), .B2(new_n528), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n525), .A2(new_n604), .A3(new_n530), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT38), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n566), .A2(new_n569), .A3(new_n531), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n605), .A2(new_n528), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(KEYINPUT81), .A3(new_n612), .A4(new_n607), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n607), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT81), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n609), .A2(new_n610), .A3(new_n613), .A4(new_n616), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n600), .A2(new_n617), .B1(new_n518), .B2(new_n571), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT36), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n580), .B2(new_n468), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n470), .A2(new_n476), .A3(new_n479), .A4(new_n619), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  AOI211_X1 g423(.A(new_n274), .B(new_n382), .C1(new_n583), .C2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n570), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g427(.A1(new_n625), .A2(new_n599), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT96), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n234), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT42), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT97), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n629), .A2(new_n234), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n629), .A2(KEYINPUT42), .A3(new_n631), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(G1325gat));
  AOI21_X1  g435(.A(new_n457), .B1(new_n477), .B2(KEYINPUT72), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n575), .B1(new_n637), .B2(new_n579), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n621), .B1(new_n638), .B2(new_n619), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n625), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n480), .A2(G15gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n640), .A2(G15gat), .B1(new_n625), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT98), .Z(G1326gat));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n518), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT43), .B(G22gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  AOI21_X1  g445(.A(new_n359), .B1(new_n583), .B2(new_n624), .ZN(new_n647));
  INV_X1    g446(.A(new_n381), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n274), .A2(new_n312), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G29gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n626), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT45), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT35), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n576), .A2(new_n580), .ZN(new_n655));
  INV_X1    g454(.A(new_n571), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND4_X1   g456(.A1(new_n609), .A2(new_n610), .A3(new_n613), .A4(new_n616), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n515), .B(new_n516), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n596), .A2(new_n565), .A3(new_n597), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n660), .B2(new_n540), .ZN(new_n661));
  OAI22_X1  g460(.A1(new_n658), .A2(new_n661), .B1(new_n659), .B2(new_n656), .ZN(new_n662));
  OAI22_X1  g461(.A1(new_n657), .A2(new_n573), .B1(new_n662), .B2(new_n639), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n354), .A2(KEYINPUT99), .A3(new_n358), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT99), .B1(new_n354), .B2(new_n358), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n647), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n649), .ZN(new_n673));
  OAI21_X1  g472(.A(G29gat), .B1(new_n673), .B2(new_n570), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n653), .A2(new_n674), .ZN(G1328gat));
  NAND3_X1  g474(.A1(new_n650), .A2(new_n206), .A3(new_n599), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT46), .Z(new_n677));
  OAI21_X1  g476(.A(G36gat), .B1(new_n673), .B2(new_n540), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1329gat));
  INV_X1    g478(.A(new_n480), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n650), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n639), .A2(G43gat), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n681), .A2(G43gat), .B1(new_n673), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g483(.A(new_n359), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n671), .B1(new_n663), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n669), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n583), .B2(new_n624), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n518), .B(new_n649), .C1(new_n686), .C2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n672), .A2(KEYINPUT101), .A3(new_n518), .A4(new_n649), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(G50gat), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n659), .A2(G50gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT100), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n650), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT48), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n689), .A2(G50gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n696), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT48), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(G50gat), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n689), .B2(new_n690), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n697), .B1(new_n707), .B2(new_n692), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT48), .B1(new_n700), .B2(new_n696), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT102), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(new_n710), .ZN(G1331gat));
  INV_X1    g510(.A(new_n312), .ZN(new_n712));
  NOR4_X1   g511(.A1(new_n273), .A2(new_n712), .A3(new_n685), .A4(new_n381), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n663), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n626), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g516(.A1(new_n714), .A2(KEYINPUT103), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(KEYINPUT103), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n599), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT49), .B(G64gat), .Z(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(G1333gat));
  NOR2_X1   g523(.A1(new_n623), .A2(new_n277), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n718), .A2(new_n719), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(KEYINPUT104), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n277), .B1(new_n714), .B2(new_n480), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(KEYINPUT104), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n728), .B1(new_n727), .B2(new_n730), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n720), .A2(new_n518), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT105), .B(G78gat), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1335gat));
  NOR2_X1   g535(.A1(new_n273), .A2(new_n312), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n647), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT107), .B(KEYINPUT51), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741));
  AOI22_X1  g540(.A1(new_n647), .A2(new_n737), .B1(new_n741), .B2(KEYINPUT51), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  OR4_X1    g542(.A1(G85gat), .A2(new_n743), .A3(new_n570), .A4(new_n381), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n273), .A2(new_n312), .A3(new_n381), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n672), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n626), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G85gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n744), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n672), .A2(new_n599), .A3(new_n745), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(KEYINPUT52), .A3(G92gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n540), .A2(G92gat), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n648), .B(new_n755), .C1(new_n740), .C2(new_n742), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n754), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n753), .A2(KEYINPUT109), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n753), .A2(KEYINPUT109), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n756), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n764), .B2(new_n757), .ZN(G1337gat));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n639), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G99gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n680), .A2(new_n648), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n768), .A2(G99gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n743), .B2(new_n769), .ZN(G1338gat));
  INV_X1    g569(.A(G106gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n518), .A2(new_n771), .ZN(new_n772));
  OR3_X1    g571(.A1(new_n743), .A2(new_n381), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n746), .B2(new_n518), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n743), .A2(new_n381), .A3(new_n772), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT53), .B1(new_n778), .B2(new_n774), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1339gat));
  NOR2_X1   g579(.A1(new_n246), .A2(new_n249), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n248), .B1(new_n260), .B2(new_n251), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n267), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n648), .A2(new_n272), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n268), .B1(new_n271), .B2(new_n261), .ZN(new_n785));
  AND4_X1   g584(.A1(new_n261), .A2(new_n250), .A3(new_n257), .A4(new_n268), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n366), .A2(new_n372), .A3(new_n367), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT111), .A4(new_n372), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n375), .B2(new_n377), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  AOI211_X1 g593(.A(KEYINPUT54), .B(new_n372), .C1(new_n366), .C2(new_n367), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n362), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n368), .A2(new_n792), .A3(new_n369), .ZN(new_n797));
  INV_X1    g596(.A(new_n362), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(KEYINPUT112), .A3(new_n798), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n791), .A2(new_n793), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n785), .A2(new_n786), .B1(new_n800), .B2(KEYINPUT55), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n378), .A2(new_n380), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n796), .A2(new_n799), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n378), .A2(KEYINPUT54), .A3(new_n791), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n784), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n668), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n800), .A2(KEYINPUT55), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n272), .A2(new_n783), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n667), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n312), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n382), .A2(new_n273), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT110), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n626), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(new_n818), .A3(new_n581), .ZN(new_n819));
  INV_X1    g618(.A(new_n802), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n800), .B2(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n273), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n667), .B1(new_n823), .B2(new_n784), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT99), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n359), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n812), .A2(new_n664), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n822), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n712), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n815), .B(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n570), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT113), .B1(new_n833), .B2(new_n655), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n540), .B1(new_n819), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n273), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n830), .A2(new_n832), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NOR4_X1   g638(.A1(new_n839), .A2(new_n570), .A3(new_n518), .A4(new_n599), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n680), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(new_n429), .A3(new_n274), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n837), .A2(new_n842), .ZN(G1340gat));
  AOI21_X1  g642(.A(G120gat), .B1(new_n836), .B2(new_n648), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n768), .A2(new_n430), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n840), .B2(new_n845), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n841), .B2(new_n712), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n312), .A2(new_n299), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n835), .B2(new_n848), .ZN(G1342gat));
  OAI21_X1  g648(.A(G134gat), .B1(new_n841), .B2(new_n359), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT114), .Z(new_n851));
  NOR2_X1   g650(.A1(new_n359), .A2(G134gat), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n836), .A2(KEYINPUT56), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT56), .B1(new_n836), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(G1343gat));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n621), .B(new_n518), .C1(new_n638), .C2(new_n619), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n817), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n833), .A2(new_n623), .A3(KEYINPUT118), .A4(new_n518), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n274), .A2(G141gat), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n540), .A4(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n623), .A2(new_n626), .A3(new_n540), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n659), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n808), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n823), .A2(KEYINPUT116), .A3(new_n784), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n359), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n312), .B1(new_n871), .B2(new_n813), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT117), .B(new_n867), .C1(new_n872), .C2(new_n816), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n838), .A2(new_n518), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n685), .B1(new_n808), .B2(new_n868), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n829), .B1(new_n878), .B2(new_n870), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n832), .B1(new_n879), .B2(new_n312), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT117), .B1(new_n880), .B2(new_n867), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n273), .B(new_n865), .C1(new_n877), .C2(new_n881), .ZN(new_n882));
  AOI211_X1 g681(.A(KEYINPUT119), .B(new_n863), .C1(G141gat), .C2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(G141gat), .ZN(new_n885));
  INV_X1    g684(.A(new_n863), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n860), .A2(new_n540), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n817), .A2(new_n857), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(new_n882), .B2(G141gat), .ZN(new_n890));
  OAI22_X1  g689(.A1(new_n883), .A2(new_n887), .B1(new_n862), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI221_X1 g692(.A(KEYINPUT120), .B1(new_n862), .B2(new_n890), .C1(new_n883), .C2(new_n887), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1344gat));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n865), .B1(new_n877), .B2(new_n881), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n896), .B(G148gat), .C1(new_n897), .C2(new_n381), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n811), .A2(new_n685), .A3(new_n812), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n878), .B2(new_n870), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n901), .A2(new_n312), .B1(new_n273), .B2(new_n382), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n902), .B2(new_n518), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n903), .A2(KEYINPUT121), .B1(new_n874), .B2(new_n875), .ZN(new_n904));
  INV_X1    g703(.A(new_n900), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n871), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n815), .B1(new_n906), .B2(new_n712), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n866), .B1(new_n907), .B2(new_n659), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n648), .B(new_n865), .C1(new_n904), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G148gat), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n899), .B1(new_n912), .B2(KEYINPUT59), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT122), .B(new_n896), .C1(new_n911), .C2(G148gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n898), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n858), .A2(new_n859), .A3(new_n540), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n916), .A2(G148gat), .A3(new_n381), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n897), .B2(new_n712), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n312), .A2(new_n307), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n916), .B2(new_n920), .ZN(G1346gat));
  NOR3_X1   g720(.A1(new_n916), .A2(G162gat), .A3(new_n359), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT123), .Z(new_n923));
  OAI21_X1  g722(.A(G162gat), .B1(new_n897), .B2(new_n668), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n626), .A2(new_n540), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n480), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n838), .A2(new_n659), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(G169gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(new_n274), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n839), .A2(new_n581), .A3(new_n927), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT124), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n273), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n930), .ZN(G1348gat));
  INV_X1    g735(.A(G176gat), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n929), .A2(new_n937), .A3(new_n381), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n648), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n937), .ZN(G1349gat));
  OR2_X1    g739(.A1(new_n929), .A2(new_n712), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n312), .A2(new_n421), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n941), .A2(G183gat), .B1(new_n932), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT125), .B(KEYINPUT60), .Z(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1350gat));
  AOI21_X1  g744(.A(new_n422), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n929), .B2(new_n359), .ZN(new_n947));
  NOR2_X1   g746(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n947), .B(new_n948), .Z(new_n949));
  NAND2_X1  g748(.A1(new_n667), .A2(new_n422), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n933), .B2(new_n950), .ZN(G1351gat));
  NAND2_X1  g750(.A1(new_n623), .A2(new_n926), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(new_n874), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n273), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n874), .A2(new_n875), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n908), .B2(new_n909), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n903), .A2(KEYINPUT121), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n273), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  INV_X1    g759(.A(new_n958), .ZN(new_n961));
  OAI21_X1  g760(.A(G204gat), .B1(new_n961), .B2(new_n381), .ZN(new_n962));
  INV_X1    g761(.A(new_n953), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n963), .A2(G204gat), .A3(new_n381), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(G1353gat));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n967));
  INV_X1    g766(.A(new_n952), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n312), .B(new_n968), .C1(new_n904), .C2(new_n910), .ZN(new_n969));
  OAI21_X1  g768(.A(G211gat), .B1(new_n969), .B2(KEYINPUT127), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n971), .B1(new_n958), .B2(new_n312), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n967), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n971), .A3(new_n312), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  OR3_X1    g776(.A1(new_n963), .A2(G211gat), .A3(new_n712), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1354gat));
  OAI21_X1  g778(.A(G218gat), .B1(new_n961), .B2(new_n359), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n668), .A2(G218gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n963), .B2(new_n981), .ZN(G1355gat));
endmodule


