//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G125), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT16), .A3(G140), .ZN(new_n189));
  XNOR2_X1  g003(.A(G125), .B(G140), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OR3_X1    g014(.A1(new_n196), .A2(KEYINPUT23), .A3(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT23), .B1(new_n196), .B2(G128), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n195), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G110), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n200), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n193), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT74), .B(G110), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n198), .B2(new_n199), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n191), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n190), .A2(new_n192), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT22), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n216), .B(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(KEYINPUT75), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n206), .A2(new_n212), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G902), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n187), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI211_X1 g039(.A(KEYINPUT25), .B(G902), .C1(new_n219), .C2(new_n222), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(G234), .B2(new_n224), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G902), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n227), .A2(new_n229), .B1(new_n223), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(G116), .B(G119), .Z(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT2), .B(G113), .Z(new_n237));
  XNOR2_X1  g051(.A(G116), .B(G119), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n238), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(KEYINPUT67), .A3(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n236), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n239), .B1(new_n236), .B2(new_n242), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT30), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(new_n249), .A3(new_n217), .A4(G134), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  OAI22_X1  g065(.A1(new_n251), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI22_X1  g067(.A1(new_n248), .A2(new_n249), .B1(new_n217), .B2(G134), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(G131), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n251), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n217), .B2(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n251), .A2(KEYINPUT66), .A3(G137), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n257), .B(new_n258), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n247), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n194), .A2(new_n192), .A3(G143), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n265), .B(G146), .C1(new_n194), .C2(KEYINPUT1), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n192), .A2(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G128), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n264), .B(new_n266), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G131), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n254), .B1(new_n252), .B2(new_n250), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n274), .B(KEYINPUT69), .C1(new_n275), .C2(G131), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n263), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n253), .A2(new_n255), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n279), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G128), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n269), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G143), .B(G146), .ZN(new_n286));
  NAND2_X1  g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n246), .B1(new_n277), .B2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n280), .A2(new_n282), .B1(new_n285), .B2(new_n288), .ZN(new_n292));
  INV_X1    g106(.A(new_n272), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n278), .A2(new_n257), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n274), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n292), .A2(new_n295), .A3(KEYINPUT30), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n245), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n239), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n241), .B1(new_n240), .B2(KEYINPUT67), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n300));
  AOI211_X1 g114(.A(new_n300), .B(KEYINPUT68), .C1(new_n237), .C2(new_n238), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n236), .A2(new_n239), .A3(new_n242), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n290), .A3(new_n277), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(G101), .ZN(new_n308));
  NOR2_X1   g122(.A1(G237), .A2(G953), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G210), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n308), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT29), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n302), .B(new_n303), .C1(new_n292), .C2(new_n295), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT28), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n277), .A2(new_n290), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(new_n245), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n305), .A2(KEYINPUT71), .A3(new_n317), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n311), .B(KEYINPUT70), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n316), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n313), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n313), .A2(new_n324), .A3(KEYINPUT72), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n224), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n305), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n304), .B1(new_n290), .B2(new_n277), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT28), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n332), .A2(new_n321), .A3(new_n322), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n333), .A2(KEYINPUT73), .A3(KEYINPUT29), .A4(new_n311), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(KEYINPUT29), .A3(new_n321), .A4(new_n322), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n312), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G472), .B1(new_n329), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(G472), .A2(G902), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n297), .A2(new_n305), .A3(new_n311), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n297), .A2(KEYINPUT31), .A3(new_n305), .A4(new_n311), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n316), .A2(new_n321), .A3(new_n322), .ZN(new_n347));
  INV_X1    g161(.A(new_n323), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n341), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n344), .A2(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n352), .A2(new_n353), .A3(new_n341), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n232), .B1(new_n339), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G214), .B1(G237), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n196), .A3(G116), .ZN(new_n360));
  OAI211_X1 g174(.A(G113), .B(new_n360), .C1(new_n233), .C2(new_n359), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n240), .ZN(new_n362));
  NOR2_X1   g176(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n363));
  INV_X1    g177(.A(G107), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(G104), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G104), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n366), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n367));
  OAI22_X1  g181(.A1(new_n366), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n368));
  INV_X1    g182(.A(G101), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n365), .A2(new_n367), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n364), .A2(G104), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n366), .A2(G107), .ZN(new_n372));
  OAI21_X1  g186(.A(G101), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n362), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n370), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n379), .A3(G101), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n375), .B1(new_n304), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(KEYINPUT81), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n384), .B(new_n375), .C1(new_n304), .C2(new_n381), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n289), .A2(G125), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(G125), .B2(new_n293), .ZN(new_n390));
  INV_X1    g204(.A(G224), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G953), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n392), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n382), .A2(new_n396), .A3(new_n385), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n388), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n393), .B(new_n394), .C1(KEYINPUT7), .C2(new_n392), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n362), .B(new_n374), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n384), .B(KEYINPUT8), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OR3_X1    g216(.A1(new_n390), .A2(KEYINPUT7), .A3(new_n392), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n399), .A2(new_n387), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n224), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G210), .B1(G237), .B2(G902), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n398), .A2(new_n224), .A3(new_n406), .A4(new_n404), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n358), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT9), .B(G234), .Z(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT76), .ZN(new_n412));
  OAI21_X1  g226(.A(G221), .B1(new_n412), .B2(G902), .ZN(new_n413));
  INV_X1    g227(.A(G469), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n272), .A2(new_n373), .A3(new_n370), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT10), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n272), .A2(KEYINPUT10), .A3(new_n373), .A4(new_n370), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n378), .A2(new_n289), .A3(new_n380), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT78), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT78), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n378), .A2(new_n289), .A3(new_n422), .A4(new_n380), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n283), .B(new_n419), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G140), .ZN(new_n425));
  INV_X1    g239(.A(G227), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G953), .ZN(new_n427));
  XOR2_X1   g241(.A(new_n425), .B(new_n427), .Z(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT79), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n283), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n423), .ZN(new_n432));
  INV_X1    g246(.A(new_n419), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n431), .A3(new_n433), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT79), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n428), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n430), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n293), .A2(new_n374), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n415), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n441), .A2(KEYINPUT12), .A3(new_n283), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT12), .B1(new_n441), .B2(new_n283), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n429), .B1(new_n424), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT80), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n439), .A2(KEYINPUT80), .A3(new_n445), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n414), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n414), .A2(new_n224), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n429), .B1(new_n434), .B2(new_n424), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n436), .B(new_n428), .C1(new_n442), .C2(new_n443), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n454), .B2(new_n414), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n410), .B(new_n413), .C1(new_n450), .C2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G113), .B(G122), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n366), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n309), .A2(G214), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n265), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n309), .A2(G143), .A3(G214), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G131), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n257), .A3(new_n463), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(KEYINPUT17), .A3(G131), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n193), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n190), .B(new_n192), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT82), .A2(KEYINPUT18), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(new_n257), .ZN(new_n473));
  OAI221_X1 g287(.A(new_n471), .B1(new_n464), .B2(new_n473), .C1(new_n465), .C2(new_n472), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n460), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(KEYINPUT85), .B(new_n460), .C1(new_n470), .C2(new_n474), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n460), .B(KEYINPUT84), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n470), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G475), .B1(new_n481), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(G475), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n465), .A2(new_n467), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT19), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT83), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n485), .A2(KEYINPUT83), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n190), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(G125), .A2(G140), .ZN(new_n489));
  NAND2_X1  g303(.A1(G125), .A2(G140), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(KEYINPUT83), .A3(new_n485), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n192), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n210), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n460), .B1(new_n474), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n483), .B(new_n224), .C1(new_n480), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT20), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n470), .A2(new_n479), .A3(new_n474), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n474), .A2(new_n494), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n460), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(KEYINPUT20), .A3(new_n483), .A4(new_n224), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n482), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n194), .B2(G143), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT86), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n194), .A2(G143), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n265), .A2(G128), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT86), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n504), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n265), .A2(KEYINPUT13), .A3(G128), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT88), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n506), .A2(new_n510), .A3(KEYINPUT87), .A4(new_n507), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G134), .ZN(new_n518));
  XNOR2_X1  g332(.A(G116), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n364), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n508), .A2(new_n507), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n251), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n521), .B(new_n251), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n519), .A2(new_n364), .ZN(new_n527));
  INV_X1    g341(.A(G116), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT14), .A3(G122), .ZN(new_n529));
  INV_X1    g343(.A(new_n519), .ZN(new_n530));
  OAI211_X1 g344(.A(G107), .B(new_n529), .C1(new_n530), .C2(KEYINPUT14), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(KEYINPUT89), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n523), .B1(new_n517), .B2(G134), .ZN(new_n535));
  INV_X1    g349(.A(new_n532), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n412), .A2(new_n228), .A3(G953), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n533), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n534), .B(new_n538), .C1(new_n535), .C2(new_n536), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n224), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  OR2_X1    g357(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n544));
  NAND2_X1  g358(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n542), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G952), .ZN(new_n548));
  AOI211_X1 g362(.A(G953), .B(new_n548), .C1(G234), .C2(G237), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT21), .B(G898), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT91), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI211_X1 g366(.A(new_n224), .B(new_n214), .C1(G234), .C2(G237), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n503), .A2(new_n547), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n356), .A2(new_n458), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(G101), .ZN(G3));
  INV_X1    g371(.A(new_n413), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n439), .A2(KEYINPUT80), .A3(new_n445), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT80), .B1(new_n439), .B2(new_n445), .ZN(new_n560));
  OAI21_X1  g374(.A(G469), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n561), .B2(new_n455), .ZN(new_n562));
  OAI21_X1  g376(.A(G472), .B1(new_n352), .B2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n350), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n562), .A2(new_n231), .A3(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n358), .B(new_n554), .C1(new_n408), .C2(new_n409), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT33), .B1(new_n540), .B2(new_n541), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT92), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n525), .B(new_n532), .C1(new_n570), .C2(new_n538), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n539), .B(KEYINPUT92), .C1(new_n535), .C2(new_n536), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(G478), .B(new_n224), .C1(new_n568), .C2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n542), .A2(new_n575), .A3(new_n543), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n542), .B2(new_n543), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n498), .A2(new_n502), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n477), .A2(new_n478), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n224), .B1(new_n581), .B2(new_n480), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n582), .B2(G475), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n567), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n566), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT34), .B(G104), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G6));
  AND2_X1   g402(.A1(new_n583), .A2(new_n547), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n567), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n566), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT35), .B(G107), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT94), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(G9));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n220), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT95), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n597), .A2(new_n221), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n221), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n230), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n227), .A2(new_n229), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n458), .A2(new_n555), .A3(new_n565), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT37), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(new_n204), .ZN(G12));
  AND2_X1   g419(.A1(new_n600), .A2(new_n601), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n339), .B2(new_n355), .ZN(new_n607));
  INV_X1    g421(.A(new_n549), .ZN(new_n608));
  INV_X1    g422(.A(new_n553), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(G900), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(KEYINPUT96), .Z(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n589), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n607), .A2(new_n458), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G128), .ZN(G30));
  NAND2_X1  g429(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n353), .B1(new_n352), .B2(new_n341), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n348), .B1(new_n330), .B2(new_n331), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n618), .A2(new_n342), .ZN(new_n619));
  OAI21_X1  g433(.A(G472), .B1(new_n619), .B2(G902), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT97), .A4(new_n620), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n503), .A2(new_n547), .A3(new_n357), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n611), .B(KEYINPUT39), .Z(new_n627));
  OAI211_X1 g441(.A(new_n413), .B(new_n627), .C1(new_n450), .C2(new_n456), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT98), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n562), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n626), .B1(new_n632), .B2(KEYINPUT40), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n629), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n408), .A2(new_n409), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT38), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n633), .A2(new_n606), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G143), .ZN(G45));
  NAND3_X1  g453(.A1(new_n578), .A2(new_n503), .A3(new_n612), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT99), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n607), .A2(new_n641), .A3(new_n458), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G146), .ZN(G48));
  NAND2_X1  g457(.A1(new_n452), .A2(new_n453), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n224), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G469), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n454), .A2(new_n414), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n413), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n356), .A2(new_n585), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT41), .B(G113), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G15));
  NAND3_X1  g467(.A1(new_n356), .A2(new_n590), .A3(new_n650), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G116), .ZN(G18));
  AND3_X1   g469(.A1(new_n410), .A2(new_n648), .A3(new_n413), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n607), .A2(new_n555), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G119), .ZN(G21));
  OAI21_X1  g472(.A(new_n346), .B1(new_n333), .B2(new_n323), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n340), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n563), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT100), .B1(new_n661), .B2(new_n232), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n231), .A2(new_n563), .A3(new_n660), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n625), .A2(new_n636), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n649), .A2(new_n554), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G122), .ZN(G24));
  NOR2_X1   g483(.A1(new_n606), .A2(new_n661), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n641), .A2(new_n656), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G125), .ZN(G27));
  AND2_X1   g486(.A1(new_n616), .A2(KEYINPUT104), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n616), .A2(KEYINPUT104), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n673), .A2(new_n674), .A3(new_n351), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n232), .B1(new_n675), .B2(new_n339), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n408), .A2(new_n357), .A3(new_n409), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n439), .A2(G469), .A3(new_n445), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n558), .B1(new_n455), .B2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n408), .A2(KEYINPUT101), .A3(new_n357), .A4(new_n409), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n676), .A2(KEYINPUT42), .A3(new_n641), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n356), .A2(new_n683), .A3(new_n641), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n687));
  AND3_X1   g501(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G131), .ZN(G33));
  AND2_X1   g505(.A1(new_n356), .A2(new_n683), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n613), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G134), .ZN(G36));
  INV_X1    g508(.A(new_n647), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n448), .A2(new_n696), .A3(new_n449), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n439), .A2(KEYINPUT45), .A3(new_n445), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(G469), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n451), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n695), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n699), .A2(KEYINPUT46), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n679), .A2(new_n682), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n705), .A2(new_n413), .A3(new_n627), .A4(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n565), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n542), .A2(new_n543), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT93), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n542), .A2(new_n575), .A3(new_n543), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n503), .B1(new_n714), .B2(new_n574), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n710), .B1(new_n715), .B2(KEYINPUT43), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n578), .A2(new_n583), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(KEYINPUT105), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n578), .A2(KEYINPUT43), .A3(new_n583), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n578), .A2(new_n583), .A3(new_n722), .A4(KEYINPUT43), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n716), .A2(new_n719), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n709), .B(new_n602), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n722), .B1(new_n715), .B2(KEYINPUT43), .ZN(new_n727));
  INV_X1    g541(.A(new_n723), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT105), .B1(new_n717), .B2(new_n718), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n710), .B(KEYINPUT43), .C1(new_n578), .C2(new_n583), .ZN(new_n730));
  OAI22_X1  g544(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT44), .B1(new_n726), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n565), .B1(new_n731), .B2(KEYINPUT107), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n724), .A2(new_n725), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n735), .A3(new_n602), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n708), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n217), .ZN(G39));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n701), .A2(new_n702), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n741), .A2(new_n647), .A3(new_n704), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n742), .B2(new_n558), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n705), .A2(KEYINPUT47), .A3(new_n413), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n355), .A2(new_n707), .A3(new_n339), .A4(new_n232), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n641), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G140), .ZN(G42));
  INV_X1    g562(.A(new_n648), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(KEYINPUT49), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(KEYINPUT49), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n357), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n637), .A3(new_n232), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n623), .A2(new_n624), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n413), .A3(new_n754), .A4(new_n715), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n607), .B(new_n458), .C1(new_n641), .C2(new_n613), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n600), .A2(KEYINPUT110), .A3(new_n601), .A4(new_n612), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n757), .A2(new_n636), .A3(new_n625), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n602), .B2(new_n611), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(new_n621), .A3(new_n681), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n756), .A2(new_n671), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT52), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n756), .A2(new_n764), .A3(new_n761), .A4(new_n671), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n763), .A2(new_n765), .B1(KEYINPUT111), .B2(new_n762), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(KEYINPUT111), .A3(new_n764), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n578), .A2(KEYINPUT108), .A3(new_n503), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT108), .B1(new_n578), .B2(new_n503), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n567), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT109), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n567), .B(new_n774), .C1(new_n770), .C2(new_n771), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n566), .A3(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(new_n556), .A3(new_n591), .A4(new_n603), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n503), .A2(new_n547), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n562), .A2(new_n607), .A3(new_n780), .A4(new_n612), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n641), .A2(new_n670), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n781), .A2(new_n707), .B1(new_n782), .B2(new_n683), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n690), .A2(new_n779), .A3(new_n693), .A4(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n668), .A2(new_n651), .A3(new_n654), .A4(new_n657), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT115), .Z(new_n786));
  NAND3_X1  g600(.A1(new_n769), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n777), .A2(new_n785), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n690), .A2(new_n791), .A3(new_n693), .A4(new_n783), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n763), .A2(new_n765), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n787), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n724), .A2(new_n608), .A3(new_n649), .A4(new_n706), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n676), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT48), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n548), .A2(G953), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n706), .A2(new_n232), .A3(new_n649), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n549), .A3(new_n754), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n584), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n798), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n724), .A2(new_n608), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(new_n665), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n803), .B1(new_n656), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n648), .A2(new_n558), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n743), .A2(new_n744), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n805), .A2(new_n707), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n650), .A2(new_n358), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n637), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n805), .A2(KEYINPUT50), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n804), .A2(new_n665), .A3(new_n813), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n818), .B1(new_n819), .B2(new_n815), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n801), .A2(new_n583), .A3(new_n579), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n796), .A2(new_n670), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n810), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n824), .A2(KEYINPUT51), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(KEYINPUT51), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n806), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n685), .A2(new_n687), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT103), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n831), .A2(new_n684), .B1(new_n613), .B2(new_n692), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n781), .A2(new_n707), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n782), .A2(new_n683), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n777), .A3(new_n785), .ZN(new_n836));
  INV_X1    g650(.A(new_n793), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n832), .A2(new_n836), .A3(new_n789), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n690), .A2(new_n791), .A3(new_n693), .A4(new_n783), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n789), .A4(new_n837), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(KEYINPUT112), .B(KEYINPUT53), .C1(new_n769), .C2(new_n840), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n793), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n832), .A2(new_n847), .A3(new_n836), .A4(new_n767), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n845), .B1(new_n848), .B2(new_n778), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n843), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n795), .B(new_n827), .C1(new_n850), .C2(KEYINPUT54), .ZN(new_n851));
  NOR2_X1   g665(.A1(G952), .A2(G953), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n755), .B1(new_n851), .B2(new_n852), .ZN(G75));
  NAND2_X1  g667(.A1(new_n787), .A2(new_n794), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(G210), .A3(G902), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n388), .A2(new_n397), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(new_n395), .Z(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT55), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(KEYINPUT117), .B2(new_n856), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n855), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(new_n855), .B2(new_n856), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n214), .A2(G952), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G51));
  NAND2_X1  g678(.A1(new_n700), .A2(KEYINPUT57), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n788), .B1(new_n787), .B2(new_n794), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n795), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n700), .A2(KEYINPUT57), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n644), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n854), .A2(G902), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(new_n699), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n863), .B1(new_n869), .B2(new_n871), .ZN(G54));
  NAND4_X1  g686(.A1(new_n854), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n873));
  INV_X1    g687(.A(new_n501), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n876), .A3(new_n863), .ZN(G60));
  NOR2_X1   g691(.A1(new_n568), .A2(new_n573), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(G478), .A2(G902), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT59), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n879), .B(new_n881), .C1(new_n795), .C2(new_n866), .ZN(new_n882));
  INV_X1    g696(.A(new_n863), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n792), .A2(new_n768), .A3(new_n766), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT112), .B1(new_n885), .B2(KEYINPUT53), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n848), .A2(new_n845), .A3(new_n778), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n788), .B1(new_n888), .B2(new_n843), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n881), .B1(new_n889), .B2(new_n795), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n884), .B1(new_n890), .B2(new_n878), .ZN(G63));
  NAND2_X1  g705(.A1(G217), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT60), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n854), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n223), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n863), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n854), .A2(new_n598), .A3(new_n599), .A4(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT61), .B1(new_n898), .B2(KEYINPUT118), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n897), .B(new_n898), .C1(KEYINPUT118), .C2(KEYINPUT61), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G66));
  OAI21_X1  g717(.A(G953), .B1(new_n552), .B2(new_n391), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n791), .B2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n857), .B1(G898), .B2(new_n214), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(G69));
  OR2_X1    g721(.A1(new_n291), .A2(new_n296), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n492), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n733), .A2(new_n737), .ZN(new_n910));
  INV_X1    g724(.A(new_n708), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n756), .A2(new_n671), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(KEYINPUT122), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n738), .B2(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n705), .A2(new_n413), .A3(new_n627), .A4(new_n666), .ZN(new_n919));
  INV_X1    g733(.A(new_n676), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT123), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n627), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n558), .B(new_n922), .C1(new_n703), .C2(new_n704), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(new_n924), .A3(new_n666), .A4(new_n676), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n832), .A2(new_n747), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(G953), .B1(new_n918), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n214), .A2(G900), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n909), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  INV_X1    g745(.A(new_n356), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n770), .A2(new_n771), .A3(new_n589), .ZN(new_n933));
  NOR4_X1   g747(.A1(new_n632), .A2(new_n932), .A3(new_n706), .A4(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n912), .A2(KEYINPUT119), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n738), .B2(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n638), .A2(new_n914), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n638), .A2(KEYINPUT62), .A3(new_n914), .ZN(new_n943));
  INV_X1    g757(.A(new_n641), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n743), .B2(new_n744), .ZN(new_n945));
  AOI22_X1  g759(.A1(new_n942), .A2(new_n943), .B1(new_n945), .B2(new_n746), .ZN(new_n946));
  AOI21_X1  g760(.A(G953), .B1(new_n939), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n931), .B1(new_n947), .B2(new_n909), .ZN(new_n948));
  INV_X1    g762(.A(new_n909), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n638), .A2(KEYINPUT62), .A3(new_n914), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT62), .B1(new_n638), .B2(new_n914), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n747), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n938), .B2(new_n936), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT120), .B(new_n949), .C1(new_n953), .C2(G953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n930), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n929), .B1(new_n426), .B2(G953), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT121), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n930), .A2(new_n948), .A3(new_n954), .A4(new_n957), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(G72));
  NAND3_X1  g775(.A1(new_n918), .A2(new_n927), .A3(new_n791), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT125), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n306), .A2(new_n311), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n962), .A2(new_n968), .A3(new_n964), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n964), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n953), .B2(new_n791), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n306), .A2(new_n311), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n967), .A3(new_n971), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT126), .Z(new_n979));
  AOI21_X1  g793(.A(new_n863), .B1(new_n850), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT124), .B1(new_n972), .B2(new_n975), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n970), .A2(new_n977), .A3(new_n980), .A4(new_n981), .ZN(G57));
endmodule


