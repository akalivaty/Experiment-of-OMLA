//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT3), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT79), .B1(new_n193), .B2(G104), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n191), .A3(G107), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT4), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n197), .A2(new_n199), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n196), .B1(new_n202), .B2(new_n195), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G116), .B(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT2), .A2(G113), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT2), .A3(G113), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT2), .A2(G113), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n207), .A2(new_n209), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G116), .ZN(new_n216));
  INV_X1    g030(.A(G116), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G119), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n213), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n210), .A2(KEYINPUT67), .A3(new_n205), .A4(new_n211), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n212), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI211_X1 g036(.A(KEYINPUT4), .B(new_n196), .C1(new_n202), .C2(new_n195), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n204), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT5), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n215), .A3(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G113), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(KEYINPUT5), .B2(new_n205), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(new_n220), .B2(new_n221), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n191), .A2(G107), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n193), .A2(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n200), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n189), .B1(new_n224), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n222), .ZN(new_n238));
  INV_X1    g052(.A(new_n203), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT4), .A3(new_n200), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G101), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n188), .A3(new_n235), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n237), .A2(new_n245), .A3(KEYINPUT6), .ZN(new_n246));
  INV_X1    g060(.A(G125), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G146), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n248), .B(new_n249), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(G146), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT0), .A4(G128), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n247), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT1), .B1(new_n250), .B2(G146), .ZN(new_n259));
  OAI211_X1 g073(.A(G128), .B(new_n259), .C1(new_n251), .C2(new_n253), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n255), .B(new_n256), .C1(KEYINPUT1), .C2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(G125), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT83), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n265));
  XNOR2_X1  g079(.A(G143), .B(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n249), .A2(new_n248), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n257), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n265), .B1(new_n269), .B2(new_n247), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G224), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n273), .B(KEYINPUT84), .Z(new_n274));
  XOR2_X1   g088(.A(new_n271), .B(new_n274), .Z(new_n275));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(new_n189), .C1(new_n224), .C2(new_n236), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n246), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n264), .A2(new_n270), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n258), .B2(new_n263), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n222), .A2(new_n223), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n284), .A2(new_n240), .B1(new_n234), .B2(new_n229), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n188), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n229), .A2(new_n234), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n188), .B(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n235), .A2(KEYINPUT85), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n289), .B(new_n290), .C1(new_n291), .C2(new_n287), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n187), .B1(new_n278), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT86), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n278), .A2(new_n293), .A3(new_n187), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n278), .A2(new_n293), .A3(KEYINPUT87), .A4(new_n187), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n243), .B(new_n269), .C1(new_n201), .C2(new_n203), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n260), .A2(new_n262), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n308), .A2(KEYINPUT10), .A3(new_n200), .A4(new_n232), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n200), .A2(new_n262), .A3(new_n260), .A4(new_n232), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT11), .ZN(new_n314));
  INV_X1    g128(.A(G134), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G137), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT11), .A3(G134), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(G137), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G131), .ZN(new_n321));
  INV_X1    g135(.A(G131), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n316), .A2(new_n318), .A3(new_n322), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n313), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n324), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n306), .A2(new_n309), .A3(new_n312), .A4(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G110), .B(G140), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT77), .ZN(new_n329));
  INV_X1    g143(.A(G227), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G953), .ZN(new_n331));
  XOR2_X1   g145(.A(new_n329), .B(new_n331), .Z(new_n332));
  NAND3_X1  g146(.A1(new_n325), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n233), .A2(new_n307), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n326), .B1(new_n334), .B2(new_n310), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(KEYINPUT12), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT12), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n337), .B(new_n326), .C1(new_n334), .C2(new_n310), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT80), .B(new_n327), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n332), .B(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n310), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n200), .A2(new_n232), .B1(new_n262), .B2(new_n260), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n324), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n337), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n335), .A2(KEYINPUT12), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT80), .B1(new_n347), .B2(new_n327), .ZN(new_n348));
  OAI211_X1 g162(.A(G469), .B(new_n333), .C1(new_n341), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(G469), .A2(G902), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n332), .B1(new_n325), .B2(new_n327), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n352), .A2(KEYINPUT82), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n327), .A2(new_n332), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n327), .A2(KEYINPUT81), .A3(new_n332), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n347), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n352), .A2(KEYINPUT82), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G469), .ZN(new_n361));
  INV_X1    g175(.A(G902), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n305), .B1(new_n351), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(G234), .A2(G237), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(G952), .A3(new_n272), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT21), .B(G898), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(G902), .A3(G953), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G214), .B1(G237), .B2(G902), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n302), .A2(new_n364), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(G475), .A2(G902), .ZN(new_n374));
  INV_X1    g188(.A(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n247), .A2(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G146), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n252), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT88), .ZN(new_n382));
  OR3_X1    g196(.A1(new_n380), .A2(KEYINPUT88), .A3(new_n252), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(G237), .A2(G953), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G214), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n250), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(G143), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT18), .A3(G131), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT18), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n387), .B(new_n388), .C1(new_n391), .C2(new_n322), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT89), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n392), .A2(new_n393), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n384), .B(new_n390), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n389), .A2(G131), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n387), .A2(new_n322), .A3(new_n388), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT16), .ZN(new_n401));
  OR3_X1    g215(.A1(new_n247), .A2(KEYINPUT16), .A3(G140), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G146), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(G146), .B1(new_n401), .B2(new_n402), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n400), .B(new_n406), .C1(new_n398), .C2(new_n397), .ZN(new_n407));
  XNOR2_X1  g221(.A(G113), .B(G122), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(new_n191), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n396), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n397), .A2(new_n399), .ZN(new_n411));
  NAND2_X1  g225(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n380), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n380), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n411), .B(new_n403), .C1(G146), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n409), .B1(new_n396), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n374), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT20), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(new_n374), .C1(new_n410), .C2(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n409), .B1(new_n396), .B2(new_n407), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n362), .B1(new_n410), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G475), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G122), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G116), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n217), .A2(G122), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G107), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n429), .A3(new_n193), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT13), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n261), .B2(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n261), .A2(G143), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n250), .A2(G128), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(new_n434), .ZN(new_n439));
  OAI21_X1  g253(.A(G134), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n436), .A3(new_n315), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n433), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G134), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n441), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n217), .A2(KEYINPUT14), .A3(G122), .ZN(new_n446));
  OAI211_X1 g260(.A(G107), .B(new_n446), .C1(new_n430), .C2(KEYINPUT14), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n432), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n303), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(G217), .A3(new_n272), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n442), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n442), .B2(new_n448), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n362), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G478), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n442), .A2(new_n448), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n450), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n442), .A2(new_n448), .A3(new_n451), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n456), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n362), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n426), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n373), .A2(KEYINPUT91), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G234), .ZN(new_n469));
  OAI21_X1  g283(.A(G217), .B1(new_n469), .B2(G902), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT71), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT72), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT22), .B(G137), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n215), .A2(G128), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n261), .A2(KEYINPUT23), .A3(G119), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n215), .A2(G128), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(KEYINPUT23), .ZN(new_n479));
  XNOR2_X1  g293(.A(G119), .B(G128), .ZN(new_n480));
  INV_X1    g294(.A(G110), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT24), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G110), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n479), .A2(G110), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n404), .B2(new_n405), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n479), .A2(G110), .B1(new_n480), .B2(new_n485), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n403), .A3(new_n381), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT73), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT73), .B1(new_n487), .B2(new_n489), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n475), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n489), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT73), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n475), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n362), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT74), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT74), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n492), .A2(new_n502), .A3(new_n497), .A4(new_n362), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n498), .A2(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT25), .B1(new_n498), .B2(KEYINPUT74), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n500), .B1(new_n507), .B2(new_n503), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n471), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n471), .A2(G902), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT76), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n492), .A2(new_n497), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n315), .A2(G137), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n317), .A2(G134), .ZN(new_n515));
  OAI21_X1  g329(.A(G131), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n323), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n323), .A2(new_n516), .A3(KEYINPUT68), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n308), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n269), .A2(new_n324), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(KEYINPUT30), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT69), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n521), .A2(new_n525), .A3(KEYINPUT30), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n307), .A2(new_n517), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n268), .B1(new_n323), .B2(new_n321), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT64), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n522), .A2(KEYINPUT64), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT65), .B(new_n528), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n522), .A2(KEYINPUT64), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(new_n531), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n529), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT65), .B1(new_n538), .B2(new_n528), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n238), .B(new_n527), .C1(new_n535), .C2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n521), .A2(new_n222), .A3(new_n522), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n385), .A2(G210), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT27), .Z(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT31), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n238), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n541), .A2(KEYINPUT28), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n541), .A2(KEYINPUT28), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n545), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT31), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n540), .A2(new_n554), .A3(new_n541), .A4(new_n546), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n548), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(G472), .A2(G902), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT70), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT32), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n222), .B1(new_n521), .B2(new_n522), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n550), .B2(new_n551), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT29), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n564), .A2(new_n565), .A3(new_n545), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G902), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n546), .B1(new_n540), .B2(new_n541), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n565), .B1(new_n552), .B2(new_n545), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n556), .A2(new_n561), .B1(new_n570), .B2(G472), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n513), .B1(new_n560), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n302), .A2(new_n467), .A3(new_n364), .A4(new_n372), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n468), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  NAND2_X1  g391(.A1(new_n556), .A2(new_n362), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G472), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n556), .A2(new_n558), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n513), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n278), .A2(new_n293), .ZN(new_n583));
  INV_X1    g397(.A(new_n187), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n297), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n370), .A3(new_n371), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n422), .A2(new_n425), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT33), .B1(new_n451), .B2(KEYINPUT92), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n461), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n461), .A2(new_n589), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n455), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n455), .A2(new_n362), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n454), .B2(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n587), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n582), .A2(new_n364), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  NAND3_X1  g415(.A1(new_n422), .A2(new_n464), .A3(new_n425), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n587), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n582), .A2(new_n364), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  AOI22_X1  g420(.A1(new_n578), .A2(G472), .B1(new_n558), .B2(new_n556), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n475), .A2(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT94), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT93), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n608), .A2(KEYINPUT94), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(KEYINPUT94), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n493), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n610), .B2(new_n614), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n511), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n509), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n468), .A2(new_n575), .A3(new_n607), .A4(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT37), .B(G110), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G12));
  NAND2_X1  g436(.A1(new_n556), .A2(new_n561), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n570), .A2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n371), .B(new_n586), .C1(new_n625), .C2(new_n559), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n369), .A2(G900), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n366), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n426), .A2(KEYINPUT95), .A3(new_n464), .A4(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n630));
  INV_X1    g444(.A(new_n628), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n630), .B1(new_n602), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n364), .A3(new_n619), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n261), .ZN(G30));
  XNOR2_X1  g450(.A(new_n628), .B(KEYINPUT39), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n364), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n302), .B(KEYINPUT38), .ZN(new_n641));
  INV_X1    g455(.A(new_n619), .ZN(new_n642));
  INV_X1    g456(.A(new_n371), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n465), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n588), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n541), .A2(new_n545), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n646), .B2(new_n563), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n540), .A2(new_n541), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(new_n545), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n556), .A2(new_n561), .B1(new_n649), .B2(G472), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n645), .B1(new_n560), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n640), .A2(new_n641), .A3(new_n642), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G143), .ZN(G45));
  INV_X1    g467(.A(new_n626), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n597), .A2(new_n631), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n619), .A2(new_n364), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G146), .ZN(G48));
  NAND2_X1  g472(.A1(new_n360), .A2(new_n362), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(KEYINPUT96), .A3(G469), .ZN(new_n660));
  NAND2_X1  g474(.A1(KEYINPUT96), .A2(G469), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n360), .A2(new_n362), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n304), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n572), .A2(new_n598), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT41), .B(G113), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G15));
  NAND3_X1  g481(.A1(new_n572), .A2(new_n603), .A3(new_n664), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G116), .ZN(G18));
  NOR3_X1   g483(.A1(new_n663), .A2(new_n587), .A3(new_n466), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n560), .A2(new_n571), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n619), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G119), .ZN(G21));
  XOR2_X1   g487(.A(KEYINPUT98), .B(G472), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n578), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n546), .B1(new_n564), .B2(KEYINPUT97), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(KEYINPUT97), .B2(new_n564), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n548), .A2(new_n555), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n558), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n513), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n586), .A2(new_n588), .A3(new_n370), .A4(new_n644), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n663), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  NAND4_X1  g499(.A1(new_n675), .A2(new_n619), .A3(new_n655), .A4(new_n679), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT99), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n586), .A2(new_n371), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n663), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n663), .A2(new_n689), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT99), .B1(new_n692), .B2(new_n686), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n585), .A2(new_n295), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n294), .A2(KEYINPUT86), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n301), .A2(new_n697), .A3(new_n698), .A4(new_n371), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT101), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n296), .A2(new_n701), .A3(new_n301), .A4(new_n371), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n333), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n333), .A2(new_n703), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n704), .B(new_n705), .C1(new_n348), .C2(new_n341), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n361), .B1(new_n706), .B2(new_n362), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n305), .B1(new_n708), .B2(new_n363), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n700), .A2(new_n702), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n655), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n623), .B(KEYINPUT102), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n559), .B1(G472), .B2(new_n570), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n513), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n696), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n681), .B1(new_n625), .B2(new_n559), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n710), .A2(new_n718), .A3(KEYINPUT42), .A4(new_n711), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n322), .ZN(G33));
  NOR2_X1   g536(.A1(new_n710), .A2(new_n718), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n633), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n726), .B1(new_n706), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n704), .A2(new_n705), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n341), .A2(new_n348), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(KEYINPUT103), .A3(KEYINPUT45), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n333), .B1(new_n341), .B2(new_n348), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n361), .B1(new_n732), .B2(new_n727), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n350), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n350), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n363), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n304), .A3(new_n637), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n422), .A2(new_n596), .A3(new_n425), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n581), .A2(KEYINPUT44), .A3(new_n619), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n619), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n745), .B1(new_n746), .B2(new_n607), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n700), .A2(new_n702), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g564(.A(KEYINPUT104), .B(G137), .Z(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G39));
  NOR3_X1   g566(.A1(new_n671), .A2(new_n681), .A3(new_n711), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n748), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n739), .A2(new_n304), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n739), .A2(KEYINPUT47), .A3(new_n304), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n375), .ZN(G42));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n464), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n457), .A2(new_n463), .A3(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n588), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT107), .Z(new_n766));
  XOR2_X1   g580(.A(new_n597), .B(KEYINPUT105), .Z(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n582), .A2(new_n768), .A3(new_n373), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n620), .A2(new_n576), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n700), .A2(new_n702), .A3(new_n709), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n723), .A2(new_n633), .B1(new_n687), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n422), .A2(new_n764), .A3(new_n425), .A4(new_n628), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n619), .A2(new_n364), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n560), .B2(new_n571), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n748), .A3(new_n778), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n305), .B(new_n774), .C1(new_n351), .C2(new_n363), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n780), .B(new_n619), .C1(new_n625), .C2(new_n559), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n700), .A2(new_n702), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT108), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n773), .A2(new_n784), .A3(KEYINPUT109), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT109), .B1(new_n773), .B2(new_n784), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n771), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n665), .A2(new_n668), .A3(new_n684), .A4(new_n672), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n717), .A2(new_n791), .A3(KEYINPUT53), .A4(new_n720), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n635), .B1(new_n691), .B2(new_n693), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n709), .A2(new_n642), .A3(KEYINPUT110), .A4(new_n628), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  INV_X1    g609(.A(new_n363), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n304), .B(new_n628), .C1(new_n796), .C2(new_n707), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n797), .B2(new_n619), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n586), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n800), .B(new_n645), .C1(new_n560), .C2(new_n650), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n799), .A2(new_n801), .B1(new_n654), .B2(new_n656), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n793), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n793), .A2(KEYINPUT52), .A3(new_n802), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n792), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT111), .B(new_n771), .C1(new_n785), .C2(new_n786), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n789), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n716), .A2(new_n790), .A3(new_n719), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n811), .B(new_n771), .C1(new_n785), .C2(new_n786), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n793), .A2(KEYINPUT52), .A3(new_n802), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(new_n793), .B2(new_n802), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n810), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n817));
  NAND3_X1  g631(.A1(new_n809), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n773), .A2(new_n784), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n773), .A2(new_n784), .A3(KEYINPUT109), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n770), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n805), .A2(new_n806), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n826), .A3(KEYINPUT53), .A4(new_n811), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n816), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT54), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n809), .A2(KEYINPUT113), .A3(new_n816), .A4(new_n817), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n782), .A2(new_n366), .A3(new_n663), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n560), .A2(new_n650), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n681), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n588), .A2(new_n596), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n743), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n680), .A2(new_n619), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n833), .A2(new_n834), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n366), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n680), .A2(new_n681), .A3(new_n839), .A4(new_n743), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n664), .A2(new_n643), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n840), .A2(new_n641), .A3(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n840), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n757), .A2(new_n758), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n659), .B(new_n661), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(new_n305), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n748), .B(new_n846), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n845), .A2(KEYINPUT51), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT51), .B1(new_n845), .B2(new_n850), .ZN(new_n852));
  INV_X1    g666(.A(G952), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n853), .B(G953), .C1(new_n846), .C2(new_n690), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n831), .A2(new_n715), .A3(new_n743), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n856));
  INV_X1    g670(.A(new_n715), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n835), .A2(KEYINPUT48), .A3(new_n857), .ZN(new_n858));
  OAI221_X1 g672(.A(new_n854), .B1(new_n597), .B2(new_n833), .C1(new_n856), .C2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n851), .A2(new_n852), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n820), .A2(new_n829), .A3(new_n830), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT114), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n829), .A2(new_n830), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n864), .A3(new_n820), .A4(new_n860), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n853), .A2(new_n272), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n741), .A2(new_n305), .A3(new_n643), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT49), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n868), .B1(new_n848), .B2(new_n869), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n513), .B(new_n870), .C1(new_n869), .C2(new_n848), .ZN(new_n871));
  INV_X1    g685(.A(new_n641), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n832), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n867), .A2(new_n873), .ZN(G75));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n809), .A2(new_n816), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(G902), .ZN(new_n877));
  INV_X1    g691(.A(G210), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n246), .A2(new_n277), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(new_n275), .Z(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n881), .B(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n879), .A2(new_n883), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n272), .A2(G952), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G51));
  NAND2_X1  g701(.A1(new_n818), .A2(KEYINPUT116), .ZN(new_n888));
  INV_X1    g702(.A(new_n817), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n876), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n809), .A2(new_n891), .A3(new_n816), .A4(new_n817), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n350), .B(KEYINPUT57), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n360), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n734), .B(KEYINPUT117), .Z(new_n897));
  NAND3_X1  g711(.A1(new_n876), .A2(G902), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n886), .B1(new_n896), .B2(new_n898), .ZN(G54));
  NOR2_X1   g713(.A1(new_n410), .A2(new_n417), .ZN(new_n900));
  NAND2_X1  g714(.A1(KEYINPUT58), .A2(G475), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n877), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n886), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n877), .A2(new_n900), .A3(new_n901), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT118), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n877), .A2(new_n900), .A3(new_n901), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n907), .A2(new_n908), .A3(new_n903), .A4(new_n902), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n906), .A2(new_n909), .ZN(G60));
  AND2_X1   g724(.A1(new_n590), .A2(new_n591), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n593), .B(KEYINPUT59), .Z(new_n912));
  NAND3_X1  g726(.A1(new_n893), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n903), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n820), .A2(new_n829), .A3(new_n830), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n915), .B2(new_n912), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT60), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n876), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n492), .A2(new_n497), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT121), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT122), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n616), .A2(new_n617), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT120), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n903), .B1(new_n920), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n920), .A2(new_n931), .A3(new_n923), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n925), .A2(new_n930), .A3(KEYINPUT61), .A4(new_n932), .ZN(new_n933));
  XOR2_X1   g747(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n921), .A2(new_n924), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n929), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(G66));
  INV_X1    g751(.A(G224), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n367), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n770), .A2(new_n790), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n880), .B1(G898), .B2(new_n272), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G69));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n715), .A2(new_n588), .A3(new_n586), .A4(new_n644), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n724), .B1(new_n945), .B2(new_n740), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n721), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n750), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n759), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n793), .A2(new_n657), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n947), .A2(new_n949), .A3(new_n272), .A4(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n527), .B1(new_n535), .B2(new_n539), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(new_n415), .ZN(new_n953));
  NAND2_X1  g767(.A1(G900), .A2(G953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n944), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n638), .B1(new_n766), .B2(new_n767), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n572), .A3(new_n748), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n740), .B2(new_n749), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT123), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n958), .C1(new_n740), .C2(new_n749), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n759), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n635), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n694), .A2(new_n652), .A3(new_n964), .A4(new_n657), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n965), .A2(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(KEYINPUT62), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n963), .A2(new_n966), .A3(KEYINPUT124), .A4(new_n967), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n956), .B1(new_n972), .B2(new_n953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT125), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n956), .B(new_n975), .C1(new_n972), .C2(new_n953), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n974), .A2(new_n976), .A3(new_n978), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  INV_X1    g798(.A(new_n568), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n547), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n828), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n988));
  INV_X1    g802(.A(new_n940), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n540), .A3(new_n646), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n903), .B(new_n987), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n970), .A2(new_n940), .A3(new_n971), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n545), .B(new_n648), .C1(new_n996), .C2(new_n984), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n995), .A2(new_n997), .ZN(G57));
endmodule


