//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1122, new_n1123, new_n1125,
    new_n1126;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(new_n452));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G567), .B1(new_n454), .B2(G2106), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT69), .B(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(new_n460), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n462), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n470), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n469), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n469), .B2(G112), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n469), .B(new_n470), .C1(new_n466), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n482), .B1(new_n483), .B2(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n479), .A2(G138), .A3(new_n469), .A4(new_n470), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n472), .A2(new_n498), .A3(G138), .A4(new_n469), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n469), .A2(G102), .A3(G2104), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n480), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n502), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT6), .B(G651), .Z(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n516), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT74), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(G543), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n528), .A2(new_n529), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n534), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(new_n525), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n510), .A2(new_n512), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n539), .A2(G90), .B1(G651), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n538), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT75), .B(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n533), .A2(new_n547), .B1(new_n525), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n549), .B(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n515), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n534), .A2(KEYINPUT9), .A3(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n541), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n539), .A2(G91), .B1(G651), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n533), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n562), .A2(new_n566), .A3(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n534), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n539), .A2(G87), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n541), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT77), .Z(new_n579));
  AOI22_X1  g154(.A1(new_n513), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n518), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n515), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT78), .Z(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n533), .A2(new_n586), .B1(new_n587), .B2(new_n525), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n588), .A2(KEYINPUT79), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(KEYINPUT79), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n585), .B1(new_n589), .B2(new_n590), .ZN(G290));
  AOI22_X1  g166(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n515), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(G54), .B2(new_n534), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n513), .A2(G92), .A3(new_n524), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT80), .B1(new_n598), .B2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  MUX2_X1   g175(.A(KEYINPUT80), .B(new_n599), .S(new_n600), .Z(G284));
  MUX2_X1   g176(.A(KEYINPUT80), .B(new_n599), .S(new_n600), .Z(G321));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT81), .B1(new_n603), .B2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  MUX2_X1   g180(.A(KEYINPUT81), .B(new_n604), .S(new_n605), .Z(G297));
  MUX2_X1   g181(.A(KEYINPUT81), .B(new_n604), .S(new_n605), .Z(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n598), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n598), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n555), .B2(G868), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND3_X1   g188(.A1(new_n472), .A2(new_n469), .A3(new_n466), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n481), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(new_n469), .B2(G111), .ZN(new_n620));
  INV_X1    g195(.A(G135), .ZN(new_n621));
  OAI221_X1 g196(.A(new_n618), .B1(new_n619), .B2(new_n620), .C1(new_n488), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n617), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT83), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2451), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT84), .Z(new_n639));
  INV_X1    g214(.A(G14), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n636), .B2(new_n637), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT17), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XOR2_X1   g221(.A(G2067), .B(G2678), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT85), .ZN(new_n649));
  INV_X1    g224(.A(new_n646), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n644), .A2(new_n647), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n650), .B(new_n651), .C1(new_n645), .C2(new_n647), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n650), .A2(new_n644), .A3(new_n647), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n661), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT87), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT22), .B(G1981), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G27), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G164), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2078), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT28), .ZN(new_n685));
  INV_X1    g260(.A(G26), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(G29), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(G29), .ZN(new_n688));
  INV_X1    g263(.A(new_n488), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n689), .A2(G140), .B1(G128), .B2(new_n481), .ZN(new_n690));
  NOR2_X1   g265(.A1(G104), .A2(G2105), .ZN(new_n691));
  OAI21_X1  g266(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n688), .B1(new_n693), .B2(G29), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n687), .B1(new_n694), .B2(new_n685), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G2067), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G19), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n555), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT89), .B(G1341), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(G29), .A2(G33), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT25), .Z(new_n704));
  AOI22_X1  g279(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n705));
  INV_X1    g280(.A(G139), .ZN(new_n706));
  OAI221_X1 g281(.A(new_n704), .B1(new_n469), .B2(new_n705), .C1(new_n488), .C2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n702), .B1(new_n707), .B2(new_n681), .ZN(new_n708));
  INV_X1    g283(.A(G2072), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n695), .A2(G2067), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n696), .A2(new_n701), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n681), .A2(G35), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n681), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT29), .Z(new_n715));
  INV_X1    g290(.A(G2090), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(KEYINPUT24), .A2(G34), .ZN(new_n718));
  NAND2_X1  g293(.A1(KEYINPUT24), .A2(G34), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n681), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G160), .B2(new_n681), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2084), .ZN(new_n722));
  OR4_X1    g297(.A1(new_n684), .A2(new_n712), .A3(new_n717), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n697), .A2(G5), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G171), .B2(new_n697), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT93), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n598), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G4), .B2(G16), .ZN(new_n729));
  INV_X1    g304(.A(G1348), .ZN(new_n730));
  OAI22_X1  g305(.A1(new_n726), .A2(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G168), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G16), .B2(G21), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n681), .B2(new_n622), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n731), .B(new_n736), .C1(new_n715), .C2(new_n716), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n726), .A2(new_n727), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n681), .A2(G32), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n689), .A2(G141), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n481), .A2(G129), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n466), .A2(G105), .A3(new_n469), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT91), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT26), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n740), .A2(new_n741), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n681), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n737), .A2(new_n738), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT23), .ZN(new_n754));
  INV_X1    g329(.A(G20), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G16), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n753), .B(new_n756), .C1(new_n603), .C2(new_n697), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1956), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n729), .A2(new_n730), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT30), .B(G28), .Z(new_n760));
  OAI221_X1 g335(.A(new_n759), .B1(G29), .B2(new_n760), .C1(new_n733), .C2(new_n734), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n723), .A2(new_n752), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n697), .A2(G23), .ZN(new_n763));
  INV_X1    g338(.A(G288), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n697), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT33), .ZN(new_n766));
  INV_X1    g341(.A(G1976), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  MUX2_X1   g344(.A(G6), .B(G305), .S(G16), .Z(new_n770));
  XOR2_X1   g345(.A(KEYINPUT32), .B(G1981), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n697), .A2(G22), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n697), .ZN(new_n774));
  INV_X1    g349(.A(G1971), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n768), .A2(new_n769), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT34), .ZN(new_n778));
  NOR2_X1   g353(.A1(G16), .A2(G24), .ZN(new_n779));
  XNOR2_X1  g354(.A(G290), .B(KEYINPUT88), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(G16), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G1986), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n777), .A2(KEYINPUT34), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n689), .A2(G131), .B1(G119), .B2(new_n481), .ZN(new_n784));
  NOR2_X1   g359(.A1(G95), .A2(G2105), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(new_n469), .B2(G107), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G25), .B(new_n787), .S(G29), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT35), .B(G1991), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n788), .B(new_n789), .Z(new_n790));
  NAND4_X1  g365(.A1(new_n778), .A2(new_n782), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT36), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n708), .A2(new_n709), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT90), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT31), .B(G11), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n762), .A2(new_n792), .A3(new_n794), .A4(new_n795), .ZN(G150));
  INV_X1    g371(.A(G150), .ZN(G311));
  AOI22_X1  g372(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(new_n515), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT95), .Z(new_n800));
  INV_X1    g375(.A(G55), .ZN(new_n801));
  INV_X1    g376(.A(G93), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n533), .A2(new_n801), .B1(new_n802), .B2(new_n525), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G860), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT37), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n554), .B(new_n804), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n597), .A2(new_n608), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT39), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n808), .B(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(G860), .ZN(G145));
  XNOR2_X1  g389(.A(new_n693), .B(new_n507), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(new_n707), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(new_n747), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n481), .A2(G130), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n469), .A2(G118), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT96), .Z(new_n821));
  INV_X1    g396(.A(G142), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n818), .B1(new_n819), .B2(new_n821), .C1(new_n488), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n615), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n787), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT97), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n817), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n622), .B(G160), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G162), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G37), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n829), .B1(new_n817), .B2(new_n826), .ZN(new_n832));
  INV_X1    g407(.A(new_n825), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n817), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n837));
  INV_X1    g412(.A(G868), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n808), .B(new_n610), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n597), .B(G299), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n840), .A2(KEYINPUT41), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT98), .B1(new_n840), .B2(KEYINPUT41), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n842), .B(new_n843), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n839), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(G290), .B(G305), .ZN(new_n849));
  XNOR2_X1  g424(.A(G288), .B(G303), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT99), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n841), .A2(KEYINPUT100), .A3(new_n845), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n853), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n848), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n846), .ZN(new_n859));
  INV_X1    g434(.A(new_n857), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n859), .B(KEYINPUT100), .C1(new_n860), .C2(new_n854), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n838), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n805), .A2(G868), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n837), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n862), .A2(KEYINPUT101), .A3(new_n864), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(G295));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n863), .B2(new_n865), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n862), .A2(KEYINPUT102), .A3(new_n864), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(G331));
  XNOR2_X1  g447(.A(G286), .B(G171), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n808), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(new_n840), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n840), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n840), .A2(KEYINPUT41), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n842), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n851), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n844), .A2(new_n874), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n875), .A2(new_n851), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n831), .A3(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT106), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(KEYINPUT106), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(KEYINPUT43), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n875), .A2(new_n884), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n882), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n831), .A3(new_n885), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n892), .A2(KEYINPUT43), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(KEYINPUT44), .A3(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n895));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n883), .A2(new_n896), .A3(new_n831), .A4(new_n885), .ZN(new_n897));
  AOI22_X1  g472(.A1(KEYINPUT104), .A2(new_n897), .B1(new_n892), .B2(KEYINPUT43), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n892), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n900), .ZN(G397));
  AOI21_X1  g476(.A(G1384), .B1(new_n500), .B2(new_n506), .ZN(new_n902));
  XNOR2_X1  g477(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(G160), .A2(G40), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT109), .ZN(new_n907));
  INV_X1    g482(.A(G2067), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n693), .B(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G1996), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(new_n747), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n906), .A2(G1996), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n907), .A2(new_n911), .B1(new_n747), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n787), .A2(new_n789), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n787), .A2(new_n789), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n907), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n906), .ZN(new_n919));
  OR2_X1    g494(.A1(G290), .A2(G1986), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT108), .ZN(new_n921));
  NAND2_X1  g496(.A1(G290), .A2(G1986), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n918), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT114), .ZN(new_n925));
  NAND2_X1  g500(.A1(G160), .A2(G40), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n902), .B2(new_n903), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n496), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT71), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n930));
  AND4_X1   g505(.A1(G138), .A2(new_n472), .A3(new_n498), .A4(new_n469), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n506), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n925), .B1(new_n937), .B2(new_n734), .ZN(new_n938));
  AOI211_X1 g513(.A(KEYINPUT114), .B(G1966), .C1(new_n927), .C2(new_n936), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n902), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n926), .B1(new_n941), .B2(KEYINPUT111), .ZN(new_n942));
  AOI211_X1 g517(.A(KEYINPUT50), .B(G1384), .C1(new_n500), .C2(new_n506), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n934), .A2(KEYINPUT50), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n938), .A2(new_n939), .B1(new_n947), .B2(G2084), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI221_X1 g525(.A(KEYINPUT122), .B1(new_n947), .B2(G2084), .C1(new_n938), .C2(new_n939), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(G168), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G8), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT51), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(KEYINPUT51), .A3(new_n951), .ZN(new_n955));
  INV_X1    g530(.A(new_n948), .ZN(new_n956));
  OAI21_X1  g531(.A(G168), .B1(new_n956), .B2(KEYINPUT51), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n957), .A3(G8), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G303), .A2(G8), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT55), .Z(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT112), .Z(new_n962));
  AOI21_X1  g537(.A(new_n926), .B1(new_n902), .B2(KEYINPUT45), .ZN(new_n963));
  INV_X1    g538(.A(new_n903), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n934), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n963), .A2(new_n965), .A3(KEYINPUT110), .ZN(new_n969));
  AOI21_X1  g544(.A(G1971), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n947), .A2(G2090), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n962), .B(G8), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G8), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n905), .B2(new_n902), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n764), .A2(G1976), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n976), .B(new_n977), .C1(G1976), .C2(new_n764), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n581), .A2(new_n578), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G1981), .ZN(new_n981));
  OAI221_X1 g556(.A(new_n981), .B1(KEYINPUT113), .B2(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n982));
  NAND2_X1  g557(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(G305), .A2(G1981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n981), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n984), .B(new_n974), .C1(new_n983), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n978), .A2(new_n979), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n969), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT110), .B1(new_n963), .B2(new_n965), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n775), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n940), .B1(new_n507), .B2(new_n928), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n993), .A2(new_n943), .A3(new_n926), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n716), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n973), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n972), .B(new_n989), .C1(new_n996), .C2(new_n961), .ZN(new_n997));
  INV_X1    g572(.A(new_n947), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(G1961), .ZN(new_n999));
  XNOR2_X1  g574(.A(G301), .B(KEYINPUT54), .ZN(new_n1000));
  INV_X1    g575(.A(G2078), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n968), .A2(new_n1001), .A3(new_n969), .ZN(new_n1002));
  NAND2_X1  g577(.A1(KEYINPUT123), .A2(KEYINPUT53), .ZN(new_n1003));
  OR2_X1    g578(.A1(KEYINPUT123), .A2(KEYINPUT53), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT124), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1002), .A2(KEYINPUT124), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n999), .B(new_n1000), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n963), .A2(new_n965), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT125), .B(G2078), .Z(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n997), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n999), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n927), .A2(new_n936), .A3(KEYINPUT53), .A4(new_n1001), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1000), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n959), .A2(new_n1013), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n905), .A2(new_n902), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT58), .B(G1341), .Z(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n966), .B2(G1996), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n555), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1022), .B2(new_n555), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT56), .B(G2072), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n963), .A2(new_n965), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(G299), .B(KEYINPUT57), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1028), .B(new_n1030), .C1(new_n994), .C2(G1956), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n946), .A2(new_n905), .A3(new_n941), .ZN(new_n1034));
  INV_X1    g609(.A(G1956), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1010), .A2(new_n1027), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1029), .B(KEYINPUT116), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1033), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1028), .B1(new_n994), .B2(G1956), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1029), .B(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1041), .A3(KEYINPUT117), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1032), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1026), .B1(new_n1043), .B2(KEYINPUT61), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n993), .A2(new_n943), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1956), .B1(new_n1047), .B2(new_n905), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n963), .A2(new_n965), .A3(new_n1027), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1046), .B(new_n1029), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1031), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1046), .B1(new_n1039), .B2(new_n1029), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1045), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT119), .B(new_n1045), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1044), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1044), .A2(new_n1055), .A3(KEYINPUT120), .A4(new_n1056), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1019), .A2(G2067), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n947), .B2(new_n730), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n598), .B1(new_n1062), .B2(KEYINPUT60), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1062), .A2(KEYINPUT60), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT121), .B(new_n598), .C1(new_n1062), .C2(KEYINPUT60), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1059), .A2(new_n1060), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n597), .B2(new_n1062), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1031), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1018), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n955), .A2(new_n957), .A3(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n952), .B2(G8), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT62), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n954), .A2(new_n1080), .A3(new_n958), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1015), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n999), .B(new_n1082), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1083), .A2(new_n997), .A3(G301), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n987), .A2(new_n767), .A3(new_n764), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n985), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n974), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n972), .B2(new_n988), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  OAI21_X1  g665(.A(G8), .B1(new_n970), .B2(new_n971), .ZN(new_n1091));
  INV_X1    g666(.A(new_n961), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n988), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n1093), .B2(KEYINPUT115), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n998), .A2(new_n716), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n973), .B1(new_n1095), .B2(new_n992), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n989), .B1(new_n1096), .B2(new_n961), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n956), .A2(new_n973), .A3(G286), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1094), .A2(new_n1099), .A3(new_n972), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1100), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1090), .B1(new_n1102), .B2(new_n997), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1089), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1085), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n924), .B1(new_n1075), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n920), .A2(new_n906), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT48), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n918), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n909), .A2(new_n747), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n907), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT127), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n912), .B(KEYINPUT46), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT47), .Z(new_n1115));
  NOR2_X1   g690(.A1(new_n693), .A2(G2067), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n913), .B2(new_n914), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT126), .Z(new_n1118));
  AOI211_X1 g693(.A(new_n1109), .B(new_n1115), .C1(new_n907), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1106), .A2(new_n1119), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g695(.A(new_n835), .B(new_n457), .C1(new_n898), .C2(new_n899), .ZN(new_n1122));
  NAND3_X1  g696(.A1(new_n642), .A2(new_n657), .A3(new_n679), .ZN(new_n1123));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n1123), .ZN(G308));
  OR2_X1    g698(.A1(new_n898), .A2(new_n899), .ZN(new_n1125));
  INV_X1    g699(.A(new_n1123), .ZN(new_n1126));
  NAND4_X1  g700(.A1(new_n1125), .A2(new_n457), .A3(new_n835), .A4(new_n1126), .ZN(G225));
endmodule


