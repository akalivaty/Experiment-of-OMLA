//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n193), .A3(new_n196), .A4(new_n191), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT76), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(KEYINPUT76), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n199), .A2(new_n202), .A3(KEYINPUT76), .A4(G104), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n205), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n207), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G101), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT1), .B1(new_n215), .B2(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(G128), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n214), .B(new_n216), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n219), .A2(new_n221), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n209), .A3(new_n211), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n198), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n226), .B(KEYINPUT12), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n209), .A2(KEYINPUT10), .A3(new_n211), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n219), .A2(KEYINPUT66), .A3(new_n221), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n233));
  AOI22_X1  g047(.A1(new_n228), .A2(new_n232), .B1(new_n225), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT76), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n206), .A2(G107), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n208), .A2(new_n207), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n235), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n204), .A2(KEYINPUT77), .A3(new_n207), .A4(new_n208), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(G101), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n240), .A2(new_n241), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(new_n205), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n214), .A2(new_n216), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G143), .B(G146), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n242), .A2(new_n243), .A3(G101), .A4(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n248), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n234), .A2(new_n257), .A3(new_n198), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n227), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G140), .ZN(new_n260));
  INV_X1    g074(.A(G227), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G953), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n260), .B(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n198), .B1(new_n234), .B2(new_n257), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G469), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n187), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n258), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n263), .B1(new_n272), .B2(new_n267), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n227), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT81), .B1(new_n258), .B2(new_n265), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n273), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n270), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n265), .B1(new_n227), .B2(new_n258), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n266), .A2(new_n267), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT80), .A3(G469), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n271), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT9), .B(G234), .ZN(new_n285));
  OAI21_X1  g099(.A(G221), .B1(new_n285), .B2(G902), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G214), .B1(G237), .B2(G902), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n288), .B(KEYINPUT82), .Z(new_n289));
  OAI21_X1  g103(.A(G210), .B1(G237), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n254), .A2(G125), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(G125), .B2(new_n222), .ZN(new_n293));
  INV_X1    g107(.A(G224), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(G953), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT86), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n293), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G110), .B(G122), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n301));
  XNOR2_X1  g115(.A(G116), .B(G119), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT2), .B(G113), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n304), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n302), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n248), .A2(new_n301), .A3(new_n308), .A4(new_n256), .ZN(new_n309));
  INV_X1    g123(.A(new_n212), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n302), .A2(KEYINPUT5), .ZN(new_n311));
  INV_X1    g125(.A(G116), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n312), .A2(KEYINPUT5), .A3(G119), .ZN(new_n313));
  INV_X1    g127(.A(G113), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n311), .A2(new_n315), .B1(new_n306), .B2(new_n302), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n309), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n308), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n244), .B2(new_n247), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n301), .B1(new_n320), .B2(new_n256), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT85), .B(new_n300), .C1(new_n318), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT6), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n248), .A2(new_n308), .A3(new_n256), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT83), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(new_n317), .A3(new_n309), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n327), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n300), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT84), .B1(new_n327), .B2(new_n300), .ZN(new_n330));
  INV_X1    g144(.A(new_n318), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT84), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n299), .A4(new_n326), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n300), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n298), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n333), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT7), .B1(new_n294), .B2(G953), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n293), .B(new_n338), .Z(new_n339));
  NOR2_X1   g153(.A1(new_n310), .A2(new_n316), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n311), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n302), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n315), .A3(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n310), .A2(new_n344), .A3(new_n307), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n340), .B1(new_n345), .B2(KEYINPUT88), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(KEYINPUT88), .B2(new_n345), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n299), .B(KEYINPUT8), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n339), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n337), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n278), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n291), .B1(new_n336), .B2(new_n351), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n330), .A2(new_n334), .A3(new_n333), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n324), .A2(new_n328), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n297), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(G902), .B1(new_n337), .B2(new_n349), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n290), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n289), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n215), .A2(G128), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n220), .A2(G143), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(new_n189), .ZN(new_n362));
  XNOR2_X1  g176(.A(G116), .B(G122), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n202), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n312), .A2(KEYINPUT14), .A3(G122), .ZN(new_n365));
  INV_X1    g179(.A(new_n363), .ZN(new_n366));
  OAI211_X1 g180(.A(G107), .B(new_n365), .C1(new_n366), .C2(KEYINPUT14), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n359), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n369), .A2(KEYINPUT13), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n360), .B1(new_n369), .B2(KEYINPUT13), .ZN(new_n371));
  OAI21_X1  g185(.A(G134), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n361), .A2(new_n189), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n363), .B(new_n202), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G217), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n285), .A2(new_n377), .A3(G953), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n368), .A2(new_n375), .A3(new_n378), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n278), .ZN(new_n384));
  INV_X1    g198(.A(G478), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT91), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT15), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(KEYINPUT15), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n384), .B(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G125), .B(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT16), .ZN(new_n393));
  INV_X1    g207(.A(G125), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n394), .A2(KEYINPUT16), .A3(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n213), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(G146), .A3(new_n395), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  INV_X1    g214(.A(G953), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(G214), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n215), .ZN(new_n403));
  NOR2_X1   g217(.A1(G237), .A2(G953), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(G143), .A3(G214), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT17), .A3(G131), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(G131), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n399), .B(new_n407), .C1(KEYINPUT17), .C2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G113), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n206), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n392), .A2(new_n213), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n392), .A2(new_n213), .ZN(new_n413));
  AND2_X1   g227(.A1(KEYINPUT18), .A2(G131), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n412), .A2(new_n413), .B1(new_n406), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n406), .A2(new_n414), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n416), .A2(KEYINPUT89), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(KEYINPUT89), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n409), .A2(new_n411), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n411), .B1(new_n409), .B2(new_n419), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n278), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G475), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n392), .B(KEYINPUT19), .Z(new_n425));
  OAI211_X1 g239(.A(new_n408), .B(new_n398), .C1(G146), .C2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n420), .B1(new_n427), .B2(new_n411), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n429));
  NOR2_X1   g243(.A1(G475), .A2(G902), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n429), .B1(new_n428), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n424), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n401), .A2(G952), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(G234), .B2(G237), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n278), .B(new_n401), .C1(G234), .C2(G237), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(G898), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n391), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n287), .A2(new_n358), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(G217), .A2(G902), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n377), .B2(G234), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n443), .B(KEYINPUT70), .Z(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT71), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n401), .A2(G221), .A3(G234), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT74), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT22), .B(G137), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT23), .ZN(new_n454));
  INV_X1    g268(.A(G119), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(G128), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(G128), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n220), .A2(KEYINPUT23), .A3(G119), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G110), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT72), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n220), .B2(G119), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(KEYINPUT72), .A3(G128), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n463), .B(new_n464), .C1(new_n455), .C2(G128), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT24), .B(G110), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT73), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n398), .A2(new_n413), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n397), .A2(new_n398), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n465), .A2(new_n466), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n459), .A2(new_n460), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n453), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n468), .B(KEYINPUT73), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n398), .A3(new_n413), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n476), .A3(new_n452), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n448), .B1(new_n482), .B2(new_n278), .ZN(new_n483));
  AOI211_X1 g297(.A(G902), .B(new_n447), .C1(new_n478), .C2(new_n481), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n446), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n444), .A2(new_n278), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n404), .A2(G210), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT27), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT26), .B(G101), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n253), .A2(KEYINPUT64), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n195), .A2(new_n197), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n250), .B(new_n496), .C1(new_n251), .C2(new_n252), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT65), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT65), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n494), .A2(new_n495), .A3(new_n500), .A4(new_n497), .ZN(new_n501));
  INV_X1    g315(.A(new_n191), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n189), .A2(G137), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n197), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n224), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n499), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n308), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n505), .B1(new_n230), .B2(new_n231), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n495), .A2(new_n254), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n319), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n493), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n219), .A2(KEYINPUT66), .A3(new_n221), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT66), .B1(new_n219), .B2(new_n221), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n506), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n511), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n308), .B1(new_n519), .B2(KEYINPUT68), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n521), .A3(new_n511), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT28), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n492), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n508), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n513), .A2(KEYINPUT30), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n308), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n492), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n514), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT29), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT68), .B1(new_n510), .B2(new_n512), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n319), .A3(new_n522), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n493), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n519), .A2(new_n308), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n319), .B1(new_n518), .B2(new_n511), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT28), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n492), .A2(KEYINPUT29), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n278), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G472), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT69), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT69), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n543), .B(G472), .C1(new_n531), .C2(new_n540), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n535), .A2(new_n529), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n546), .B1(new_n528), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n498), .A2(KEYINPUT65), .B1(new_n506), .B2(new_n224), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n319), .B1(new_n549), .B2(new_n501), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT28), .B1(new_n550), .B2(new_n535), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n492), .B1(new_n551), .B2(new_n534), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n528), .A2(new_n546), .A3(new_n547), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT67), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n528), .A2(KEYINPUT67), .A3(new_n546), .A4(new_n547), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n548), .B(new_n552), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(G472), .A2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT32), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n556), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n552), .A2(new_n548), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT32), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n558), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n488), .B1(new_n545), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n441), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT92), .B(G101), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(G3));
  NAND2_X1  g384(.A1(new_n352), .A2(new_n357), .ZN(new_n571));
  INV_X1    g385(.A(new_n289), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n383), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n379), .A2(KEYINPUT33), .A3(new_n380), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n385), .A2(G902), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n384), .A2(new_n385), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n434), .A2(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n573), .A2(new_n439), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G472), .B1(new_n557), .B2(G902), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n559), .B2(new_n557), .ZN(new_n584));
  INV_X1    g398(.A(new_n488), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n284), .A3(new_n286), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT34), .B(G104), .Z(new_n589));
  XOR2_X1   g403(.A(new_n589), .B(KEYINPUT93), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n588), .B(new_n590), .ZN(G6));
  INV_X1    g405(.A(new_n434), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n391), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n573), .A2(new_n439), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n587), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT94), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G107), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  NAND2_X1  g412(.A1(new_n480), .A2(new_n476), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n278), .A3(new_n444), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n485), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n584), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n441), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT37), .B(G110), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT95), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n605), .B(new_n607), .ZN(G12));
  AOI211_X1 g422(.A(new_n289), .B(new_n603), .C1(new_n352), .C2(new_n357), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n564), .B1(new_n563), .B2(new_n558), .ZN(new_n610));
  AOI211_X1 g424(.A(KEYINPUT32), .B(new_n559), .C1(new_n561), .C2(new_n562), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n544), .B(new_n542), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G900), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n436), .B1(new_n437), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n593), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n609), .A2(new_n612), .A3(new_n287), .A4(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT96), .B(G128), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G30));
  XOR2_X1   g432(.A(new_n614), .B(KEYINPUT39), .Z(new_n619));
  NAND2_X1  g433(.A1(new_n287), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT99), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n571), .B(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n535), .A2(new_n536), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n278), .B1(new_n628), .B2(new_n492), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n529), .B1(new_n528), .B2(new_n514), .ZN(new_n630));
  OAI21_X1  g444(.A(G472), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT98), .B1(new_n566), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(KEYINPUT98), .B(new_n631), .C1(new_n610), .C2(new_n611), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n391), .A2(new_n434), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n603), .A2(new_n636), .A3(new_n572), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n623), .A2(new_n626), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n215), .ZN(G45));
  INV_X1    g454(.A(new_n614), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n434), .A2(new_n580), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n609), .A2(new_n612), .A3(new_n287), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G146), .ZN(G48));
  NAND2_X1  g459(.A1(new_n612), .A2(new_n585), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n277), .A2(new_n270), .A3(new_n278), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n648));
  INV_X1    g462(.A(new_n286), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n582), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT41), .B(G113), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G15));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n594), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G116), .ZN(G18));
  AND3_X1   g471(.A1(new_n612), .A2(new_n440), .A3(new_n650), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n609), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G119), .ZN(G21));
  AOI21_X1  g474(.A(new_n492), .B1(new_n534), .B2(new_n537), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n548), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n514), .A2(new_n492), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n510), .A2(new_n512), .A3(new_n525), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n525), .B2(new_n508), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n663), .B1(new_n665), .B2(new_n308), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT67), .B1(new_n666), .B2(new_n546), .ZN(new_n667));
  INV_X1    g481(.A(new_n556), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n558), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n585), .A2(new_n583), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n439), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n650), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n571), .A2(new_n572), .A3(new_n636), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G122), .ZN(G24));
  NAND2_X1  g491(.A1(new_n485), .A2(new_n602), .ZN(new_n678));
  INV_X1    g492(.A(G472), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n561), .B2(new_n562), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n670), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n583), .A2(KEYINPUT100), .A3(new_n678), .A4(new_n670), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n336), .A2(new_n351), .A3(new_n291), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n290), .B1(new_n355), .B2(new_n356), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n650), .B(new_n572), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n428), .A2(new_n430), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n431), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n692), .A2(new_n424), .B1(new_n578), .B2(new_n579), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(KEYINPUT101), .A3(new_n641), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n642), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n685), .A2(new_n689), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  NAND2_X1  g513(.A1(new_n282), .A2(G469), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n649), .B1(new_n279), .B2(new_n700), .ZN(new_n701));
  AND4_X1   g515(.A1(new_n572), .A2(new_n352), .A3(new_n357), .A4(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n612), .A3(new_n585), .A4(new_n697), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n567), .A2(KEYINPUT42), .A3(new_n697), .A4(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G131), .ZN(G33));
  NAND4_X1  g522(.A1(new_n702), .A2(new_n612), .A3(new_n585), .A4(new_n615), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G134), .ZN(G36));
  XNOR2_X1  g524(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n592), .B2(new_n580), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n434), .B1(new_n579), .B2(new_n578), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(KEYINPUT43), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT104), .B1(new_n714), .B2(new_n711), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n584), .A3(new_n678), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT105), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n264), .A2(new_n268), .A3(KEYINPUT45), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT102), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT45), .B1(new_n264), .B2(new_n268), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n270), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n270), .A2(new_n278), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n722), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n279), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n728), .A2(new_n722), .A3(new_n729), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n286), .B(new_n619), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n352), .A2(new_n357), .A3(new_n572), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n718), .B2(new_n719), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n721), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G137), .ZN(G39));
  OAI21_X1  g552(.A(new_n286), .B1(new_n731), .B2(new_n732), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(KEYINPUT106), .B2(KEYINPUT47), .ZN(new_n740));
  AND2_X1   g554(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n741));
  NOR2_X1   g555(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n742));
  OAI221_X1 g556(.A(new_n286), .B1(new_n741), .B2(new_n742), .C1(new_n731), .C2(new_n732), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n612), .A2(new_n735), .A3(new_n585), .A4(new_n642), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G140), .ZN(G42));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n694), .A2(new_n696), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n683), .B2(new_n684), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT107), .A3(new_n702), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n685), .A2(new_n697), .A3(new_n702), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n735), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n603), .A2(new_n391), .A3(new_n434), .A4(new_n614), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n612), .A4(new_n287), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n709), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n707), .A2(new_n750), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n652), .B1(new_n582), .B2(new_n594), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n441), .B1(new_n567), .B2(new_n604), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n658), .A2(new_n609), .B1(new_n675), .B2(new_n674), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n573), .A2(new_n439), .ZN(new_n762));
  INV_X1    g576(.A(new_n593), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n762), .B(new_n587), .C1(new_n693), .C2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n603), .A2(new_n701), .A3(new_n641), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n675), .B(new_n768), .C1(new_n632), .C2(new_n634), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n698), .A3(new_n616), .A4(new_n644), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(KEYINPUT108), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n631), .B1(new_n610), .B2(new_n611), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT98), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n767), .B1(new_n776), .B2(new_n633), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n612), .A2(new_n287), .A3(new_n643), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n777), .A2(new_n675), .B1(new_n778), .B2(new_n609), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n612), .A2(new_n287), .A3(new_n615), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n609), .A2(new_n780), .B1(new_n749), .B2(new_n689), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n747), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n770), .A2(KEYINPUT108), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n782), .B1(new_n779), .B2(new_n781), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n773), .A2(new_n783), .A3(KEYINPUT52), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(KEYINPUT53), .A3(new_n766), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n785), .A2(KEYINPUT109), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(KEYINPUT109), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(KEYINPUT54), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  INV_X1    g609(.A(new_n436), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n715), .B2(new_n716), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n735), .A2(new_n651), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(KEYINPUT112), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n685), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n488), .A2(new_n796), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n635), .A2(new_n798), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n592), .A3(new_n579), .A4(new_n578), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n647), .A2(new_n648), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n286), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n740), .B2(new_n743), .ZN(new_n812));
  INV_X1    g626(.A(new_n671), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n797), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n735), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT110), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n804), .B(new_n808), .C1(new_n812), .C2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n626), .A2(new_n289), .A3(new_n650), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n814), .B1(new_n818), .B2(KEYINPUT111), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n626), .A2(new_n289), .A3(new_n650), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(KEYINPUT50), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n824));
  INV_X1    g638(.A(new_n822), .ZN(new_n825));
  INV_X1    g639(.A(new_n814), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n820), .B2(new_n821), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n824), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n795), .B1(new_n817), .B2(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n812), .A2(new_n816), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n823), .A2(new_n828), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n808), .A2(new_n804), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(KEYINPUT51), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n435), .B1(new_n826), .B2(new_n689), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n581), .B2(new_n806), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT113), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n835), .B(new_n838), .C1(new_n581), .C2(new_n806), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n803), .A2(new_n567), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT48), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT48), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n830), .A2(new_n834), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n766), .A2(new_n790), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n747), .B1(new_n849), .B2(new_n784), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n789), .A2(KEYINPUT53), .A3(new_n766), .A4(new_n771), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n794), .A2(new_n848), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(G952), .A2(G953), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT115), .Z(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n585), .A2(new_n714), .A3(new_n572), .A4(new_n286), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n635), .A3(new_n626), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT116), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n857), .A2(new_n865), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(G75));
  NOR2_X1   g681(.A1(new_n401), .A2(G952), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n278), .B1(new_n850), .B2(new_n852), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n870), .B2(G210), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n353), .A2(new_n354), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n298), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n355), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT55), .Z(new_n875));
  OAI21_X1  g689(.A(new_n869), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n850), .A2(new_n852), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT117), .B1(new_n877), .B2(G902), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n879), .B(new_n278), .C1(new_n850), .C2(new_n852), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n291), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n875), .B(KEYINPUT118), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n876), .B1(new_n882), .B2(new_n884), .ZN(G51));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n881), .B2(new_n728), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT120), .A4(new_n727), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n853), .A2(KEYINPUT119), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n853), .A2(KEYINPUT119), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n729), .B(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n277), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n868), .B1(new_n889), .B2(new_n896), .ZN(G54));
  AND2_X1   g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n881), .A2(new_n428), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n428), .B1(new_n881), .B2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n868), .ZN(G60));
  AND2_X1   g715(.A1(new_n575), .A2(new_n576), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n385), .A2(new_n278), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n893), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n794), .A2(new_n853), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n902), .B1(new_n907), .B2(new_n905), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n868), .A3(new_n908), .ZN(G63));
  XOR2_X1   g723(.A(new_n442), .B(KEYINPUT60), .Z(new_n910));
  NAND3_X1  g724(.A1(new_n877), .A2(new_n601), .A3(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n877), .A2(new_n910), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n869), .B(new_n911), .C1(new_n912), .C2(new_n482), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g728(.A1(new_n765), .A2(new_n401), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n438), .B2(new_n294), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(KEYINPUT122), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(KEYINPUT122), .B2(new_n915), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n872), .B1(G898), .B2(new_n401), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n918), .B(new_n919), .Z(G69));
  NAND3_X1  g734(.A1(new_n734), .A2(new_n567), .A3(new_n675), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n921), .A2(new_n709), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n781), .A2(new_n644), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n705), .B2(new_n706), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n922), .A2(new_n737), .A3(new_n745), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n401), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n613), .A2(G953), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n665), .B(KEYINPUT123), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(new_n425), .Z(new_n931));
  OR2_X1    g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(KEYINPUT124), .ZN(new_n933));
  OR3_X1    g747(.A1(new_n639), .A2(KEYINPUT62), .A3(new_n923), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT62), .B1(new_n639), .B2(new_n923), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n763), .A2(new_n693), .ZN(new_n936));
  OR4_X1    g750(.A1(new_n646), .A2(new_n620), .A3(new_n735), .A4(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n737), .A2(new_n745), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n939), .B2(G953), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n261), .B2(new_n613), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G72));
  NAND2_X1  g758(.A1(G472), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT63), .Z(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n925), .B2(new_n765), .ZN(new_n947));
  INV_X1    g761(.A(new_n530), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n946), .B1(new_n950), .B2(new_n765), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n951), .A2(KEYINPUT126), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n630), .B1(new_n951), .B2(KEYINPUT126), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n946), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n948), .A2(new_n630), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT127), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n792), .A2(new_n793), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n954), .A2(new_n958), .ZN(G57));
endmodule


