//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g024(.A(G2106), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT64), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n450), .B1(new_n458), .B2(new_n455), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(G137), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  XNOR2_X1  g057(.A(KEYINPUT66), .B(KEYINPUT4), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n462), .A2(new_n483), .A3(G138), .A4(new_n461), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n461), .ZN(new_n485));
  OR2_X1    g060(.A1(KEYINPUT66), .A2(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n471), .A2(new_n473), .A3(G126), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n461), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n470), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G102), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n499), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT69), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  INV_X1    g095(.A(new_n507), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(new_n520), .A3(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  XOR2_X1   g100(.A(KEYINPUT70), .B(KEYINPUT7), .Z(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n518), .A2(new_n521), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n519), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n518), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n529), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n516), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n507), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n522), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n519), .A2(G43), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n550), .A2(G860), .A3(new_n551), .A4(new_n552), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND4_X1  g133(.A1(new_n515), .A2(G53), .A3(G543), .A4(new_n517), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n518), .A2(G91), .A3(new_n521), .ZN(new_n564));
  XNOR2_X1  g139(.A(KEYINPUT73), .B(G65), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n521), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n516), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g143(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  OAI21_X1  g146(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n572));
  INV_X1    g147(.A(G49), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI221_X1 g149(.A(new_n572), .B1(new_n539), .B2(new_n573), .C1(new_n574), .C2(new_n529), .ZN(G288));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT74), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n507), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n519), .A2(G48), .B1(G651), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n529), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n507), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n539), .B2(new_n587), .C1(new_n588), .C2(new_n529), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n529), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n591), .A2(new_n594), .B1(G54), .B2(new_n519), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT75), .Z(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n507), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT76), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n590), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n590), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n602), .B2(new_n609), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n601), .A2(KEYINPUT76), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(new_n595), .B2(new_n600), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(KEYINPUT77), .ZN(new_n617));
  OAI21_X1  g192(.A(G868), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n605), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n462), .A2(new_n493), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT13), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n475), .A2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n477), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n626), .A2(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(KEYINPUT15), .B(G2435), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT79), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2430), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT78), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n640), .B(new_n646), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n647), .A2(G14), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT17), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n657), .B(new_n658), .C1(new_n656), .C2(new_n652), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n664), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  AOI22_X1  g245(.A1(new_n668), .A2(KEYINPUT20), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n664), .A3(new_n667), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n671), .B(new_n673), .C1(KEYINPUT20), .C2(new_n668), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT80), .B(G1986), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1981), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(G229));
  MUX2_X1   g256(.A(G24), .B(G290), .S(G16), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1986), .ZN(new_n683));
  OAI21_X1  g258(.A(KEYINPUT83), .B1(G16), .B2(G23), .ZN(new_n684));
  OR3_X1    g259(.A1(KEYINPUT83), .A2(G16), .A3(G23), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n684), .B(new_n685), .C1(G288), .C2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT84), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT33), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT32), .B(G1981), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G6), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G16), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G305), .B2(G16), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n696), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n692), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n699), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n701), .A2(new_n697), .A3(new_n691), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n686), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n686), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n690), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n683), .B1(new_n708), .B2(KEYINPUT34), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n475), .A2(G119), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n477), .A2(G131), .ZN(new_n712));
  NOR2_X1   g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G25), .B(new_n715), .S(G29), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT35), .B(G1991), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT81), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n690), .A2(new_n703), .A3(new_n720), .A4(new_n707), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n709), .A2(new_n710), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(KEYINPUT85), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n709), .A2(new_n719), .A3(new_n721), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n723), .B(KEYINPUT36), .C1(KEYINPUT85), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n726), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT29), .B(G2090), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n722), .A2(KEYINPUT85), .A3(new_n731), .ZN(new_n732));
  AOI22_X1  g307(.A1(G129), .A2(new_n475), .B1(new_n477), .B2(G141), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n493), .A2(G105), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT26), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n743), .B(new_n744), .C1(G29), .C2(G32), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n744), .B2(new_n743), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT27), .B(G1996), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G5), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G171), .B2(G16), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT24), .A2(G34), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n751), .A2(new_n726), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G160), .B2(new_n726), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n748), .B1(G1961), .B2(new_n750), .C1(G2084), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT93), .ZN(new_n756));
  NOR2_X1   g331(.A1(G4), .A2(G16), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n602), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1348), .ZN(new_n759));
  INV_X1    g334(.A(G1341), .ZN(new_n760));
  OR2_X1    g335(.A1(G16), .A2(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n619), .B2(new_n686), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n746), .A2(new_n747), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n760), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n686), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT94), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT23), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n569), .B2(new_n686), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT95), .B(G1956), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n686), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n686), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n726), .A2(G26), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT89), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT28), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n477), .A2(G140), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT87), .Z(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT88), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n475), .A2(G128), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2067), .ZN(new_n786));
  INV_X1    g361(.A(G1961), .ZN(new_n787));
  INV_X1    g362(.A(new_n750), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n726), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n726), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n493), .A2(G103), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT25), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n477), .A2(G139), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n795), .B(new_n796), .C1(new_n461), .C2(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G33), .B(new_n798), .S(G29), .Z(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(G2072), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(KEYINPUT90), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(KEYINPUT90), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT31), .B(G11), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n754), .A2(G2084), .ZN(new_n804));
  INV_X1    g379(.A(G28), .ZN(new_n805));
  AOI21_X1  g380(.A(G29), .B1(new_n805), .B2(KEYINPUT30), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(KEYINPUT30), .B2(new_n805), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n631), .B2(new_n726), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n799), .B2(G2072), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n789), .A2(new_n801), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n764), .A2(new_n770), .A3(new_n774), .A4(new_n811), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n756), .A2(new_n759), .A3(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n725), .A2(new_n730), .A3(new_n732), .A4(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n816), .A2(new_n539), .B1(new_n529), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n516), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n602), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n619), .A2(new_n821), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n619), .A2(new_n821), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT39), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n826), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(G860), .ZN(G145));
  XNOR2_X1  g407(.A(new_n631), .B(G160), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n481), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n475), .A2(G130), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n477), .A2(G142), .ZN(new_n836));
  NOR2_X1   g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n742), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n742), .A2(new_n839), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n624), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n741), .B(new_n839), .ZN(new_n843));
  INV_X1    g418(.A(new_n624), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n492), .B2(new_n495), .ZN(new_n848));
  INV_X1    g423(.A(new_n491), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n462), .B2(G126), .ZN(new_n850));
  OAI211_X1 g425(.A(KEYINPUT96), .B(new_n494), .C1(new_n850), .C2(new_n461), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n852), .A2(new_n853), .A3(new_n489), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n853), .B1(new_n852), .B2(new_n489), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n846), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n798), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n784), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n715), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n842), .B(new_n845), .C1(new_n855), .C2(new_n854), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n857), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n861), .B1(new_n857), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n834), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT99), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n863), .A2(new_n864), .A3(new_n834), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(new_n834), .C1(new_n863), .C2(new_n864), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g447(.A(new_n601), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n569), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n601), .A2(G299), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT100), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n602), .A2(new_n611), .A3(new_n609), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n616), .A2(KEYINPUT77), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n829), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n829), .B1(new_n878), .B2(new_n879), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n827), .A2(new_n828), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n612), .B2(new_n617), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n876), .A2(new_n886), .A3(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n874), .A2(new_n889), .A3(new_n875), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT102), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n885), .A2(new_n887), .A3(new_n880), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT101), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n885), .A2(new_n880), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT101), .B1(new_n895), .B2(new_n877), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G288), .B(G290), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G303), .B(G305), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n902), .A2(new_n901), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(KEYINPUT104), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n909), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n894), .A2(new_n897), .A3(new_n910), .A4(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n883), .B2(new_n892), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n912), .B(new_n911), .C1(new_n916), .C2(new_n896), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(G868), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n822), .A2(new_n605), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n914), .A2(new_n917), .A3(new_n921), .A4(G868), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(G295));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(G331));
  NAND2_X1  g499(.A1(new_n891), .A2(new_n887), .ZN(new_n925));
  NAND2_X1  g500(.A1(G171), .A2(KEYINPUT106), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n926), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n884), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(G171), .A2(KEYINPUT106), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n829), .A2(G168), .A3(new_n926), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n925), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n931), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n876), .B1(new_n935), .B2(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n937), .B2(new_n906), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n935), .A2(new_n932), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n888), .A3(new_n890), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n940), .B(new_n905), .C1(new_n877), .C2(new_n939), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n938), .A2(new_n941), .A3(KEYINPUT43), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n936), .A3(new_n905), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT43), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT44), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n938), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n938), .B2(new_n943), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n949), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g525(.A(KEYINPUT127), .B(KEYINPUT46), .Z(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n854), .B2(new_n855), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  AND2_X1   g529(.A1(G160), .A2(G40), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n953), .A2(KEYINPUT107), .A3(new_n954), .A4(new_n955), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n951), .B1(new_n961), .B2(G1996), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n784), .B(G2067), .Z(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n741), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT127), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n960), .B(new_n966), .C1(new_n967), .C2(KEYINPUT46), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n962), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n961), .A2(G1986), .A3(G290), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT48), .Z(new_n972));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n960), .A2(new_n973), .A3(G1996), .A4(new_n741), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n963), .B1(G1996), .B2(new_n741), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n960), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n958), .A2(G1996), .A3(new_n741), .A4(new_n959), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT108), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n974), .A2(KEYINPUT109), .A3(new_n976), .A4(new_n978), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n715), .A2(new_n717), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n715), .A2(new_n717), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n960), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n972), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT126), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n985), .B(KEYINPUT125), .Z(new_n989));
  NAND3_X1  g564(.A1(new_n981), .A2(new_n982), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n784), .A2(G2067), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n992), .B2(new_n960), .ZN(new_n993));
  AOI211_X1 g568(.A(KEYINPUT126), .B(new_n961), .C1(new_n990), .C2(new_n991), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n970), .B(new_n987), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT45), .B(new_n952), .C1(new_n854), .C2(new_n855), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n497), .A2(new_n952), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n954), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n955), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n706), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n488), .B1(new_n848), .B2(new_n851), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(G1384), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n955), .ZN(new_n1010));
  OR3_X1    g585(.A1(new_n1010), .A2(KEYINPUT112), .A3(G2090), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1000), .A2(KEYINPUT110), .A3(new_n706), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT112), .B1(new_n1010), .B2(G2090), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1003), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT55), .Z(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1016), .A3(G8), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT113), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .A4(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n954), .B1(new_n1004), .B2(G1384), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1022), .A2(KEYINPUT118), .A3(new_n955), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT118), .B1(new_n1022), .B2(new_n955), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n998), .A2(new_n954), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT119), .B1(new_n1026), .B2(G1966), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT120), .B(G2084), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1010), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1022), .A2(new_n955), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1025), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1022), .A2(KEYINPUT118), .A3(new_n955), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n773), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1027), .A2(new_n1029), .A3(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1038), .A2(G8), .A3(G168), .ZN(new_n1039));
  OR2_X1    g614(.A1(G305), .A2(G1981), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT114), .B(G86), .Z(new_n1041));
  OAI21_X1  g616(.A(new_n580), .B1(new_n529), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G1981), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(new_n1046), .A3(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1005), .A2(new_n955), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(G288), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1048), .A2(new_n1050), .B1(KEYINPUT52), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G288), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G1976), .ZN(new_n1055));
  OR3_X1    g630(.A1(new_n1052), .A2(KEYINPUT52), .A3(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1016), .B1(new_n1014), .B2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT63), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1021), .A2(new_n1039), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT63), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1021), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1057), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G288), .A2(G1976), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT115), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1040), .B1(new_n1048), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1050), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1062), .A2(new_n1064), .A3(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1027), .A2(G168), .A3(new_n1029), .A4(new_n1037), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT123), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(G8), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(KEYINPUT123), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1038), .A2(G8), .A3(G286), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1074), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1070), .A2(G8), .A3(new_n1072), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1026), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n997), .A2(new_n792), .A3(new_n955), .A4(new_n999), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1082), .A2(new_n1083), .B1(new_n787), .B2(new_n1010), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(G301), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1075), .A2(new_n1087), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1080), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1021), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1039), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n997), .A2(new_n792), .A3(new_n955), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n953), .A2(new_n954), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1084), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1096), .B2(G171), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1085), .A2(G301), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1049), .A2(G2067), .ZN(new_n1103));
  INV_X1    g678(.A(G1348), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n1010), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n873), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n997), .A2(new_n966), .A3(new_n955), .A4(new_n999), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1049), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n619), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1107), .B1(KEYINPUT59), .B2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1111), .A2(KEYINPUT59), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1006), .B1(new_n1004), .B2(G1384), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n955), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1119), .A3(new_n955), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1956), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n561), .A2(new_n1124), .A3(new_n562), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1130));
  OAI21_X1  g705(.A(G299), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1130), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n569), .A3(new_n1128), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n997), .A2(new_n955), .A3(new_n999), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1123), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1123), .A2(new_n1134), .A3(KEYINPUT61), .A4(new_n1136), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1105), .A2(new_n601), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1105), .A2(new_n601), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1114), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1123), .A2(new_n1136), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(new_n1133), .A3(new_n1131), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1096), .A2(G171), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1092), .B1(new_n1086), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1102), .A2(new_n1149), .A3(new_n1079), .A4(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1089), .A2(new_n1091), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1001), .B1(new_n1121), .B2(G2090), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1016), .B1(G8), .B2(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1057), .A2(KEYINPUT117), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1057), .A2(KEYINPUT117), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1155), .B(new_n1063), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1069), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(G290), .B(G1986), .Z(new_n1160));
  OAI211_X1 g735(.A(new_n983), .B(new_n986), .C1(new_n961), .C2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n996), .B1(new_n1159), .B2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g737(.A(G319), .ZN(new_n1164));
  NOR2_X1   g738(.A1(G227), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g739(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g740(.A1(G401), .A2(G229), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n871), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g742(.A(new_n948), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n938), .A2(new_n941), .A3(new_n946), .ZN(new_n1170));
  AOI211_X1 g744(.A(new_n1166), .B(new_n1168), .C1(new_n1169), .C2(new_n1170), .ZN(G308));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1172));
  NAND4_X1  g746(.A1(new_n1172), .A2(new_n871), .A3(new_n1165), .A4(new_n1167), .ZN(G225));
endmodule


