//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928;
  XOR2_X1   g000(.A(KEYINPUT31), .B(G50gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(KEYINPUT22), .B2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G211gat), .B(G218gat), .Z(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(KEYINPUT2), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218));
  INV_X1    g017(.A(G148gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G141gat), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(G141gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT2), .B1(new_n225), .B2(KEYINPUT78), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(new_n214), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n213), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(G228gat), .B2(G233gat), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n228), .B(KEYINPUT80), .Z(new_n233));
  AOI21_X1  g032(.A(KEYINPUT3), .B1(new_n213), .B2(new_n230), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n228), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g036(.A(G228gat), .B(G233gat), .C1(new_n237), .C2(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n206), .B1(new_n239), .B2(G22gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G22gat), .B2(new_n239), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n204), .A2(new_n205), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT84), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n241), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G64gat), .B(G92gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT76), .ZN(new_n247));
  XNOR2_X1  g046(.A(G8gat), .B(G36gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT68), .B1(KEYINPUT69), .B2(G183gat), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(KEYINPUT27), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT67), .B(G190gat), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(KEYINPUT27), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT68), .A2(KEYINPUT27), .A3(G183gat), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT27), .B(G183gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT67), .B(G190gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(new_n257), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT26), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR3_X1   g065(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n270), .A2(new_n264), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n264), .B1(new_n272), .B2(KEYINPUT23), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n273), .A3(new_n263), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT24), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n262), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G183gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n253), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT25), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n269), .A2(new_n281), .ZN(new_n282));
  OAI221_X1 g081(.A(new_n277), .B1(G183gat), .B2(G190gat), .C1(new_n276), .C2(KEYINPUT64), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(KEYINPUT64), .B2(new_n276), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n274), .A2(KEYINPUT25), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n230), .ZN(new_n291));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(G226gat), .A3(G233gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n213), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n290), .A2(new_n230), .B1(G226gat), .B2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(G226gat), .ZN(new_n297));
  INV_X1    g096(.A(G233gat), .ZN(new_n298));
  AOI211_X1 g097(.A(new_n297), .B(new_n298), .C1(new_n282), .C2(new_n289), .ZN(new_n299));
  INV_X1    g098(.A(new_n213), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n250), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n293), .A2(new_n213), .A3(new_n294), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n296), .B2(new_n299), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n249), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(KEYINPUT30), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n303), .A2(new_n304), .A3(new_n307), .A4(new_n249), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n310), .B(KEYINPUT79), .Z(new_n311));
  XNOR2_X1  g110(.A(G127gat), .B(G134gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G113gat), .B2(G120gat), .ZN(new_n316));
  XOR2_X1   g115(.A(KEYINPUT70), .B(G113gat), .Z(new_n317));
  AOI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(G113gat), .B2(G120gat), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(new_n312), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(new_n228), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT81), .ZN(new_n324));
  INV_X1    g123(.A(new_n322), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n324), .B1(new_n325), .B2(new_n236), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(KEYINPUT81), .A3(new_n228), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n311), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n311), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n233), .A2(new_n325), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n229), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT4), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n323), .A2(KEYINPUT4), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT39), .ZN(new_n337));
  OR3_X1    g136(.A1(new_n328), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  INV_X1    g138(.A(G85gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT0), .B(G57gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n336), .B2(new_n337), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n338), .A2(KEYINPUT40), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT40), .B1(new_n338), .B2(new_n344), .ZN(new_n346));
  INV_X1    g145(.A(new_n343), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n326), .A2(new_n311), .A3(new_n327), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n323), .B1(new_n332), .B2(KEYINPUT4), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n329), .B1(new_n330), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n348), .B(KEYINPUT5), .C1(new_n349), .C2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n311), .A2(KEYINPUT5), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n335), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n347), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n345), .A2(new_n346), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n245), .B1(new_n309), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT37), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n302), .B1(new_n358), .B2(new_n249), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT38), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT37), .B1(new_n295), .B2(new_n301), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT85), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n303), .B2(new_n304), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT85), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n359), .A2(new_n360), .A3(new_n362), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n303), .A2(new_n304), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n250), .B1(new_n367), .B2(KEYINPUT37), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT38), .B1(new_n368), .B2(new_n363), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n370));
  AOI211_X1 g169(.A(new_n370), .B(new_n347), .C1(new_n352), .C2(new_n354), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n355), .A2(KEYINPUT6), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n347), .A3(new_n354), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n366), .A2(new_n305), .A3(new_n369), .A4(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n357), .A2(new_n375), .A3(KEYINPUT86), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT86), .B1(new_n357), .B2(new_n375), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n290), .A2(new_n322), .ZN(new_n379));
  INV_X1    g178(.A(G227gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(new_n298), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n282), .A2(new_n325), .A3(new_n289), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n379), .A2(new_n383), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT72), .B1(new_n388), .B2(new_n381), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT72), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n390), .B(new_n382), .C1(new_n379), .C2(new_n383), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT32), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n389), .B2(new_n391), .ZN(new_n394));
  XNOR2_X1  g193(.A(G15gat), .B(G43gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G71gat), .B(G99gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  OAI221_X1 g198(.A(KEYINPUT32), .B1(new_n393), .B2(new_n399), .C1(new_n389), .C2(new_n391), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n387), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT36), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n387), .A3(new_n400), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n402), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n387), .A2(KEYINPUT73), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n398), .A2(new_n400), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n409), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(KEYINPUT36), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n355), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n370), .A3(new_n373), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n371), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n372), .A2(KEYINPUT82), .A3(new_n373), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n309), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n245), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n378), .A2(new_n414), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT35), .ZN(new_n426));
  INV_X1    g225(.A(new_n374), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n406), .A2(new_n405), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n401), .A2(new_n402), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT87), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n403), .A2(new_n432), .A3(new_n405), .A4(new_n406), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n245), .B(new_n428), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n245), .B1(new_n410), .B2(new_n411), .ZN(new_n435));
  INV_X1    g234(.A(new_n423), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n426), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n425), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(G99gat), .B(G106gat), .Z(new_n440));
  INV_X1    g239(.A(KEYINPUT7), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n441), .A2(KEYINPUT98), .B1(G85gat), .B2(G92gat), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT99), .B1(new_n441), .B2(KEYINPUT98), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT98), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT99), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT7), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT8), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(G99gat), .B2(G106gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(KEYINPUT100), .A2(G92gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(KEYINPUT100), .A2(G92gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n340), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n442), .B1(new_n443), .B2(new_n446), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n440), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT100), .B(G92gat), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n449), .B1(new_n457), .B2(new_n340), .ZN(new_n458));
  NAND2_X1  g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n444), .B2(KEYINPUT7), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n445), .B1(new_n444), .B2(KEYINPUT7), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n441), .A2(KEYINPUT98), .A3(KEYINPUT99), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n440), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n458), .A2(new_n463), .A3(new_n464), .A4(new_n447), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT101), .B1(new_n456), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(KEYINPUT101), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G29gat), .A2(G36gat), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT14), .ZN(new_n471));
  INV_X1    g270(.A(G29gat), .ZN(new_n472));
  INV_X1    g271(.A(G36gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(new_n474), .B2(KEYINPUT89), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  NOR2_X1   g275(.A1(G29gat), .A2(G36gat), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n471), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n469), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT15), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT90), .B(G50gat), .Z(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(G43gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(KEYINPUT15), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n474), .A2(new_n470), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n469), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G232gat), .A2(G233gat), .ZN(new_n490));
  XOR2_X1   g289(.A(new_n490), .B(KEYINPUT97), .Z(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT41), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n481), .A2(new_n487), .A3(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n489), .B(new_n493), .C1(new_n468), .C2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G134gat), .B(G162gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n492), .A2(KEYINPUT41), .ZN(new_n501));
  XNOR2_X1  g300(.A(G190gat), .B(G218gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n500), .A2(new_n503), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(G1gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n508), .B1(new_n510), .B2(G1gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n507), .A3(new_n511), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT9), .ZN(new_n516));
  INV_X1    g315(.A(G64gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G57gat), .ZN(new_n518));
  INV_X1    g317(.A(G57gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G64gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n516), .B1(new_n521), .B2(KEYINPUT93), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(KEYINPUT93), .B2(new_n521), .ZN(new_n523));
  XOR2_X1   g322(.A(G71gat), .B(G78gat), .Z(new_n524));
  INV_X1    g323(.A(new_n521), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(KEYINPUT94), .ZN(new_n526));
  NAND2_X1  g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  INV_X1    g326(.A(G71gat), .ZN(new_n528));
  INV_X1    g327(.A(G78gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT9), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n525), .A2(KEYINPUT94), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n523), .A2(new_n524), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n515), .B1(new_n532), .B2(KEYINPUT21), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT21), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n532), .B(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n535), .B2(new_n515), .ZN(new_n536));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT96), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT19), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT20), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n536), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT95), .ZN(new_n543));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n541), .B(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n506), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n548));
  INV_X1    g347(.A(new_n514), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(new_n512), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n513), .A2(KEYINPUT91), .A3(new_n514), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT92), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n495), .A4(new_n496), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n495), .A2(new_n496), .A3(new_n550), .A4(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT92), .ZN(new_n556));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n515), .A2(new_n488), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n554), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n515), .B(new_n488), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n557), .B(KEYINPUT13), .Z(new_n562));
  AOI22_X1  g361(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G169gat), .B(G197gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT12), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n555), .A2(KEYINPUT92), .B1(new_n488), .B2(new_n515), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n570), .A2(KEYINPUT18), .A3(new_n557), .A4(new_n554), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n569), .B1(new_n563), .B2(new_n571), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n456), .A2(new_n465), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT101), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n532), .ZN(new_n579));
  INV_X1    g378(.A(new_n467), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n532), .A2(new_n576), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT10), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n584));
  NOR4_X1   g383(.A1(new_n579), .A2(new_n466), .A3(new_n584), .A4(new_n467), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n575), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n575), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n581), .A2(new_n587), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G120gat), .B(G148gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n547), .A2(new_n574), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n439), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n421), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g401(.A1(new_n439), .A2(new_n422), .A3(new_n598), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT42), .B1(new_n603), .B2(new_n507), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT16), .B(G8gat), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  MUX2_X1   g405(.A(KEYINPUT42), .B(new_n604), .S(new_n606), .Z(G1325gat));
  NAND2_X1  g406(.A1(new_n431), .A2(new_n433), .ZN(new_n608));
  AOI21_X1  g407(.A(G15gat), .B1(new_n599), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n413), .A2(G15gat), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n599), .B2(new_n610), .ZN(G1326gat));
  NAND2_X1  g410(.A1(new_n599), .A2(new_n245), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT43), .B(G22gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(G1327gat));
  INV_X1    g413(.A(new_n546), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n572), .A2(new_n573), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n615), .A2(new_n616), .A3(new_n596), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n438), .A2(new_n506), .A3(new_n617), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n618), .A2(G29gat), .A3(new_n421), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT45), .Z(new_n620));
  OAI211_X1 g419(.A(new_n412), .B(new_n407), .C1(new_n376), .C2(new_n377), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n424), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n423), .A2(KEYINPUT102), .A3(new_n245), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI22_X1  g424(.A1(new_n434), .A2(new_n437), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n626), .A2(new_n627), .A3(new_n506), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n438), .B2(new_n506), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n617), .ZN(new_n631));
  OAI21_X1  g430(.A(G29gat), .B1(new_n631), .B2(new_n421), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n620), .A2(new_n632), .ZN(G1328gat));
  OAI21_X1  g432(.A(G36gat), .B1(new_n631), .B2(new_n422), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n618), .A2(G36gat), .A3(new_n422), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT46), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(G1329gat));
  OAI21_X1  g436(.A(G43gat), .B1(new_n631), .B2(new_n414), .ZN(new_n638));
  INV_X1    g437(.A(new_n608), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n618), .A2(G43gat), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(KEYINPUT47), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT47), .ZN(new_n643));
  INV_X1    g442(.A(G43gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n645));
  INV_X1    g444(.A(new_n617), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n647), .B2(new_n413), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n643), .B1(new_n648), .B2(new_n640), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n642), .A2(new_n649), .ZN(G1330gat));
  INV_X1    g449(.A(new_n245), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n483), .B1(new_n631), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n483), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n245), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n618), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT48), .B1(new_n655), .B2(KEYINPUT103), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n652), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n653), .B1(new_n647), .B2(new_n245), .ZN(new_n659));
  INV_X1    g458(.A(new_n655), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(G1331gat));
  AND4_X1   g461(.A1(new_n616), .A2(new_n626), .A3(new_n547), .A4(new_n596), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n600), .A2(KEYINPUT104), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n600), .A2(KEYINPUT104), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g467(.A(new_n422), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT105), .ZN(new_n671));
  OR2_X1    g470(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1333gat));
  NAND3_X1  g472(.A1(new_n663), .A2(new_n528), .A3(new_n608), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n663), .A2(new_n413), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(new_n528), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g476(.A1(new_n663), .A2(new_n245), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT106), .B(G78gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1335gat));
  NAND2_X1  g479(.A1(new_n616), .A2(new_n546), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT107), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(new_n596), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n630), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G85gat), .B1(new_n684), .B2(new_n421), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n245), .B1(new_n431), .B2(new_n433), .ZN(new_n686));
  INV_X1    g485(.A(new_n428), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n437), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n621), .A2(new_n625), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n506), .B(new_n682), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT51), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n626), .A2(KEYINPUT51), .A3(new_n506), .A4(new_n682), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n600), .A2(new_n340), .A3(new_n596), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n685), .B1(new_n695), .B2(new_n696), .ZN(G1336gat));
  NAND3_X1  g496(.A1(new_n692), .A2(KEYINPUT108), .A3(new_n693), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n690), .A2(new_n699), .A3(new_n691), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n422), .A2(new_n597), .A3(G92gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n698), .A2(new_n704), .A3(new_n700), .A4(new_n701), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n309), .B(new_n683), .C1(new_n628), .C2(new_n629), .ZN(new_n706));
  INV_X1    g505(.A(new_n457), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT52), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT52), .B1(new_n694), .B2(new_n701), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1337gat));
  OAI21_X1  g512(.A(G99gat), .B1(new_n684), .B2(new_n414), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n639), .A2(G99gat), .A3(new_n597), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT110), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n695), .B2(new_n716), .ZN(G1338gat));
  NOR3_X1   g516(.A1(new_n651), .A2(G106gat), .A3(new_n597), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT111), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n698), .A2(new_n700), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT112), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n698), .A2(new_n722), .A3(new_n700), .A4(new_n719), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n245), .B(new_n683), .C1(new_n628), .C2(new_n629), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G106gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT53), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT53), .B1(new_n694), .B2(new_n718), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1339gat));
  INV_X1    g529(.A(new_n506), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n592), .B1(new_n586), .B2(KEYINPUT54), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n466), .A2(new_n532), .A3(new_n467), .ZN(new_n733));
  INV_X1    g532(.A(new_n582), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n584), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n468), .A2(KEYINPUT10), .A3(new_n532), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n736), .A3(new_n587), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n586), .A2(KEYINPUT54), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n586), .A2(new_n737), .A3(KEYINPUT113), .A4(KEYINPUT54), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n732), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n593), .B1(new_n742), .B2(KEYINPUT55), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT114), .B1(new_n742), .B2(KEYINPUT55), .ZN(new_n744));
  INV_X1    g543(.A(new_n732), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT54), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n735), .A2(new_n736), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(new_n575), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT113), .B1(new_n748), .B2(new_n737), .ZN(new_n749));
  AND4_X1   g548(.A1(KEYINPUT113), .A2(new_n586), .A3(KEYINPUT54), .A4(new_n737), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n743), .A2(new_n744), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n743), .A2(new_n744), .A3(new_n754), .A4(KEYINPUT115), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n616), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n557), .B1(new_n570), .B2(new_n554), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n561), .A2(new_n562), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n568), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n596), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n731), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n506), .A2(new_n760), .A3(new_n763), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n757), .B2(new_n758), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n615), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n547), .A2(new_n616), .A3(new_n597), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n773), .A2(new_n422), .A3(new_n666), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n435), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT117), .ZN(new_n776));
  INV_X1    g575(.A(new_n317), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n574), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n773), .A2(new_n686), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n421), .A2(new_n309), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n574), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n784), .A3(G113gat), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n783), .B2(G113gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n778), .B1(new_n786), .B2(new_n787), .ZN(G1340gat));
  INV_X1    g587(.A(G120gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n776), .A2(new_n789), .A3(new_n596), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n782), .A2(new_n596), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(KEYINPUT118), .A3(G120gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT118), .B1(new_n791), .B2(G120gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(G1341gat));
  INV_X1    g594(.A(G127gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n796), .A3(new_n546), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n774), .A2(new_n435), .A3(new_n615), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n796), .ZN(G1342gat));
  OR3_X1    g598(.A1(new_n775), .A2(G134gat), .A3(new_n731), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n800), .A2(KEYINPUT56), .ZN(new_n801));
  OAI21_X1  g600(.A(G134gat), .B1(new_n781), .B2(new_n731), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(KEYINPUT56), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(G1343gat));
  NAND2_X1  g603(.A1(new_n414), .A2(new_n780), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n773), .A2(new_n245), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n651), .A2(new_n807), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n751), .A2(new_n753), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n743), .A2(new_n574), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n506), .B1(new_n812), .B2(new_n764), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n546), .B1(new_n768), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n810), .B1(new_n814), .B2(new_n771), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT119), .Z(new_n816));
  AOI21_X1  g615(.A(new_n805), .B1(new_n808), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n221), .B1(new_n817), .B2(new_n574), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n413), .A2(new_n651), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n774), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(G141gat), .A3(new_n616), .ZN(new_n821));
  OR3_X1    g620(.A1(new_n818), .A2(KEYINPUT58), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT58), .B1(new_n818), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1344gat));
  INV_X1    g623(.A(new_n820), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n219), .A3(new_n596), .ZN(new_n826));
  AOI211_X1 g625(.A(KEYINPUT59), .B(new_n219), .C1(new_n817), .C2(new_n596), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828));
  OAI211_X1 g627(.A(KEYINPUT57), .B(new_n245), .C1(new_n770), .C2(new_n772), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n755), .A2(new_n767), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n546), .B1(new_n813), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n651), .B1(new_n832), .B2(new_n771), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n833), .B2(KEYINPUT57), .ZN(new_n834));
  INV_X1    g633(.A(new_n767), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(new_n754), .A3(new_n743), .A4(new_n744), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n616), .B1(new_n753), .B2(new_n751), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n765), .B1(new_n837), .B2(new_n743), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n838), .B2(new_n506), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n772), .B1(new_n839), .B2(new_n546), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT120), .B(new_n807), .C1(new_n840), .C2(new_n651), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n834), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n829), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(new_n414), .A3(new_n596), .A4(new_n780), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n828), .B1(new_n844), .B2(G148gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n826), .B1(new_n827), .B2(new_n845), .ZN(G1345gat));
  XNOR2_X1  g645(.A(KEYINPUT78), .B(G155gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n825), .A2(new_n615), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n817), .A2(new_n615), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n847), .ZN(G1346gat));
  INV_X1    g649(.A(G162gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n825), .A2(new_n851), .A3(new_n506), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n817), .A2(new_n506), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(G1347gat));
  NAND2_X1  g653(.A1(new_n773), .A2(new_n421), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n422), .B1(new_n855), .B2(KEYINPUT121), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n773), .A2(new_n857), .A3(new_n421), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n435), .ZN(new_n860));
  INV_X1    g659(.A(G169gat), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n574), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n422), .B1(new_n664), .B2(new_n665), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n773), .A2(new_n686), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G169gat), .B1(new_n866), .B2(new_n616), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n867), .ZN(G1348gat));
  NAND2_X1  g667(.A1(new_n860), .A2(new_n596), .ZN(new_n869));
  INV_X1    g668(.A(G176gat), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n864), .B(KEYINPUT122), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n597), .A2(new_n870), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n869), .A2(new_n870), .B1(new_n871), .B2(new_n872), .ZN(G1349gat));
  OAI21_X1  g672(.A(G183gat), .B1(new_n866), .B2(new_n546), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n615), .A2(new_n258), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n435), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT60), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n874), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n860), .A2(new_n253), .A3(new_n506), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n871), .A2(new_n506), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(new_n884), .A3(G190gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n883), .B2(G190gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(G1351gat));
  AND2_X1   g686(.A1(new_n859), .A2(new_n819), .ZN(new_n888));
  INV_X1    g687(.A(G197gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n574), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n414), .A2(new_n863), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n843), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n829), .A2(new_n842), .A3(KEYINPUT123), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G197gat), .B1(new_n895), .B2(new_n616), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n890), .A2(new_n896), .ZN(G1352gat));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n895), .B2(new_n597), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n893), .A2(KEYINPUT125), .A3(new_n596), .A4(new_n894), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(G204gat), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n597), .A2(G204gat), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n856), .A2(new_n819), .A3(new_n858), .A4(new_n902), .ZN(new_n903));
  OR3_X1    g702(.A1(new_n903), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(KEYINPUT62), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT124), .B1(new_n903), .B2(KEYINPUT62), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n901), .A2(new_n904), .A3(new_n905), .A4(new_n906), .ZN(G1353gat));
  NOR2_X1   g706(.A1(new_n546), .A2(G211gat), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n856), .A2(new_n819), .A3(new_n858), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n414), .A2(new_n863), .A3(new_n615), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n843), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n208), .B1(new_n912), .B2(KEYINPUT126), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT126), .B(new_n910), .C1(new_n829), .C2(new_n842), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT63), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n829), .B2(new_n842), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918));
  OAI21_X1  g717(.A(G211gat), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(new_n914), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n909), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT127), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n924), .B(new_n909), .C1(new_n916), .C2(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1354gat));
  NOR3_X1   g725(.A1(new_n895), .A2(new_n209), .A3(new_n731), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n888), .A2(new_n506), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n209), .ZN(G1355gat));
endmodule


