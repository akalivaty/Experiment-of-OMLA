//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(KEYINPUT23), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(G169gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(G176gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(KEYINPUT25), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT67), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n213), .A2(new_n218), .A3(new_n214), .A4(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n214), .A2(KEYINPUT24), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n221), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT68), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226));
  AOI211_X1 g025(.A(new_n226), .B(new_n223), .C1(new_n217), .C2(new_n219), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n212), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT69), .B(new_n212), .C1(new_n225), .C2(new_n227), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n224), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT64), .B(G176gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n232), .B(new_n207), .C1(new_n209), .C2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n230), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT27), .B(G183gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT28), .B1(new_n242), .B2(KEYINPUT70), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NOR2_X1   g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247));
  NOR4_X1   g046(.A1(KEYINPUT71), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n249), .B1(new_n247), .B2(new_n246), .ZN(new_n250));
  OAI221_X1 g049(.A(new_n203), .B1(new_n246), .B2(new_n247), .C1(new_n248), .C2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n244), .A2(new_n245), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT29), .B1(new_n237), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT76), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n202), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n255), .ZN(new_n257));
  INV_X1    g056(.A(new_n252), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n228), .A2(new_n229), .B1(new_n235), .B2(new_n234), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(new_n231), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT77), .B(new_n257), .C1(new_n260), .C2(KEYINPUT29), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(G211gat), .A2(G218gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G211gat), .ZN(new_n267));
  INV_X1    g066(.A(G218gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n263), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(new_n262), .A3(new_n265), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n218), .B1(new_n240), .B2(new_n214), .ZN(new_n275));
  INV_X1    g074(.A(new_n219), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n224), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n226), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n220), .A2(KEYINPUT68), .A3(new_n224), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n211), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n236), .B1(new_n280), .B2(KEYINPUT69), .ZN(new_n281));
  INV_X1    g080(.A(new_n231), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n252), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n274), .B1(new_n283), .B2(new_n255), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n256), .A2(new_n261), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT78), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n255), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n253), .B2(new_n255), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n274), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT78), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n256), .A2(new_n261), .A3(new_n290), .A4(new_n284), .ZN(new_n291));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  NAND4_X1  g093(.A1(new_n286), .A2(new_n289), .A3(new_n291), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n291), .A2(new_n289), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n298), .A2(KEYINPUT30), .A3(new_n286), .A4(new_n294), .ZN(new_n299));
  INV_X1    g098(.A(new_n294), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n285), .A2(KEYINPUT78), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n291), .A2(new_n289), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n305));
  XNOR2_X1  g104(.A(G1gat), .B(G29gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT0), .ZN(new_n307));
  XOR2_X1   g106(.A(G57gat), .B(G85gat), .Z(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G148gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G141gat), .ZN(new_n311));
  INV_X1    g110(.A(G141gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G148gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n315), .A2(KEYINPUT81), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n315), .A2(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n314), .A2(KEYINPUT80), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(KEYINPUT80), .B2(new_n314), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(KEYINPUT79), .B2(new_n322), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n312), .A2(KEYINPUT82), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G141gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n328), .A3(G148gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT83), .B1(new_n329), .B2(new_n311), .ZN(new_n330));
  NOR2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n322), .B1(new_n315), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n329), .A2(KEYINPUT83), .A3(new_n311), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n325), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G127gat), .B(G134gat), .Z(new_n337));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT72), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(KEYINPUT1), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n342), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT4), .B1(new_n336), .B2(new_n345), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n319), .A2(new_n324), .B1(new_n333), .B2(new_n334), .ZN(new_n347));
  INV_X1    g146(.A(new_n345), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(KEYINPUT85), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n336), .B2(KEYINPUT3), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n347), .A2(new_n348), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT4), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n309), .B1(new_n362), .B2(KEYINPUT39), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n336), .A2(new_n345), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n356), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT39), .B1(new_n365), .B2(new_n361), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(new_n359), .B2(new_n361), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n305), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n368), .A2(KEYINPUT40), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT5), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n365), .B2(new_n361), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n347), .A2(new_n348), .A3(new_n372), .A4(new_n349), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n360), .A3(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n346), .A2(KEYINPUT84), .A3(new_n350), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n361), .B1(new_n352), .B2(new_n354), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n377), .A2(new_n351), .A3(new_n370), .A4(new_n358), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n309), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n368), .B2(KEYINPUT40), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n369), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n304), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n274), .A2(KEYINPUT29), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n383), .A2(KEYINPUT88), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n353), .B1(new_n383), .B2(KEYINPUT88), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n336), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n354), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n274), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n386), .A2(G228gat), .A3(new_n389), .A4(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(G22gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n273), .B1(new_n354), .B2(new_n387), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n270), .A2(KEYINPUT87), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n394), .B(new_n387), .C1(new_n395), .C2(new_n273), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n347), .B1(new_n396), .B2(new_n353), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n392), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n390), .A2(new_n391), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n391), .B1(new_n390), .B2(new_n398), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT31), .B(G50gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT86), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OR4_X1    g204(.A1(KEYINPUT89), .A2(new_n399), .A3(new_n400), .A4(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT89), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n404), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n400), .B2(new_n399), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT38), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n300), .A2(KEYINPUT37), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n303), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n286), .A2(new_n289), .A3(new_n291), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT37), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT37), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n288), .B2(new_n273), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n256), .A2(new_n261), .A3(new_n274), .A4(new_n287), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT38), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(new_n300), .C1(new_n414), .C2(KEYINPUT37), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n376), .A2(new_n309), .A3(new_n378), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n422), .A2(new_n379), .A3(KEYINPUT6), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424));
  AOI211_X1 g223(.A(new_n424), .B(new_n309), .C1(new_n376), .C2(new_n378), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n426), .A3(new_n295), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n382), .B(new_n410), .C1(new_n416), .C2(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n423), .A2(new_n425), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(new_n297), .A3(new_n303), .A4(new_n299), .ZN(new_n430));
  INV_X1    g229(.A(new_n410), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT74), .B(G71gat), .ZN(new_n433));
  INV_X1    g232(.A(G99gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G15gat), .B(G43gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n348), .B(new_n252), .C1(new_n281), .C2(new_n282), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n237), .A2(KEYINPUT73), .A3(new_n348), .A4(new_n252), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n283), .A2(new_n345), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G227gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n437), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n348), .B1(new_n237), .B2(new_n252), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n439), .B2(new_n438), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT34), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n444), .A4(new_n441), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n440), .A2(new_n442), .A3(new_n444), .A4(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT34), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n446), .A2(KEYINPUT32), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT33), .B1(new_n443), .B2(new_n445), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n454), .B(new_n452), .C1(new_n459), .C2(new_n437), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n458), .B1(new_n456), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT75), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n465), .ZN(new_n467));
  NAND2_X1  g266(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(new_n468), .C1(new_n461), .C2(new_n462), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n428), .A2(new_n432), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n456), .A2(new_n460), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n457), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n410), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT91), .B1(new_n474), .B2(new_n430), .ZN(new_n475));
  AND4_X1   g274(.A1(new_n429), .A2(new_n297), .A3(new_n303), .A4(new_n299), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n463), .A3(new_n477), .A4(new_n410), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n478), .A3(KEYINPUT35), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT91), .B(new_n480), .C1(new_n474), .C2(new_n430), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n470), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT18), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT96), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT95), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(G43gat), .A2(G50gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(G43gat), .A2(G50gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(KEYINPUT93), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n499));
  AOI21_X1  g298(.A(G36gat), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n497), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n500), .A2(new_n501), .B1(KEYINPUT15), .B2(new_n489), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT94), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n491), .B(new_n494), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n503), .B2(new_n505), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n486), .B(new_n487), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n505), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT94), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT17), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n509), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT95), .B1(new_n513), .B2(new_n487), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n508), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G1gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G1gat), .B2(new_n516), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(G8gat), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n520), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n510), .A2(new_n511), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n485), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n526), .B(KEYINPUT13), .Z(new_n529));
  INV_X1    g328(.A(new_n524), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n522), .A2(new_n523), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n521), .A2(new_n526), .A3(new_n524), .A4(new_n484), .ZN(new_n533));
  XOR2_X1   g332(.A(G113gat), .B(G141gat), .Z(new_n534));
  XNOR2_X1  g333(.A(G169gat), .B(G197gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  XOR2_X1   g337(.A(new_n538), .B(KEYINPUT12), .Z(new_n539));
  NAND4_X1  g338(.A1(new_n528), .A2(new_n532), .A3(new_n533), .A4(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n539), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n532), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n530), .B1(new_n515), .B2(new_n520), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n484), .B1(new_n543), .B2(new_n526), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n482), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  OR2_X1    g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n552));
  INV_X1    g351(.A(G57gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(G64gat), .ZN(new_n554));
  INV_X1    g353(.A(G64gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(G57gat), .B2(new_n555), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n552), .A2(new_n553), .A3(G64gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n551), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n553), .A2(G64gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n555), .A2(G57gat), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT9), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n548), .A3(new_n549), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G127gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n563), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n522), .B1(KEYINPUT21), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n567), .B(G127gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n571), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n577));
  INV_X1    g376(.A(G155gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n576), .B(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT101), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT7), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(G85gat), .A3(G92gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n592), .B2(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n597), .A2(new_n601), .A3(new_n599), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(KEYINPUT98), .A3(new_n602), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(new_n610));
  OAI22_X1  g409(.A1(new_n609), .A2(new_n610), .B1(new_n506), .B2(new_n507), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n589), .A2(new_n590), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT100), .B1(new_n609), .B2(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n606), .A2(new_n608), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT99), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI211_X1 g420(.A(new_n591), .B(new_n613), .C1(new_n621), .C2(new_n515), .ZN(new_n622));
  INV_X1    g421(.A(new_n591), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n515), .A2(new_n614), .A3(new_n619), .ZN(new_n624));
  INV_X1    g423(.A(new_n613), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n588), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n487), .B1(new_n506), .B2(new_n507), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n628), .B(KEYINPUT95), .C1(new_n487), .C2(new_n513), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n620), .B1(new_n629), .B2(new_n508), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n591), .B1(new_n630), .B2(new_n613), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n624), .A2(new_n623), .A3(new_n625), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(new_n587), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n603), .A2(new_n605), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n563), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n615), .A2(new_n563), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT10), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n570), .A2(KEYINPUT10), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n616), .B2(new_n618), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n635), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT102), .ZN(new_n644));
  INV_X1    g443(.A(new_n635), .ZN(new_n645));
  OAI211_X1 g444(.A(KEYINPUT10), .B(new_n570), .C1(new_n609), .C2(new_n610), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n570), .B1(new_n606), .B2(new_n608), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n637), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n648), .A2(new_n637), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n645), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  AND2_X1   g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n644), .A2(new_n652), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n657), .B1(new_n643), .B2(new_n654), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n583), .A2(new_n634), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n547), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n429), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT103), .B(G1gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1324gat));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(KEYINPUT104), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n547), .A2(new_n304), .A3(new_n664), .ZN(new_n673));
  AOI211_X1 g472(.A(new_n672), .B(new_n673), .C1(KEYINPUT104), .C2(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(G8gat), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n670), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n671), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n674), .B1(new_n675), .B2(new_n677), .ZN(G1325gat));
  NAND2_X1  g477(.A1(new_n466), .A2(new_n469), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n665), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n463), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n665), .B2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n665), .A2(new_n410), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  OR2_X1    g486(.A1(new_n660), .A2(new_n661), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n583), .A2(new_n688), .A3(new_n634), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n547), .A2(new_n497), .A3(new_n426), .A4(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT45), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n583), .B(KEYINPUT105), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n546), .A3(new_n662), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT106), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n627), .A2(new_n633), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n482), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n699), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n482), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n696), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n497), .B1(new_n707), .B2(new_n426), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n691), .A2(new_n708), .ZN(G1328gat));
  NAND2_X1  g508(.A1(new_n547), .A2(new_n689), .ZN(new_n710));
  INV_X1    g509(.A(new_n304), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(G36gat), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT46), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n482), .A2(new_n702), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n706), .B1(new_n714), .B2(new_n701), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n304), .A3(new_n695), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n707), .A2(KEYINPUT108), .A3(new_n304), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(G36gat), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n720), .ZN(G1329gat));
  AND3_X1   g520(.A1(new_n482), .A2(new_n702), .A3(new_n705), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n679), .B(new_n695), .C1(new_n722), .C2(new_n703), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n715), .A2(KEYINPUT110), .A3(new_n679), .A4(new_n695), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n726), .A3(G43gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n682), .A2(G43gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n547), .A2(new_n689), .A3(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n723), .A2(G43gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n547), .A2(KEYINPUT109), .A3(new_n689), .A4(new_n728), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n732), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n731), .A2(new_n738), .ZN(G1330gat));
  OAI211_X1 g538(.A(new_n431), .B(new_n695), .C1(new_n722), .C2(new_n703), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT111), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n410), .A2(G50gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n547), .A2(new_n689), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n741), .B(new_n744), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  XNOR2_X1  g548(.A(new_n576), .B(new_n581), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n546), .A2(new_n702), .A3(new_n750), .A4(new_n662), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n482), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n429), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(new_n553), .ZN(G1332gat));
  NOR2_X1   g553(.A1(new_n752), .A2(new_n711), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n752), .B2(new_n680), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n682), .A2(G71gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n752), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g562(.A1(new_n752), .A2(new_n410), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g564(.A1(new_n546), .A2(new_n583), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n688), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n704), .B2(new_n706), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n426), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G85gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n482), .A2(new_n702), .A3(new_n766), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n482), .A2(KEYINPUT51), .A3(new_n702), .A4(new_n766), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n773), .A2(KEYINPUT112), .A3(new_n774), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n688), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n426), .A2(new_n592), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n770), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  NOR3_X1   g580(.A1(new_n711), .A2(G92gat), .A3(new_n662), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(new_n775), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n767), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n304), .B(new_n784), .C1(new_n722), .C2(new_n703), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n783), .B1(new_n593), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n771), .A2(new_n788), .A3(KEYINPUT51), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT51), .B1(new_n771), .B2(new_n788), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n791), .A2(new_n782), .B1(G92gat), .B2(new_n785), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(G1337gat));
  NAND2_X1  g593(.A1(new_n768), .A2(new_n679), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G99gat), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n463), .A2(new_n434), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n779), .B2(new_n797), .ZN(G1338gat));
  OAI211_X1 g597(.A(new_n431), .B(new_n784), .C1(new_n722), .C2(new_n703), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n410), .A2(G106gat), .A3(new_n662), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n789), .A2(new_n790), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n775), .A2(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT114), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n799), .B2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n775), .A2(new_n808), .A3(new_n801), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(new_n810), .ZN(G1339gat));
  NOR2_X1   g610(.A1(new_n702), .A2(new_n750), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n540), .A2(new_n545), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n662), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT115), .B1(new_n663), .B2(new_n546), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n525), .A2(new_n527), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n530), .A2(new_n531), .A3(new_n529), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n538), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n542), .A2(new_n544), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n539), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n646), .A2(new_n649), .A3(new_n645), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n644), .A3(new_n652), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n657), .B1(new_n650), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n827), .A3(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n827), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n660), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n822), .A2(new_n702), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n830), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(new_n659), .A3(new_n828), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n702), .A4(new_n822), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n835), .A2(new_n546), .B1(new_n822), .B2(new_n688), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n833), .B(new_n837), .C1(new_n838), .C2(new_n702), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n817), .B1(new_n693), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n429), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n474), .A2(new_n304), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n546), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n840), .A2(new_n431), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n846), .A2(new_n426), .A3(new_n711), .A4(new_n463), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT117), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n546), .A2(G113gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(G1340gat));
  AOI21_X1  g649(.A(G120gat), .B1(new_n844), .B2(new_n688), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n688), .A2(G120gat), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n848), .B2(new_n852), .ZN(G1341gat));
  INV_X1    g652(.A(new_n848), .ZN(new_n854));
  OAI21_X1  g653(.A(G127gat), .B1(new_n854), .B2(new_n693), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n844), .A2(new_n568), .A3(new_n583), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  OAI21_X1  g656(.A(G134gat), .B1(new_n854), .B2(new_n634), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n843), .A2(G134gat), .A3(new_n634), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT56), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1343gat));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n840), .B2(new_n429), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n839), .A2(new_n693), .ZN(new_n865));
  INV_X1    g664(.A(new_n817), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n426), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n679), .A2(new_n410), .A3(new_n304), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n813), .A2(G141gat), .ZN(new_n871));
  AND4_X1   g670(.A1(new_n864), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n817), .B1(new_n750), .B2(new_n839), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT57), .B1(new_n873), .B2(new_n410), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(new_n820), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n688), .A2(new_n540), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n834), .A2(new_n659), .A3(new_n828), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n813), .B2(new_n878), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n879), .A2(new_n634), .B1(new_n832), .B2(KEYINPUT116), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n692), .B1(new_n880), .B2(new_n837), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n875), .B(new_n431), .C1(new_n881), .C2(new_n817), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n679), .A2(new_n429), .A3(new_n304), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n874), .A2(new_n546), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n326), .A2(new_n328), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n872), .B1(new_n887), .B2(KEYINPUT118), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n884), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n863), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n872), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n862), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n890), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n889), .B1(new_n884), .B2(new_n886), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n897), .A2(new_n898), .A3(new_n872), .ZN(new_n899));
  OAI211_X1 g698(.A(KEYINPUT121), .B(new_n894), .C1(new_n899), .C2(new_n863), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n874), .A2(new_n882), .A3(new_n883), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n902), .B(G148gat), .C1(new_n903), .C2(new_n662), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT57), .B(new_n431), .C1(new_n881), .C2(new_n817), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n867), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n431), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n832), .B1(new_n838), .B2(new_n702), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n909), .A2(new_n750), .B1(new_n813), .B2(new_n664), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n875), .B1(new_n910), .B2(new_n410), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n688), .A3(new_n883), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G148gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT123), .B1(new_n914), .B2(KEYINPUT59), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  AOI211_X1 g715(.A(new_n916), .B(new_n902), .C1(new_n913), .C2(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n904), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n869), .A2(new_n864), .A3(new_n870), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n919), .A2(G148gat), .A3(new_n662), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1345gat));
  OAI21_X1  g720(.A(G155gat), .B1(new_n903), .B2(new_n693), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n583), .A2(new_n578), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n919), .B2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n903), .B2(new_n634), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n634), .A2(G162gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n919), .B2(new_n926), .ZN(G1347gat));
  NAND2_X1  g726(.A1(new_n304), .A2(new_n429), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n682), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n846), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(new_n208), .A3(new_n813), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n840), .A2(new_n426), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT124), .B1(new_n474), .B2(new_n711), .ZN(new_n933));
  OR3_X1    g732(.A1(new_n474), .A2(new_n711), .A3(KEYINPUT124), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n546), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n931), .B1(new_n937), .B2(new_n208), .ZN(G1348gat));
  AOI21_X1  g737(.A(G176gat), .B1(new_n936), .B2(new_n688), .ZN(new_n939));
  INV_X1    g738(.A(new_n930), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n688), .A2(new_n233), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G1349gat));
  OAI21_X1  g741(.A(G183gat), .B1(new_n930), .B2(new_n693), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n583), .A2(new_n241), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n935), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n936), .A2(new_n240), .A3(new_n702), .ZN(new_n947));
  OAI21_X1  g746(.A(G190gat), .B1(new_n930), .B2(new_n634), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT125), .ZN(G1351gat));
  NOR4_X1   g751(.A1(new_n840), .A2(new_n679), .A3(new_n410), .A4(new_n928), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n546), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n679), .A2(new_n928), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT126), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n912), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n546), .A2(G197gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1352gat));
  AOI21_X1  g758(.A(G204gat), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n953), .A2(new_n688), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n912), .A2(new_n956), .A3(new_n688), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G204gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1353gat));
  NAND3_X1  g765(.A1(new_n953), .A2(new_n267), .A3(new_n583), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n267), .B1(new_n957), .B2(new_n583), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT63), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  NAND3_X1  g770(.A1(new_n953), .A2(new_n268), .A3(new_n702), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n957), .A2(new_n702), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n268), .ZN(G1355gat));
endmodule


