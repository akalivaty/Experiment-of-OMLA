

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592;

  XNOR2_X1 U326 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U327 ( .A(G183GAT), .ZN(n446) );
  XNOR2_X1 U328 ( .A(n454), .B(n453), .ZN(n536) );
  XOR2_X1 U329 ( .A(G85GAT), .B(KEYINPUT72), .Z(n294) );
  INV_X1 U330 ( .A(KEYINPUT46), .ZN(n399) );
  INV_X1 U331 ( .A(KEYINPUT54), .ZN(n413) );
  INV_X1 U332 ( .A(KEYINPUT23), .ZN(n428) );
  XNOR2_X1 U333 ( .A(n413), .B(KEYINPUT121), .ZN(n414) );
  XNOR2_X1 U334 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U335 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U336 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U337 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U338 ( .A(n449), .B(n448), .ZN(n452) );
  XNOR2_X1 U339 ( .A(n381), .B(n380), .ZN(n582) );
  XOR2_X1 U340 ( .A(n436), .B(n435), .Z(n468) );
  INV_X1 U341 ( .A(G190GAT), .ZN(n456) );
  XOR2_X1 U342 ( .A(KEYINPUT110), .B(n480), .Z(n532) );
  XOR2_X1 U343 ( .A(KEYINPUT28), .B(n468), .Z(n539) );
  XNOR2_X1 U344 ( .A(n456), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U345 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U346 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U347 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n491), .B(n490), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(G92GAT), .B(KEYINPUT11), .Z(n296) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n312) );
  XOR2_X1 U352 ( .A(KEYINPUT76), .B(KEYINPUT79), .Z(n298) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U355 ( .A(n299), .B(KEYINPUT75), .Z(n304) );
  XOR2_X1 U356 ( .A(G29GAT), .B(G43GAT), .Z(n301) );
  XNOR2_X1 U357 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n396) );
  XNOR2_X1 U359 ( .A(G99GAT), .B(G106GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n294), .B(n302), .ZN(n369) );
  XNOR2_X1 U361 ( .A(n396), .B(n369), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U363 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n306) );
  XOR2_X1 U364 ( .A(G50GAT), .B(G162GAT), .Z(n420) );
  XOR2_X1 U365 ( .A(G36GAT), .B(G190GAT), .Z(n332) );
  XNOR2_X1 U366 ( .A(n420), .B(n332), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U368 ( .A(n308), .B(n307), .Z(n310) );
  XNOR2_X1 U369 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n547) );
  INV_X1 U372 ( .A(n547), .ZN(n561) );
  XOR2_X1 U373 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n314) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(KEYINPUT91), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n331) );
  XNOR2_X1 U376 ( .A(G113GAT), .B(G134GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n315), .B(KEYINPUT0), .ZN(n450) );
  XNOR2_X1 U378 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n316), .B(KEYINPUT2), .ZN(n427) );
  XNOR2_X1 U380 ( .A(n450), .B(n427), .ZN(n329) );
  XOR2_X1 U381 ( .A(G85GAT), .B(G155GAT), .Z(n318) );
  XNOR2_X1 U382 ( .A(G29GAT), .B(G162GAT), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U384 ( .A(G57GAT), .B(G148GAT), .Z(n320) );
  XNOR2_X1 U385 ( .A(G127GAT), .B(G120GAT), .ZN(n319) );
  XNOR2_X1 U386 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U387 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U388 ( .A(KEYINPUT1), .B(KEYINPUT90), .Z(n324) );
  NAND2_X1 U389 ( .A1(G225GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U390 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U391 ( .A(KEYINPUT6), .B(n325), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n526) );
  XOR2_X1 U395 ( .A(G169GAT), .B(G8GAT), .Z(n395) );
  XNOR2_X1 U396 ( .A(n395), .B(n332), .ZN(n346) );
  XOR2_X1 U397 ( .A(G183GAT), .B(KEYINPUT80), .Z(n360) );
  XOR2_X1 U398 ( .A(KEYINPUT92), .B(n360), .Z(n334) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n337) );
  XOR2_X1 U401 ( .A(G64GAT), .B(G92GAT), .Z(n336) );
  XNOR2_X1 U402 ( .A(G176GAT), .B(G204GAT), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n375) );
  XOR2_X1 U404 ( .A(n337), .B(n375), .Z(n344) );
  XOR2_X1 U405 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n339) );
  XNOR2_X1 U406 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U408 ( .A(KEYINPUT17), .B(n340), .Z(n454) );
  XOR2_X1 U409 ( .A(G211GAT), .B(KEYINPUT21), .Z(n342) );
  XNOR2_X1 U410 ( .A(G197GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U411 ( .A(n342), .B(n341), .ZN(n433) );
  XNOR2_X1 U412 ( .A(n454), .B(n433), .ZN(n343) );
  XNOR2_X1 U413 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n346), .B(n345), .ZN(n529) );
  XNOR2_X1 U415 ( .A(KEYINPUT120), .B(n529), .ZN(n412) );
  XOR2_X1 U416 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n404) );
  XOR2_X1 U417 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n352) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n348) );
  XNOR2_X1 U419 ( .A(KEYINPUT81), .B(KEYINPUT83), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n348), .B(n347), .ZN(n350) );
  XNOR2_X1 U421 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n349), .B(KEYINPUT13), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n350), .B(n366), .ZN(n351) );
  XNOR2_X1 U424 ( .A(n352), .B(n351), .ZN(n359) );
  XOR2_X1 U425 ( .A(KEYINPUT82), .B(G64GAT), .Z(n354) );
  XNOR2_X1 U426 ( .A(G211GAT), .B(G78GAT), .ZN(n353) );
  XNOR2_X1 U427 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U428 ( .A(n355), .B(G71GAT), .Z(n357) );
  XOR2_X1 U429 ( .A(KEYINPUT67), .B(G1GAT), .Z(n393) );
  XNOR2_X1 U430 ( .A(G8GAT), .B(n393), .ZN(n356) );
  XNOR2_X1 U431 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U432 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U433 ( .A(G15GAT), .B(G127GAT), .Z(n441) );
  XOR2_X1 U434 ( .A(G22GAT), .B(G155GAT), .Z(n419) );
  XOR2_X1 U435 ( .A(n419), .B(n360), .Z(n362) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U437 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U438 ( .A(n441), .B(n363), .ZN(n364) );
  XOR2_X1 U439 ( .A(n365), .B(n364), .Z(n571) );
  INV_X1 U440 ( .A(n571), .ZN(n586) );
  XOR2_X1 U441 ( .A(KEYINPUT70), .B(KEYINPUT32), .Z(n368) );
  XOR2_X1 U442 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XNOR2_X1 U443 ( .A(n442), .B(n366), .ZN(n367) );
  XOR2_X1 U444 ( .A(n368), .B(n367), .Z(n373) );
  XOR2_X1 U445 ( .A(n369), .B(KEYINPUT69), .Z(n371) );
  NAND2_X1 U446 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U447 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U448 ( .A(n373), .B(n372), .ZN(n381) );
  XNOR2_X1 U449 ( .A(G78GAT), .B(KEYINPUT71), .ZN(n374) );
  XOR2_X1 U450 ( .A(n374), .B(G148GAT), .Z(n434) );
  XOR2_X1 U451 ( .A(n434), .B(n375), .Z(n379) );
  XOR2_X1 U452 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n377) );
  XNOR2_X1 U453 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n376) );
  XOR2_X1 U454 ( .A(n377), .B(n376), .Z(n378) );
  XOR2_X1 U455 ( .A(KEYINPUT41), .B(n582), .Z(n555) );
  XOR2_X1 U456 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n383) );
  NAND2_X1 U457 ( .A1(G229GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U458 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U459 ( .A(n384), .B(KEYINPUT30), .Z(n392) );
  XOR2_X1 U460 ( .A(G22GAT), .B(G141GAT), .Z(n386) );
  XNOR2_X1 U461 ( .A(G50GAT), .B(G36GAT), .ZN(n385) );
  XNOR2_X1 U462 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U463 ( .A(KEYINPUT66), .B(G15GAT), .Z(n388) );
  XNOR2_X1 U464 ( .A(G197GAT), .B(G113GAT), .ZN(n387) );
  XNOR2_X1 U465 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U466 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U467 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U468 ( .A(n394), .B(n393), .Z(n398) );
  XNOR2_X1 U469 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U470 ( .A(n398), .B(n397), .Z(n579) );
  INV_X1 U471 ( .A(n579), .ZN(n563) );
  OR2_X1 U472 ( .A1(n555), .A2(n563), .ZN(n400) );
  XNOR2_X1 U473 ( .A(n400), .B(n399), .ZN(n401) );
  NOR2_X1 U474 ( .A1(n586), .A2(n401), .ZN(n402) );
  NAND2_X1 U475 ( .A1(n402), .A2(n561), .ZN(n403) );
  XNOR2_X1 U476 ( .A(n404), .B(n403), .ZN(n409) );
  XOR2_X1 U477 ( .A(KEYINPUT36), .B(n561), .Z(n589) );
  NAND2_X1 U478 ( .A1(n586), .A2(n589), .ZN(n405) );
  XNOR2_X1 U479 ( .A(KEYINPUT45), .B(n405), .ZN(n407) );
  NAND2_X1 U480 ( .A1(n582), .A2(n563), .ZN(n406) );
  NOR2_X1 U481 ( .A1(n407), .A2(n406), .ZN(n408) );
  NOR2_X1 U482 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U483 ( .A(n410), .B(KEYINPUT48), .ZN(n535) );
  INV_X1 U484 ( .A(n535), .ZN(n411) );
  NAND2_X1 U485 ( .A1(n412), .A2(n411), .ZN(n415) );
  NOR2_X1 U486 ( .A1(n526), .A2(n416), .ZN(n576) );
  XOR2_X1 U487 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n418) );
  XNOR2_X1 U488 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n417) );
  XNOR2_X1 U489 ( .A(n418), .B(n417), .ZN(n424) );
  XOR2_X1 U490 ( .A(KEYINPUT22), .B(G106GAT), .Z(n422) );
  XNOR2_X1 U491 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U492 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U493 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U494 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U495 ( .A(n426), .B(n425), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n427), .B(KEYINPUT87), .ZN(n429) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n436) );
  INV_X1 U498 ( .A(n434), .ZN(n435) );
  NAND2_X1 U499 ( .A1(n576), .A2(n468), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n437), .B(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U501 ( .A(KEYINPUT64), .B(G176GAT), .Z(n439) );
  XNOR2_X1 U502 ( .A(G169GAT), .B(G43GAT), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n445) );
  XOR2_X1 U504 ( .A(G99GAT), .B(G190GAT), .Z(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U507 ( .A(n445), .B(n444), .Z(n449) );
  NAND2_X1 U508 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n450), .B(KEYINPUT20), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U511 ( .A1(n455), .A2(n536), .ZN(n570) );
  NOR2_X1 U512 ( .A1(n561), .A2(n570), .ZN(n458) );
  XOR2_X1 U513 ( .A(n555), .B(KEYINPUT105), .Z(n565) );
  NOR2_X1 U514 ( .A1(n579), .A2(n565), .ZN(n459) );
  XOR2_X1 U515 ( .A(n459), .B(KEYINPUT106), .Z(n514) );
  INV_X1 U516 ( .A(n514), .ZN(n479) );
  NAND2_X1 U517 ( .A1(n536), .A2(n529), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n460), .A2(n468), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT94), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT25), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n536), .A2(n468), .ZN(n463) );
  XNOR2_X1 U522 ( .A(KEYINPUT26), .B(n463), .ZN(n577) );
  XNOR2_X1 U523 ( .A(n529), .B(KEYINPUT27), .ZN(n469) );
  AND2_X1 U524 ( .A1(n577), .A2(n469), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n466), .A2(n526), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT95), .ZN(n474) );
  INV_X1 U528 ( .A(n539), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n469), .A2(n526), .ZN(n470) );
  XOR2_X1 U530 ( .A(KEYINPUT93), .B(n470), .Z(n534) );
  NOR2_X1 U531 ( .A1(n536), .A2(n534), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n493) );
  NAND2_X1 U534 ( .A1(n493), .A2(n571), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(KEYINPUT99), .ZN(n476) );
  NAND2_X1 U536 ( .A1(n476), .A2(n589), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT100), .B(KEYINPUT37), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n486) );
  NAND2_X1 U539 ( .A1(n479), .A2(n486), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n532), .A2(n539), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n482) );
  XNOR2_X1 U542 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1339GAT) );
  NAND2_X1 U544 ( .A1(n579), .A2(n582), .ZN(n495) );
  INV_X1 U545 ( .A(n495), .ZN(n485) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT38), .B(n487), .Z(n510) );
  NAND2_X1 U548 ( .A1(n510), .A2(n536), .ZN(n491) );
  XOR2_X1 U549 ( .A(KEYINPUT102), .B(KEYINPUT40), .Z(n489) );
  INV_X1 U550 ( .A(G43GAT), .ZN(n488) );
  NOR2_X1 U551 ( .A1(n547), .A2(n571), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT16), .ZN(n494) );
  NAND2_X1 U553 ( .A1(n494), .A2(n493), .ZN(n513) );
  NOR2_X1 U554 ( .A1(n495), .A2(n513), .ZN(n503) );
  NAND2_X1 U555 ( .A1(n526), .A2(n503), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(KEYINPUT34), .ZN(n497) );
  XNOR2_X1 U557 ( .A(G1GAT), .B(n497), .ZN(G1324GAT) );
  NAND2_X1 U558 ( .A1(n503), .A2(n529), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n498), .B(KEYINPUT96), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G8GAT), .B(n499), .ZN(G1325GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n501) );
  NAND2_X1 U562 ( .A1(n503), .A2(n536), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U564 ( .A(G15GAT), .B(n502), .Z(G1326GAT) );
  NAND2_X1 U565 ( .A1(n539), .A2(n503), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(KEYINPUT98), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  XOR2_X1 U568 ( .A(G29GAT), .B(KEYINPUT39), .Z(n507) );
  NAND2_X1 U569 ( .A1(n510), .A2(n526), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  XOR2_X1 U571 ( .A(G36GAT), .B(KEYINPUT101), .Z(n509) );
  NAND2_X1 U572 ( .A1(n529), .A2(n510), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1329GAT) );
  XOR2_X1 U574 ( .A(G50GAT), .B(KEYINPUT103), .Z(n512) );
  NAND2_X1 U575 ( .A1(n510), .A2(n539), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(G1331GAT) );
  NOR2_X1 U577 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n526), .A2(n522), .ZN(n518) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n516) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n522), .A2(n529), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n536), .A2(n522), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(KEYINPUT108), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G71GAT), .B(n521), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n524) );
  NAND2_X1 U589 ( .A1(n522), .A2(n539), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U591 ( .A(G78GAT), .B(n525), .Z(G1335GAT) );
  XOR2_X1 U592 ( .A(G85GAT), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U593 ( .A1(n532), .A2(n526), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT112), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n536), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(G99GAT), .ZN(G1338GAT) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n551), .A2(n536), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT116), .B(n537), .ZN(n538) );
  NOR2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n579), .A2(n548), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 U606 ( .A(n548), .ZN(n541) );
  NOR2_X1 U607 ( .A1(n565), .A2(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n545) );
  NAND2_X1 U611 ( .A1(n548), .A2(n586), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n577), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n563), .A2(n560), .ZN(n552) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n555), .A2(n560), .ZN(n556) );
  XOR2_X1 U624 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U625 ( .A1(n571), .A2(n560), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n570), .ZN(n564) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  XNOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n565), .A2(n570), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT59), .B(n575), .Z(n581) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT123), .ZN(n590) );
  NAND2_X1 U645 ( .A1(n590), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U648 ( .A(n582), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n590), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n590), .A2(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT126), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

