//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT0), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT0), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n193), .B(KEYINPUT64), .C1(new_n195), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT0), .B(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(KEYINPUT0), .A3(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n192), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n196), .B2(new_n193), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n190), .A2(new_n192), .A3(new_n206), .A4(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n205), .B1(G125), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G224), .ZN(new_n213));
  XOR2_X1   g027(.A(new_n213), .B(KEYINPUT87), .Z(new_n214));
  XNOR2_X1  g028(.A(new_n211), .B(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G119), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(G113), .B1(new_n218), .B2(KEYINPUT5), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n220));
  INV_X1    g034(.A(G119), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G116), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(KEYINPUT68), .A3(G119), .ZN(new_n223));
  AOI211_X1 g037(.A(KEYINPUT69), .B(new_n217), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n223), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n218), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n219), .B1(new_n228), .B2(KEYINPUT5), .ZN(new_n229));
  INV_X1    g043(.A(G107), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT82), .B1(new_n230), .B2(G104), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(G104), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n230), .A2(KEYINPUT82), .A3(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(G101), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n230), .A2(G104), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n237));
  INV_X1    g051(.A(G104), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G107), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n230), .A2(KEYINPUT3), .A3(G104), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n236), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n226), .A2(new_n218), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT2), .B(G113), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT84), .B1(new_n229), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n246), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n228), .B2(new_n251), .ZN(new_n252));
  OR3_X1    g066(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n242), .ZN(new_n253));
  INV_X1    g067(.A(new_n241), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G101), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT4), .A3(new_n243), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT84), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n235), .A2(new_n243), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(new_n247), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n245), .A2(KEYINPUT69), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n217), .B1(new_n222), .B2(new_n223), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n225), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n261), .A2(KEYINPUT5), .A3(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n258), .B(new_n260), .C1(new_n264), .C2(new_n219), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n250), .A2(new_n257), .A3(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(G110), .B(G122), .Z(new_n267));
  XOR2_X1   g081(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(KEYINPUT85), .A3(new_n267), .ZN(new_n270));
  INV_X1    g084(.A(new_n267), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n250), .A2(new_n257), .A3(new_n265), .A4(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(KEYINPUT6), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT85), .B1(new_n266), .B2(new_n267), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n215), .B(new_n269), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n213), .A2(KEYINPUT7), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n211), .B(new_n277), .Z(new_n278));
  OAI21_X1  g092(.A(new_n259), .B1(new_n229), .B2(new_n247), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n282), .B(KEYINPUT88), .Z(new_n283));
  OAI21_X1  g097(.A(new_n260), .B1(new_n283), .B2(new_n219), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n280), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n267), .B(KEYINPUT8), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n272), .B(new_n278), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n275), .A2(new_n276), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G210), .B1(G237), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n275), .A2(new_n288), .A3(new_n276), .A4(new_n290), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n188), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G125), .ZN(new_n295));
  OAI21_X1  g109(.A(G140), .B1(new_n295), .B2(KEYINPUT77), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(G125), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n299), .A3(KEYINPUT16), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT16), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n298), .A4(G125), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n298), .A3(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT78), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n189), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n300), .A2(G146), .A3(new_n303), .A4(new_n305), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT24), .B(G110), .Z(new_n310));
  XNOR2_X1  g124(.A(G119), .B(G128), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n221), .B2(G128), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n221), .A2(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G110), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(KEYINPUT76), .A3(G110), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n309), .A2(new_n312), .A3(new_n322), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n317), .A2(G110), .B1(new_n310), .B2(new_n311), .ZN(new_n324));
  XNOR2_X1  g138(.A(G125), .B(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n189), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n308), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n212), .A2(G221), .A3(G234), .ZN(new_n330));
  XOR2_X1   g144(.A(new_n329), .B(new_n330), .Z(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n323), .A2(new_n327), .A3(new_n331), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n276), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT79), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n333), .A2(new_n338), .A3(new_n276), .A4(new_n334), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n335), .A2(new_n337), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n336), .A2(KEYINPUT80), .A3(new_n337), .A4(new_n339), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(G234), .B2(new_n276), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n333), .A2(new_n334), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n347), .A2(G902), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n345), .A2(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G469), .ZN(new_n352));
  INV_X1    g166(.A(new_n204), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n256), .A2(new_n353), .A3(new_n253), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n209), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n200), .A2(KEYINPUT83), .A3(new_n206), .A4(G128), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n208), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n355), .B1(new_n359), .B2(new_n259), .ZN(new_n360));
  INV_X1    g174(.A(G137), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT11), .A3(G134), .ZN(new_n362));
  INV_X1    g176(.A(G134), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G137), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT11), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT65), .B(new_n366), .C1(new_n363), .C2(G137), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n361), .A2(G134), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT65), .B1(new_n369), .B2(new_n366), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n365), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G131), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT66), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n362), .A2(new_n364), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n363), .A2(G137), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(KEYINPUT11), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n378), .B2(new_n367), .ZN(new_n379));
  INV_X1    g193(.A(new_n373), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n244), .A2(KEYINPUT10), .A3(new_n210), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n354), .A2(new_n360), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G110), .B(G140), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT81), .ZN(new_n387));
  INV_X1    g201(.A(G227), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G953), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n387), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n359), .A2(new_n259), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n244), .A2(new_n210), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT12), .B(new_n382), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n382), .B1(new_n392), .B2(new_n393), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n391), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n354), .A2(new_n360), .A3(new_n384), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n382), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n390), .B1(new_n400), .B2(new_n385), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n352), .B(new_n276), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(G469), .A2(G902), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n385), .A3(new_n390), .ZN(new_n404));
  INV_X1    g218(.A(new_n399), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n397), .A2(new_n394), .B1(new_n405), .B2(new_n383), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n404), .B(G469), .C1(new_n406), .C2(new_n390), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G221), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT9), .B(G234), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(new_n276), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n294), .A2(new_n351), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT91), .B(G104), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n296), .A2(new_n299), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT19), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(KEYINPUT19), .B2(new_n325), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n189), .ZN(new_n422));
  INV_X1    g236(.A(G237), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n212), .A3(G214), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(new_n191), .ZN(new_n425));
  NOR2_X1   g239(.A1(G237), .A2(G953), .ZN(new_n426));
  AOI21_X1  g240(.A(G143), .B1(new_n426), .B2(G214), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n372), .ZN(new_n429));
  OAI21_X1  g243(.A(G131), .B1(new_n425), .B2(new_n427), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n422), .A2(new_n308), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(KEYINPUT18), .A2(G131), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n428), .B(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n326), .B1(new_n419), .B2(new_n189), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT90), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n435), .A2(KEYINPUT90), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n418), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT17), .B(G131), .C1(new_n425), .C2(new_n427), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n307), .A2(new_n308), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT92), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT17), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n429), .A2(new_n444), .A3(new_n430), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n307), .A2(KEYINPUT92), .A3(new_n308), .A4(new_n440), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n437), .A2(new_n436), .ZN(new_n448));
  INV_X1    g262(.A(new_n434), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n418), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n439), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G475), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n276), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT93), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n451), .B1(new_n447), .B2(new_n450), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n276), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G475), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n453), .A2(new_n462), .A3(new_n454), .A4(new_n276), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n464));
  AOI21_X1  g278(.A(G475), .B1(new_n439), .B2(new_n452), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(new_n465), .B2(new_n276), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n457), .B(new_n461), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n410), .A2(new_n346), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n216), .A2(G122), .ZN(new_n470));
  INV_X1    g284(.A(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G116), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n472), .A3(new_n230), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n191), .A2(G128), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n196), .A2(G143), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n363), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n476), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G134), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT95), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n216), .B2(G122), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n216), .A2(G122), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n471), .A2(G116), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n482), .ZN(new_n487));
  OAI211_X1 g301(.A(KEYINPUT95), .B(new_n472), .C1(new_n486), .C2(new_n482), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI221_X4 g303(.A(new_n474), .B1(new_n478), .B2(new_n480), .C1(new_n489), .C2(G107), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n478), .A2(KEYINPUT94), .ZN(new_n491));
  OAI21_X1  g305(.A(G107), .B1(new_n486), .B2(new_n484), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n473), .ZN(new_n493));
  OR3_X1    g307(.A1(new_n479), .A2(KEYINPUT94), .A3(G134), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT13), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n191), .A3(G128), .ZN(new_n496));
  OAI211_X1 g310(.A(G134), .B(new_n496), .C1(new_n479), .C2(new_n495), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n469), .B1(new_n490), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n489), .A2(G107), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n478), .A2(new_n480), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(new_n473), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n498), .A3(new_n468), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n276), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT96), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n506), .B(new_n512), .Z(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n467), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(G472), .A2(G902), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n261), .A2(new_n263), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n247), .B1(new_n517), .B2(new_n246), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n365), .B(new_n372), .C1(new_n368), .C2(new_n370), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n364), .A2(new_n369), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G131), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(KEYINPUT67), .A3(new_n521), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n210), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n382), .A2(new_n353), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n210), .A2(new_n521), .A3(new_n519), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n204), .B1(new_n374), .B2(new_n381), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT30), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n518), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n518), .A3(new_n530), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n426), .A2(G210), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n242), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n534), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT74), .B1(new_n531), .B2(new_n532), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n528), .A2(new_n545), .A3(new_n530), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n546), .A3(new_n518), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n519), .A2(KEYINPUT67), .A3(new_n521), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT67), .B1(new_n519), .B2(new_n521), .ZN(new_n551));
  INV_X1    g365(.A(new_n210), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n252), .B1(new_n553), .B2(new_n532), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n526), .A2(new_n528), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT73), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n252), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n535), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n549), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n540), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n543), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT70), .B1(new_n541), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n529), .A2(new_n533), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n252), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n535), .A3(new_n562), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT31), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n516), .B1(new_n563), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT32), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT32), .B(new_n516), .C1(new_n563), .C2(new_n571), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n562), .B1(new_n567), .B2(new_n535), .ZN(new_n576));
  AOI211_X1 g390(.A(KEYINPUT29), .B(new_n576), .C1(new_n561), .C2(new_n562), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n547), .A2(new_n548), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n252), .B1(new_n531), .B2(new_n532), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n535), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n580), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT75), .B1(new_n580), .B2(KEYINPUT28), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n562), .A2(KEYINPUT29), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n276), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G472), .B1(new_n577), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n574), .A2(new_n575), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n212), .A2(G952), .ZN(new_n588));
  NAND2_X1  g402(.A1(G234), .A2(G237), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT21), .B(G898), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(G902), .A3(G953), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n591), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n415), .A2(new_n515), .A3(new_n587), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NAND2_X1  g413(.A1(new_n345), .A2(new_n347), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n349), .A2(new_n350), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n414), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n276), .B1(new_n563), .B2(new_n571), .ZN(new_n603));
  INV_X1    g417(.A(new_n560), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n557), .B1(new_n556), .B2(new_n252), .ZN(new_n605));
  AOI211_X1 g419(.A(KEYINPUT73), .B(new_n518), .C1(new_n526), .C2(new_n528), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n607), .B2(new_n535), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n540), .B1(new_n608), .B2(new_n549), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n609), .A2(new_n543), .A3(new_n565), .A4(new_n570), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n603), .A2(G472), .B1(new_n610), .B2(new_n516), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n602), .A2(new_n611), .A3(KEYINPUT97), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT97), .B1(new_n602), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI211_X1 g428(.A(new_n188), .B(new_n596), .C1(new_n292), .C2(new_n293), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n505), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n507), .A2(G902), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n505), .B2(KEYINPUT98), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n503), .A2(new_n498), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT98), .B1(new_n621), .B2(new_n469), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n619), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n500), .B2(new_n504), .ZN(new_n626));
  NOR4_X1   g440(.A1(new_n626), .A2(new_n622), .A3(KEYINPUT99), .A4(new_n616), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n617), .B(new_n618), .C1(new_n624), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n506), .A2(new_n507), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n467), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n615), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n614), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NOR2_X1   g451(.A1(new_n467), .A2(new_n513), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n615), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n614), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NAND2_X1  g456(.A1(new_n408), .A2(new_n413), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n328), .B(KEYINPUT100), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n332), .A2(KEYINPUT36), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n644), .B(new_n645), .Z(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n350), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n643), .B1(new_n600), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n615), .A2(new_n515), .A3(new_n611), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  OAI21_X1  g465(.A(new_n590), .B1(G900), .B2(new_n594), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n638), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n587), .A2(new_n294), .A3(new_n648), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  XNOR2_X1  g469(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n652), .B(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n643), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT40), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n467), .A2(new_n514), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n659), .A2(new_n187), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n580), .A2(new_n540), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n568), .A2(G472), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(G472), .A2(G902), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(KEYINPUT101), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(KEYINPUT101), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n574), .A2(new_n575), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n600), .A2(new_n647), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n292), .A2(new_n293), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT38), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n661), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  AND3_X1   g489(.A1(new_n630), .A2(new_n467), .A3(new_n652), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n672), .A2(new_n676), .A3(new_n187), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n294), .A2(KEYINPUT103), .A3(new_n676), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n587), .A3(new_n648), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  NAND2_X1  g496(.A1(new_n587), .A2(new_n351), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n276), .B1(new_n398), .B2(new_n401), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n413), .A3(new_n402), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n683), .A2(new_n633), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT41), .B(G113), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  INV_X1    g503(.A(new_n683), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n691));
  INV_X1    g505(.A(new_n686), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n690), .A2(new_n639), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n587), .A2(new_n615), .A3(new_n351), .A4(new_n638), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT104), .B1(new_n694), .B2(new_n686), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  NAND3_X1  g511(.A1(new_n587), .A2(new_n515), .A3(new_n597), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n188), .B(new_n686), .C1(new_n292), .C2(new_n293), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n669), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n221), .ZN(G21));
  NAND2_X1  g516(.A1(new_n603), .A2(G472), .ZN(new_n703));
  AOI22_X1  g517(.A1(new_n583), .A2(new_n540), .B1(KEYINPUT31), .B2(new_n568), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n543), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n516), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n351), .A2(new_n703), .A3(new_n597), .A4(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n294), .A2(new_n660), .A3(new_n692), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  AOI22_X1  g524(.A1(new_n603), .A2(G472), .B1(new_n516), .B2(new_n705), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n699), .A2(new_n669), .A3(new_n711), .A4(new_n676), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT32), .B1(new_n610), .B2(new_n516), .ZN(new_n715));
  INV_X1    g529(.A(new_n575), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n575), .A2(KEYINPUT105), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n586), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n676), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n414), .A2(new_n292), .A3(new_n187), .A4(new_n293), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n719), .A2(new_n351), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n721), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n587), .A2(new_n725), .A3(new_n351), .A4(new_n676), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n722), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NAND4_X1  g543(.A1(new_n690), .A2(KEYINPUT106), .A3(new_n653), .A4(new_n725), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n587), .A2(new_n725), .A3(new_n351), .A4(new_n653), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  NAND2_X1  g549(.A1(new_n703), .A2(new_n572), .ZN(new_n736));
  INV_X1    g550(.A(new_n467), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n630), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(new_n740), .A3(new_n630), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n736), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT44), .B1(new_n742), .B2(new_n669), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n739), .A2(new_n741), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT44), .A3(new_n736), .A4(new_n669), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n672), .A2(new_n188), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n742), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n669), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT108), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n747), .A2(new_n752), .A3(new_n749), .A4(new_n748), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n743), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n404), .B1(new_n406), .B2(new_n390), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT45), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(G469), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT46), .B1(new_n757), .B2(new_n403), .ZN(new_n758));
  INV_X1    g572(.A(new_n402), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n403), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n412), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n657), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n754), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  OR2_X1    g580(.A1(new_n762), .A2(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n762), .A2(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n587), .A2(new_n351), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n720), .A2(new_n188), .A3(new_n672), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  AND4_X1   g587(.A1(new_n351), .A2(new_n744), .A3(new_n591), .A4(new_n711), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n188), .B1(KEYINPUT113), .B2(KEYINPUT50), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n673), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n692), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n774), .A2(new_n692), .A3(new_n778), .A4(new_n776), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n591), .A2(new_n744), .A3(new_n692), .A4(new_n748), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n669), .A3(new_n711), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n748), .A2(new_n351), .A3(new_n692), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n590), .A3(new_n668), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n737), .A3(new_n629), .A4(new_n628), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n780), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n685), .A2(new_n402), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n412), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n767), .A2(new_n768), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n767), .A2(KEYINPUT115), .A3(new_n768), .A4(new_n790), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n774), .A2(new_n748), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n788), .A2(new_n796), .A3(KEYINPUT51), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n788), .A2(new_n796), .A3(KEYINPUT116), .A4(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n791), .A2(new_n795), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n787), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT114), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n719), .A2(new_n351), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n782), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT48), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n774), .A2(new_n294), .A3(new_n692), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(KEYINPUT117), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n809), .A2(KEYINPUT117), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n808), .B(new_n588), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n804), .B2(KEYINPUT114), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n801), .A2(new_n805), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n785), .A2(new_n632), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n587), .A2(new_n515), .A3(new_n648), .A4(new_n652), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n711), .A2(new_n648), .A3(new_n676), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n748), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n734), .A2(new_n728), .A3(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n414), .A2(new_n672), .A3(new_n187), .A4(new_n660), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n670), .A3(new_n652), .A4(new_n668), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n681), .A2(new_n822), .A3(new_n654), .A4(new_n712), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n414), .A2(new_n294), .A3(new_n652), .A4(new_n660), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n671), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n654), .A3(new_n681), .A4(new_n712), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n598), .A2(new_n649), .A3(new_n709), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT109), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n737), .A2(new_n831), .A3(new_n514), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT109), .B1(new_n467), .B2(new_n513), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n631), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n615), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n612), .A2(new_n613), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n830), .A2(new_n836), .A3(new_n687), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n701), .B1(new_n693), .B2(new_n695), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n820), .A2(new_n829), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  OR3_X1    g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n654), .A2(new_n712), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT110), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n681), .A3(new_n827), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n825), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n837), .A2(new_n838), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n820), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n841), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n733), .A2(new_n730), .B1(new_n724), .B2(new_n727), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n837), .A2(new_n854), .A3(new_n819), .A4(new_n838), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n825), .A2(new_n828), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n853), .B(new_n841), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n853), .B1(new_n839), .B2(new_n841), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n846), .A2(KEYINPUT53), .A3(new_n820), .A4(new_n847), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n814), .A2(new_n815), .A3(new_n852), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(G952), .B2(G953), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n789), .B(KEYINPUT49), .Z(new_n866));
  NOR3_X1   g680(.A1(new_n673), .A2(new_n738), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n351), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n668), .A2(new_n868), .A3(new_n188), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n413), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n870), .ZN(G75));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n841), .B1(new_n855), .B2(new_n856), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT112), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n862), .A3(new_n857), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(G902), .ZN(new_n876));
  INV_X1    g690(.A(G210), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(new_n215), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT118), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(KEYINPUT119), .B2(new_n872), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n878), .A2(new_n883), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n212), .A2(G952), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G51));
  XNOR2_X1  g701(.A(new_n875), .B(new_n861), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n403), .B(KEYINPUT57), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n888), .A2(new_n889), .B1(new_n401), .B2(new_n398), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n875), .A2(G469), .A3(G902), .A4(new_n756), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT120), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n890), .B2(new_n892), .ZN(G54));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n876), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n453), .B1(new_n895), .B2(G475), .ZN(new_n896));
  INV_X1    g710(.A(new_n453), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n876), .A2(new_n894), .A3(new_n454), .A4(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n886), .A3(new_n898), .ZN(G60));
  INV_X1    g713(.A(new_n886), .ZN(new_n900));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT59), .Z(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n852), .B2(new_n863), .ZN(new_n903));
  INV_X1    g717(.A(new_n624), .ZN(new_n904));
  INV_X1    g718(.A(new_n627), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n904), .A2(new_n905), .B1(new_n616), .B2(new_n505), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n900), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n906), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n888), .A2(new_n908), .A3(new_n902), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT60), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n875), .A2(new_n646), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n860), .B2(new_n862), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n900), .B(new_n914), .C1(new_n915), .C2(new_n349), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT121), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(KEYINPUT121), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n875), .A2(new_n913), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n886), .B1(new_n921), .B2(new_n348), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(KEYINPUT121), .A3(new_n917), .A4(new_n914), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n920), .A2(new_n923), .ZN(G66));
  INV_X1    g738(.A(G224), .ZN(new_n925));
  OAI21_X1  g739(.A(G953), .B1(new_n593), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n847), .B2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n879), .B1(G898), .B2(new_n212), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT122), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n927), .B(new_n929), .ZN(G69));
  INV_X1    g744(.A(G900), .ZN(new_n931));
  OAI21_X1  g745(.A(G953), .B1(new_n388), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n566), .B(new_n421), .ZN(new_n933));
  AND4_X1   g747(.A1(new_n763), .A2(new_n690), .A3(new_n725), .A4(new_n834), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n844), .A2(new_n674), .A3(new_n681), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n844), .A2(KEYINPUT62), .A3(new_n674), .A4(new_n681), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n772), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n754), .B2(new_n764), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n941), .A3(KEYINPUT124), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT124), .B1(new_n939), .B2(new_n941), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n212), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n933), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n764), .A2(new_n806), .A3(new_n294), .A4(new_n660), .ZN(new_n948));
  AND4_X1   g762(.A1(new_n681), .A2(new_n948), .A3(new_n844), .A4(new_n854), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n212), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n931), .A2(G953), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT125), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n933), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n945), .B2(KEYINPUT123), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n932), .B1(new_n947), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n955), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n939), .A2(new_n941), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(G953), .B1(new_n961), .B2(new_n942), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n958), .B1(new_n962), .B2(new_n946), .ZN(new_n963));
  INV_X1    g777(.A(new_n933), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n962), .B2(KEYINPUT123), .ZN(new_n965));
  INV_X1    g779(.A(new_n932), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n957), .A2(new_n967), .ZN(G72));
  NAND3_X1  g782(.A1(new_n961), .A2(new_n847), .A3(new_n942), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n664), .B(KEYINPUT63), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n534), .A2(new_n536), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(new_n540), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n941), .A2(new_n847), .A3(new_n949), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n971), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n534), .A2(new_n536), .A3(new_n562), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n886), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n541), .A2(KEYINPUT126), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n576), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n851), .A2(new_n971), .A3(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n975), .A2(KEYINPUT127), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n984));
  INV_X1    g798(.A(new_n974), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n969), .B2(new_n971), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n979), .A2(new_n982), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n983), .A2(new_n988), .ZN(G57));
endmodule


