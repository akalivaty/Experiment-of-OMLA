//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT73), .Z(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT10), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G104), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G107), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT74), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT3), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(new_n194), .A3(KEYINPUT3), .A4(G104), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n196), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(new_n194), .A3(G104), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n201), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT75), .A3(new_n196), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(G128), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(G143), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n218), .A2(G143), .ZN(new_n221));
  OAI22_X1  g035(.A1(new_n219), .A2(new_n220), .B1(new_n213), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT78), .B1(new_n194), .B2(G104), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT77), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n197), .B2(G107), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT78), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n197), .A3(G107), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n194), .A2(KEYINPUT77), .A3(G104), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n223), .A2(new_n225), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n217), .A2(new_n222), .B1(new_n229), .B2(G101), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT79), .B1(new_n211), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT75), .B1(new_n209), .B2(new_n196), .ZN(new_n232));
  AOI211_X1 g046(.A(new_n204), .B(new_n195), .C1(new_n208), .C2(new_n201), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n230), .B(KEYINPUT79), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n192), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G137), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(KEYINPUT65), .B(new_n237), .C1(new_n238), .C2(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n238), .A2(G137), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n238), .A2(G137), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(KEYINPUT11), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n243), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n247), .B1(new_n243), .B2(new_n246), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n208), .A2(new_n201), .B1(new_n197), .B2(G107), .ZN(new_n251));
  OAI221_X1 g065(.A(KEYINPUT4), .B1(new_n193), .B2(new_n251), .C1(new_n232), .C2(new_n233), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n213), .A2(new_n221), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT64), .B1(new_n212), .B2(G146), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n213), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n255), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n251), .A2(new_n193), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n205), .A2(new_n210), .B1(G101), .B2(new_n229), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n215), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n214), .B1(new_n269), .B2(new_n256), .ZN(new_n270));
  OAI21_X1  g084(.A(G128), .B1(new_n213), .B2(new_n216), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n192), .B1(new_n272), .B2(new_n217), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n252), .A2(new_n266), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n236), .A2(new_n250), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT80), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n236), .A2(new_n277), .A3(new_n274), .A4(new_n250), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G110), .B(G140), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n281), .A2(G227), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n280), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n285));
  NAND2_X1  g099(.A1(new_n272), .A2(new_n217), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n267), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n287), .A2(new_n288), .B1(new_n291), .B2(new_n234), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n285), .B1(new_n292), .B2(new_n250), .ZN(new_n293));
  INV_X1    g107(.A(new_n250), .ZN(new_n294));
  NOR2_X1   g108(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n231), .A2(new_n235), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n267), .A2(new_n286), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n294), .B(new_n295), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n279), .A2(new_n284), .A3(new_n293), .A4(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n274), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT10), .B1(new_n291), .B2(new_n234), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT82), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n236), .A2(new_n303), .A3(new_n274), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n304), .A3(new_n294), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n284), .B1(new_n279), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT83), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI211_X1 g122(.A(KEYINPUT83), .B(new_n284), .C1(new_n279), .C2(new_n305), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n190), .B(new_n191), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n279), .A2(new_n305), .A3(new_n284), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n293), .A2(new_n298), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n278), .B2(new_n276), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n311), .B(G469), .C1(new_n313), .C2(new_n284), .ZN(new_n314));
  NAND2_X1  g128(.A1(G469), .A2(G902), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n189), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G478), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT15), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT94), .ZN(new_n320));
  INV_X1    g134(.A(G217), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n187), .A2(new_n321), .A3(G953), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT91), .ZN(new_n324));
  XNOR2_X1  g138(.A(G128), .B(G143), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n238), .ZN(new_n326));
  INV_X1    g140(.A(G122), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G116), .ZN(new_n328));
  INV_X1    g142(.A(G116), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G122), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G107), .ZN(new_n332));
  XNOR2_X1  g146(.A(G116), .B(G122), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(new_n194), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n326), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT13), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n220), .B2(G143), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n212), .A2(KEYINPUT13), .A3(G128), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n337), .B(new_n338), .C1(G128), .C2(new_n212), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(G134), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n324), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n331), .A2(G107), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n333), .A2(new_n194), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n342), .A2(new_n343), .B1(new_n325), .B2(new_n238), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(G134), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(KEYINPUT91), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n343), .B(KEYINPUT92), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n325), .B(new_n238), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n329), .A2(KEYINPUT14), .A3(G122), .ZN(new_n351));
  OAI211_X1 g165(.A(G107), .B(new_n351), .C1(new_n331), .C2(KEYINPUT14), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n347), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n348), .B1(new_n347), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n323), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n346), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT91), .B1(new_n344), .B2(new_n345), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT93), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n347), .A2(new_n348), .A3(new_n353), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n322), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n320), .B1(new_n363), .B2(new_n191), .ZN(new_n364));
  AOI211_X1 g178(.A(KEYINPUT94), .B(G902), .C1(new_n356), .C2(new_n362), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n319), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n354), .A2(new_n355), .A3(new_n323), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n322), .B1(new_n360), .B2(new_n361), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n191), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT94), .ZN(new_n370));
  INV_X1    g184(.A(new_n319), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G140), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G125), .ZN(new_n375));
  INV_X1    g189(.A(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G140), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n375), .A2(new_n377), .A3(new_n218), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n218), .B1(new_n375), .B2(new_n377), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT88), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(new_n377), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G146), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n375), .A2(new_n377), .A3(new_n218), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G237), .ZN(new_n388));
  INV_X1    g202(.A(G237), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(KEYINPUT68), .ZN(new_n390));
  OAI211_X1 g204(.A(G214), .B(new_n281), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n212), .A2(KEYINPUT87), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(KEYINPUT68), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n387), .A2(G237), .ZN(new_n396));
  AOI21_X1  g210(.A(G953), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(G214), .A3(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT18), .A2(G131), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n386), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n402));
  AOI211_X1 g216(.A(new_n402), .B(new_n247), .C1(new_n394), .C2(new_n398), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT89), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n391), .A2(new_n393), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n392), .B1(new_n397), .B2(G214), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT18), .B(G131), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n386), .A4(new_n400), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G113), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n197), .ZN(new_n412));
  OAI21_X1  g226(.A(G131), .B1(new_n405), .B2(new_n406), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT17), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n394), .A2(new_n247), .A3(new_n398), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G125), .B(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT16), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n375), .A2(KEYINPUT16), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(G146), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT71), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n419), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT72), .B1(new_n423), .B2(new_n218), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT72), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n425), .B(G146), .C1(new_n418), .C2(new_n419), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(KEYINPUT17), .B(G131), .C1(new_n405), .C2(new_n406), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n416), .A2(new_n422), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n410), .A2(new_n412), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n412), .B1(new_n410), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n191), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G475), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n281), .A2(G952), .ZN(new_n434));
  NAND2_X1  g248(.A1(G234), .A2(G237), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(G898), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(G902), .A3(G953), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n420), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT90), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n381), .B1(new_n444), .B2(KEYINPUT19), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n381), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n443), .B1(new_n447), .B2(new_n218), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n413), .A2(new_n415), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n386), .A2(new_n400), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n408), .B1(new_n451), .B2(new_n407), .ZN(new_n452));
  AND4_X1   g266(.A1(new_n408), .A2(new_n407), .A3(new_n386), .A4(new_n400), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n412), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n412), .B(new_n429), .C1(new_n452), .C2(new_n453), .ZN(new_n457));
  AOI211_X1 g271(.A(KEYINPUT20), .B(new_n442), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n404), .A2(new_n409), .B1(new_n449), .B2(new_n448), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n412), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n461), .B2(new_n441), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n433), .B(new_n440), .C1(new_n458), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n373), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G214), .B1(G237), .B2(G902), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT84), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n287), .A2(new_n376), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n263), .A2(G125), .ZN(new_n472));
  INV_X1    g286(.A(G224), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT7), .B1(new_n473), .B2(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n471), .A2(KEYINPUT85), .A3(new_n472), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n471), .A2(new_n472), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n474), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT5), .ZN(new_n483));
  INV_X1    g297(.A(G119), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(G116), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n329), .B2(G119), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(KEYINPUT67), .A3(G116), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n329), .A2(G119), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(G113), .B(new_n485), .C1(new_n490), .C2(new_n483), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT2), .B(G113), .Z(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n267), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT8), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n490), .B(new_n492), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n264), .B2(new_n265), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n252), .A2(new_n499), .B1(new_n267), .B2(new_n494), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n495), .A2(new_n497), .B1(new_n500), .B2(new_n496), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n482), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n252), .A2(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n267), .A2(new_n494), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n496), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n496), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(KEYINPUT6), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n473), .A2(G953), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n480), .B(new_n510), .ZN(new_n511));
  OR3_X1    g325(.A1(new_n500), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n470), .B1(new_n502), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n502), .A2(new_n513), .A3(new_n470), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n466), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n464), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n317), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT29), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n243), .A2(new_n246), .A3(new_n247), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n244), .B2(new_n245), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n286), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n270), .A2(new_n261), .B1(new_n253), .B2(new_n254), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n248), .B2(new_n249), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n525), .A3(new_n498), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT28), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n286), .A2(new_n521), .A3(new_n522), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT66), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT66), .B(new_n524), .C1(new_n248), .C2(new_n249), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n528), .B(new_n530), .C1(new_n498), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n397), .A2(G210), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(G101), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n520), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n498), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT30), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n544), .C1(new_n535), .C2(KEYINPUT30), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n526), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n542), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n523), .A2(new_n525), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n543), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n526), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(KEYINPUT69), .A3(new_n543), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n530), .B1(new_n553), .B2(new_n529), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n540), .A2(KEYINPUT29), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n191), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G472), .B1(new_n547), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n545), .A2(new_n540), .A3(new_n526), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT31), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n536), .A2(new_n541), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT31), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n545), .A2(new_n561), .A3(new_n540), .A4(new_n526), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT32), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n557), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n321), .B1(G234), .B2(new_n191), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT22), .B(G137), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n422), .A2(new_n427), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT23), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n484), .B2(G128), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n220), .A2(KEYINPUT23), .A3(G119), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n577), .B(new_n578), .C1(G119), .C2(new_n220), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G110), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(KEYINPUT70), .A3(G110), .ZN(new_n583));
  XNOR2_X1  g397(.A(G119), .B(G128), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT24), .B(G110), .Z(new_n585));
  AOI22_X1  g399(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n575), .A2(new_n586), .ZN(new_n587));
  OAI22_X1  g401(.A1(new_n579), .A2(G110), .B1(new_n584), .B2(new_n585), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n420), .A3(new_n384), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n574), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n589), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n573), .B(new_n591), .C1(new_n575), .C2(new_n586), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT25), .B1(new_n593), .B2(new_n191), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  NOR4_X1   g409(.A1(new_n590), .A2(new_n592), .A3(new_n595), .A4(G902), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n570), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n570), .A2(G902), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n569), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n519), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n193), .ZN(G3));
  NAND2_X1  g418(.A1(new_n310), .A2(new_n316), .ZN(new_n605));
  INV_X1    g419(.A(new_n189), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n563), .A2(new_n565), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n563), .B2(new_n191), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n608), .A2(new_n610), .A3(new_n600), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT95), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n317), .A2(new_n614), .A3(new_n611), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n502), .A2(new_n513), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n467), .A2(KEYINPUT96), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n467), .A2(KEYINPUT96), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n502), .A2(new_n513), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n619), .A2(new_n465), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT97), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n619), .A2(new_n625), .A3(new_n465), .A4(new_n622), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n433), .B1(new_n458), .B2(new_n462), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n367), .B2(new_n368), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n356), .A2(KEYINPUT33), .A3(new_n362), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n318), .A2(G902), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT98), .B(G478), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n369), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n628), .A2(new_n637), .A3(new_n440), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n616), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND3_X1  g457(.A1(new_n363), .A2(new_n320), .A3(new_n191), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n371), .B1(new_n370), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n364), .A2(new_n319), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT99), .B1(new_n647), .B2(new_n463), .ZN(new_n648));
  INV_X1    g462(.A(new_n628), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n373), .A2(new_n649), .A3(new_n650), .A4(new_n440), .ZN(new_n651));
  AND4_X1   g465(.A1(new_n626), .A2(new_n648), .A3(new_n651), .A4(new_n624), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n616), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT100), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT35), .B(G107), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  INV_X1    g470(.A(new_n610), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n607), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n587), .A2(new_n589), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n659), .B(new_n660), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n598), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n597), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n519), .A2(new_n658), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n607), .A2(KEYINPUT32), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n566), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n664), .B1(new_n669), .B2(new_n557), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n317), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n436), .B1(G900), .B2(new_n439), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n433), .B(new_n672), .C1(new_n458), .C2(new_n462), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n647), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n671), .A2(new_n627), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n220), .ZN(G30));
  INV_X1    g490(.A(new_n317), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n672), .B(KEYINPUT39), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OR3_X1    g493(.A1(new_n677), .A2(KEYINPUT40), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT40), .B1(new_n677), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n553), .A2(new_n541), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n191), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n541), .B1(new_n545), .B2(new_n526), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n669), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n663), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n515), .A2(new_n516), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n465), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n691), .A2(new_n692), .A3(new_n649), .A4(new_n647), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n680), .A2(new_n681), .A3(new_n688), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND3_X1  g509(.A1(new_n628), .A2(new_n637), .A3(new_n672), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n628), .A2(new_n637), .A3(KEYINPUT102), .A4(new_n672), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n671), .A2(new_n627), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  OAI21_X1  g515(.A(new_n191), .B1(new_n308), .B2(new_n309), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G469), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n606), .A3(new_n310), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n602), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n703), .A2(KEYINPUT103), .A3(new_n606), .A4(new_n310), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n640), .A2(new_n706), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n706), .A2(new_n707), .A3(new_n652), .A4(new_n708), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n329), .ZN(G18));
  AND3_X1   g529(.A1(new_n569), .A2(new_n464), .A3(new_n663), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n706), .A2(new_n716), .A3(new_n627), .A4(new_n708), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  NOR2_X1   g532(.A1(new_n647), .A2(new_n649), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n624), .A3(new_n440), .A4(new_n626), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n554), .A2(new_n541), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n559), .A3(new_n562), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n565), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n657), .A2(new_n601), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n706), .A2(new_n725), .A3(new_n708), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  AND2_X1   g541(.A1(new_n706), .A2(new_n708), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n698), .A2(new_n699), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n657), .A2(new_n663), .A3(new_n723), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n698), .A2(KEYINPUT105), .A3(new_n699), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n728), .A2(KEYINPUT106), .A3(new_n627), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n706), .A2(new_n627), .A3(new_n708), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n698), .A2(KEYINPUT105), .A3(new_n699), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT105), .B1(new_n698), .B2(new_n699), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n732), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n736), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n731), .A2(new_n733), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT107), .B1(new_n313), .B2(new_n284), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n276), .A2(new_n278), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n748), .B(new_n283), .C1(new_n749), .C2(new_n312), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n747), .A2(new_n750), .A3(G469), .A4(new_n311), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n310), .A2(new_n315), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n689), .A2(new_n189), .A3(new_n692), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n569), .A3(new_n601), .A4(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n745), .B1(new_n746), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n516), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n756), .A2(new_n514), .A3(new_n692), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n606), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n751), .A2(new_n315), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n759), .B2(new_n310), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n707), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n755), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n707), .A3(new_n674), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  OAI21_X1  g579(.A(new_n283), .B1(new_n749), .B2(new_n312), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT45), .B1(new_n766), .B2(new_n311), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n190), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n747), .A2(new_n750), .A3(KEYINPUT45), .A4(new_n311), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n768), .A2(new_n769), .B1(G469), .B2(G902), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT108), .B1(new_n771), .B2(new_n310), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(KEYINPUT108), .A3(new_n310), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n773), .B(new_n774), .C1(KEYINPUT46), .C2(new_n770), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n606), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n776), .A2(KEYINPUT109), .A3(new_n679), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT109), .B1(new_n776), .B2(new_n679), .ZN(new_n778));
  INV_X1    g592(.A(new_n637), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n628), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT43), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n658), .A3(new_n663), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  INV_X1    g599(.A(new_n757), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n777), .A2(new_n778), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  XOR2_X1   g603(.A(new_n776), .B(KEYINPUT47), .Z(new_n790));
  NOR4_X1   g604(.A1(new_n729), .A2(new_n569), .A3(new_n601), .A4(new_n786), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND2_X1  g607(.A1(new_n728), .A2(new_n757), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n794), .A2(new_n600), .A3(new_n436), .A4(new_n686), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n649), .A2(new_n779), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n436), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n781), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n724), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n797), .B(new_n434), .C1(new_n737), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n794), .A2(new_n799), .ZN(new_n803));
  AND4_X1   g617(.A1(KEYINPUT118), .A2(new_n803), .A3(KEYINPUT48), .A4(new_n707), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n803), .B2(new_n707), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n703), .A2(new_n310), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n790), .B1(new_n189), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n786), .A3(new_n801), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n465), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n728), .A2(new_n691), .A3(new_n800), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n812), .A2(new_n813), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n815), .B(new_n816), .Z(new_n817));
  NAND2_X1  g631(.A1(new_n803), .A2(new_n732), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n795), .A2(new_n649), .A3(new_n779), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(KEYINPUT51), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n811), .A2(new_n820), .ZN(new_n824));
  OAI221_X1 g638(.A(new_n807), .B1(new_n811), .B2(new_n823), .C1(new_n824), .C2(KEYINPUT51), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  INV_X1    g640(.A(new_n673), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT112), .B1(new_n645), .B2(new_n646), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n366), .A2(new_n372), .A3(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n827), .A2(new_n757), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n734), .A2(new_n760), .B1(new_n671), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n762), .A2(new_n832), .A3(new_n764), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n709), .A2(new_n717), .A3(new_n726), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n714), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n466), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n689), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(KEYINPUT111), .A3(new_n638), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n639), .B2(new_n517), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n613), .A2(new_n615), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n828), .A2(new_n830), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n517), .A2(new_n440), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n844), .A3(new_n628), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n613), .A2(new_n615), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n658), .A2(new_n664), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n518), .B(new_n317), .C1(new_n707), .C2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n842), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n842), .A2(new_n846), .A3(KEYINPUT113), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT114), .B1(new_n835), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n712), .A2(KEYINPUT104), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n712), .A2(KEYINPUT104), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n834), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n833), .ZN(new_n858));
  AND4_X1   g672(.A1(KEYINPUT114), .A2(new_n853), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n675), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n627), .A2(new_n719), .ZN(new_n862));
  INV_X1    g676(.A(new_n672), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n862), .A2(new_n189), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n688), .A3(new_n752), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n743), .A2(new_n861), .A3(new_n700), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT52), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n675), .B1(new_n735), .B2(new_n742), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n700), .A4(new_n865), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n826), .B1(new_n860), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n835), .A2(KEYINPUT114), .A3(new_n853), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n867), .A2(new_n870), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n743), .A2(new_n861), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n826), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n872), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT115), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n881), .A2(new_n835), .A3(KEYINPUT53), .A4(new_n853), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n871), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n872), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n891), .A3(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n825), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(G952), .A2(G953), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n780), .A2(new_n601), .A3(new_n606), .A4(new_n836), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT110), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n691), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n687), .A3(new_n901), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n894), .A2(new_n895), .B1(new_n896), .B2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n871), .A2(new_n888), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n879), .B2(new_n826), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n191), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(G210), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n509), .A2(new_n512), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n511), .ZN(new_n909));
  XNOR2_X1  g723(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n907), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n281), .A2(G952), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G51));
  NAND2_X1  g730(.A1(new_n872), .A2(new_n889), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(G902), .A3(new_n769), .A4(new_n768), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n315), .B(KEYINPUT57), .Z(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n872), .A2(new_n921), .A3(new_n887), .A4(new_n889), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT53), .B1(new_n877), .B2(new_n878), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT54), .B1(new_n923), .B2(new_n904), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n905), .B2(new_n887), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n308), .ZN(new_n928));
  INV_X1    g742(.A(new_n309), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n919), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT122), .B1(new_n931), .B2(new_n915), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n933));
  INV_X1    g747(.A(new_n915), .ZN(new_n934));
  INV_X1    g748(.A(new_n930), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n890), .A2(KEYINPUT121), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(new_n924), .A3(new_n922), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n920), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n933), .B(new_n934), .C1(new_n938), .C2(new_n919), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n932), .A2(new_n939), .ZN(G54));
  NAND3_X1  g754(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n941));
  INV_X1    g755(.A(new_n461), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n944), .A3(new_n915), .ZN(G60));
  AND2_X1   g759(.A1(new_n630), .A2(new_n631), .ZN(new_n946));
  XNOR2_X1  g760(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n318), .A2(new_n191), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n893), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n937), .A2(new_n946), .A3(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n915), .A3(new_n951), .ZN(G63));
  XNOR2_X1  g766(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT60), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n917), .A2(KEYINPUT124), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n905), .B2(new_n956), .ZN(new_n960));
  INV_X1    g774(.A(new_n593), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n934), .ZN(new_n963));
  INV_X1    g777(.A(new_n661), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n958), .B2(new_n960), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n954), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n965), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n967), .A2(new_n934), .A3(new_n962), .A4(new_n953), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(G66));
  AOI21_X1  g783(.A(new_n281), .B1(new_n438), .B2(G224), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n853), .A2(new_n857), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n281), .ZN(new_n972));
  INV_X1    g786(.A(G898), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n908), .B1(new_n973), .B2(G953), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G69));
  AND2_X1   g789(.A1(new_n792), .A2(new_n788), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n862), .A2(new_n602), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n777), .A2(new_n778), .A3(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n868), .A2(new_n700), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n762), .A2(new_n978), .A3(new_n764), .A4(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n980), .A3(new_n281), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n544), .B1(new_n535), .B2(KEYINPUT30), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(new_n447), .Z(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(G900), .B2(G953), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n979), .A2(new_n694), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT62), .Z(new_n988));
  NOR2_X1   g802(.A1(new_n843), .A2(new_n628), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n757), .B1(new_n989), .B2(new_n796), .ZN(new_n990));
  OR4_X1    g804(.A1(new_n602), .A2(new_n990), .A3(new_n677), .A4(new_n679), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n976), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n983), .B1(new_n992), .B2(new_n281), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n986), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n994), .B(new_n995), .Z(G72));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT127), .ZN(new_n998));
  XNOR2_X1  g812(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n976), .A2(new_n980), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n971), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n546), .A2(new_n540), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n915), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n546), .A2(new_n541), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n558), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n884), .A2(new_n1000), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1000), .B1(new_n992), .B2(new_n971), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n684), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1004), .A2(new_n1007), .A3(new_n1009), .ZN(G57));
endmodule


