//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  NAND2_X1  g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT92), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n209), .B2(KEYINPUT91), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT91), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(new_n206), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n204), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n209), .A2(new_n205), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n219), .A2(new_n216), .A3(new_n204), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT17), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G1gat), .B2(new_n224), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G8gat), .ZN(new_n228));
  INV_X1    g027(.A(G8gat), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n226), .B(new_n229), .C1(G1gat), .C2(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n234), .B(KEYINPUT93), .Z(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n222), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT94), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT94), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n231), .A2(new_n239), .A3(new_n222), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n233), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT97), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n246));
  XNOR2_X1  g045(.A(G169gat), .B(G197gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n231), .A2(new_n222), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n253), .A2(KEYINPUT95), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(KEYINPUT95), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n241), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n235), .B(KEYINPUT13), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n223), .A2(new_n232), .B1(new_n238), .B2(new_n240), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(KEYINPUT18), .A3(new_n236), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n245), .A2(new_n252), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT18), .B1(new_n259), .B2(new_n236), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(new_n243), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT98), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n262), .A2(new_n243), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n251), .B1(new_n262), .B2(new_n243), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n258), .A2(new_n260), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT98), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n258), .A2(new_n260), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n251), .B1(new_n270), .B2(new_n262), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT96), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT96), .B(new_n251), .C1(new_n270), .C2(new_n262), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n264), .A2(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT99), .ZN(new_n277));
  INV_X1    g076(.A(G57gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(G64gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(G64gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G71gat), .B(G78gat), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n282), .ZN(new_n284));
  OR3_X1    g083(.A1(new_n278), .A2(KEYINPUT100), .A3(G64gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT100), .B1(new_n278), .B2(G64gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n277), .B(new_n284), .C1(new_n279), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n232), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(G183gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G231gat), .A2(G233gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G155gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT20), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n294), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n290), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(G211gat), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n298), .B(new_n300), .Z(new_n301));
  OR2_X1    g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n297), .A2(new_n301), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT103), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT102), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(G85gat), .A3(G92gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT7), .ZN(new_n308));
  INV_X1    g107(.A(G85gat), .ZN(new_n309));
  INV_X1    g108(.A(G92gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G99gat), .ZN(new_n312));
  INV_X1    g111(.A(G106gat), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT8), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G99gat), .B(G106gat), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n315), .A2(new_n317), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n305), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n320), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(KEYINPUT103), .A3(new_n318), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n223), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT104), .ZN(new_n325));
  AND2_X1   g124(.A1(G232gat), .A2(G233gat), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n324), .A2(new_n325), .B1(KEYINPUT41), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n321), .A2(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n222), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n327), .B(new_n329), .C1(new_n325), .C2(new_n324), .ZN(new_n330));
  XNOR2_X1  g129(.A(G190gat), .B(G218gat), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n326), .A2(KEYINPUT41), .ZN(new_n333));
  XNOR2_X1  g132(.A(G134gat), .B(G162gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n331), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n332), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G230gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT106), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n316), .A2(KEYINPUT105), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n315), .B(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n283), .A2(new_n288), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n322), .A2(new_n289), .A3(new_n318), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT106), .B1(new_n344), .B2(new_n345), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n348), .A2(KEYINPUT10), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n328), .A2(KEYINPUT10), .A3(new_n345), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n341), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n341), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n348), .B2(new_n349), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G120gat), .B(G148gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(G176gat), .B(G204gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n353), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n304), .A2(new_n340), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT70), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n367));
  AND2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  INV_X1    g167(.A(G169gat), .ZN(new_n369));
  INV_X1    g168(.A(G176gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OR2_X1    g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT64), .B1(new_n380), .B2(KEYINPUT23), .ZN(new_n381));
  AND4_X1   g180(.A1(KEYINPUT64), .A2(new_n369), .A3(new_n370), .A4(KEYINPUT23), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n373), .B(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT65), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n387));
  OAI221_X1 g186(.A(new_n377), .B1(new_n387), .B2(new_n375), .C1(new_n376), .C2(KEYINPUT66), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n380), .A2(KEYINPUT23), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(KEYINPUT25), .A3(new_n373), .A4(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n383), .A2(new_n391), .A3(new_n384), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT27), .B(G183gat), .ZN(new_n394));
  INV_X1    g193(.A(G190gat), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT67), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT28), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n371), .A2(KEYINPUT26), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n371), .A2(KEYINPUT26), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n400), .B(new_n401), .C1(new_n369), .C2(new_n370), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n397), .A2(KEYINPUT28), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n399), .A2(new_n374), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n393), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G127gat), .B(G134gat), .Z(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT1), .ZN(new_n408));
  INV_X1    g207(.A(G120gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(G113gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT68), .B(G120gat), .ZN(new_n411));
  INV_X1    g210(.A(G113gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n408), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n412), .A2(G120gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n407), .B1(new_n416), .B2(KEYINPUT1), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n367), .B1(new_n406), .B2(new_n419), .ZN(new_n420));
  AOI211_X1 g219(.A(KEYINPUT69), .B(new_n418), .C1(new_n393), .C2(new_n405), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n393), .A2(new_n418), .A3(new_n405), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n366), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n419), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT69), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n406), .A2(new_n367), .A3(new_n419), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n425), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(KEYINPUT70), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G15gat), .B(G43gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n424), .A2(new_n366), .A3(new_n425), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT70), .B1(new_n430), .B2(new_n431), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT32), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT34), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n443), .A3(new_n425), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n428), .A2(new_n422), .A3(new_n425), .A4(new_n429), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT34), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n433), .B2(KEYINPUT32), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n439), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G78gat), .B(G106gat), .ZN(new_n452));
  INV_X1    g251(.A(G22gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(KEYINPUT31), .B(G50gat), .Z(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT3), .ZN(new_n458));
  INV_X1    g257(.A(G148gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(G141gat), .ZN(new_n460));
  INV_X1    g259(.A(G141gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G148gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT73), .B(KEYINPUT2), .ZN(new_n464));
  INV_X1    g263(.A(G162gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G155gat), .ZN(new_n466));
  INV_X1    g265(.A(G155gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G162gat), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n463), .A2(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n467), .A2(G162gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n465), .A2(G155gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT75), .ZN(new_n475));
  OR2_X1    g274(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n476));
  OR2_X1    g275(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n474), .A2(new_n475), .B1(new_n480), .B2(KEYINPUT2), .ZN(new_n481));
  OR3_X1    g280(.A1(new_n459), .A2(KEYINPUT74), .A3(G141gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n462), .A2(KEYINPUT74), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n460), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT78), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n474), .A2(new_n475), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n476), .A2(new_n478), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT77), .B(G162gat), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT2), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND4_X1   g288(.A1(KEYINPUT78), .A2(new_n486), .A3(new_n484), .A4(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n458), .B(new_n470), .C1(new_n485), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT79), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n486), .A2(new_n489), .A3(new_n484), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT78), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT78), .A4(new_n484), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n469), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT79), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n458), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT29), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G211gat), .ZN(new_n501));
  INV_X1    g300(.A(G218gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT22), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(G211gat), .B2(G218gat), .ZN(new_n506));
  XOR2_X1   g305(.A(G197gat), .B(G204gat), .Z(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G211gat), .A2(G218gat), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(new_n503), .C1(new_n507), .C2(new_n504), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n500), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G228gat), .A2(G233gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n515), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n508), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT29), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(KEYINPUT85), .A3(new_n519), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n458), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n470), .B1(new_n485), .B2(new_n490), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(KEYINPUT86), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n514), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n519), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n497), .B1(new_n458), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n513), .B1(new_n512), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n457), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n527), .A2(new_n528), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n535), .B(new_n456), .C1(new_n536), .C2(new_n514), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n442), .A2(new_n448), .ZN(new_n539));
  INV_X1    g338(.A(new_n438), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n540), .B1(new_n433), .B2(new_n434), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n433), .A2(KEYINPUT32), .A3(new_n447), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n451), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n511), .ZN(new_n545));
  INV_X1    g344(.A(G226gat), .ZN(new_n546));
  INV_X1    g345(.A(G233gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n406), .B2(new_n519), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n546), .B(new_n547), .C1(new_n393), .C2(new_n405), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n406), .A2(new_n548), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT29), .B1(new_n393), .B2(new_n405), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n552), .B(new_n511), .C1(new_n548), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G8gat), .B(G36gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n310), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT72), .B(G64gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n551), .A2(new_n554), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(KEYINPUT30), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n551), .A2(new_n564), .A3(new_n554), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n418), .B(new_n470), .C1(new_n485), .C2(new_n490), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(KEYINPUT80), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT80), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n570), .B1(new_n497), .B2(new_n418), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT4), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n418), .B1(new_n525), .B2(KEYINPUT3), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n491), .A2(KEYINPUT79), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n498), .B1(new_n497), .B2(new_n458), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT4), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n568), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n572), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n580));
  NAND2_X1  g379(.A1(G225gat), .A2(G233gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT80), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n497), .A2(new_n570), .A3(new_n418), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n577), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n497), .A2(KEYINPUT4), .A3(new_n418), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n576), .A2(new_n581), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT82), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n525), .A2(new_n419), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n581), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n580), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n589), .B1(new_n588), .B2(new_n593), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n583), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G1gat), .B(G29gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G85gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT0), .B(G57gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n600), .B(new_n583), .C1(new_n594), .C2(new_n595), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n596), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n567), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n544), .A2(KEYINPUT35), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT35), .B1(new_n544), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n591), .A2(new_n592), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT87), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT87), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n579), .B2(new_n592), .ZN(new_n615));
  OAI211_X1 g414(.A(KEYINPUT39), .B(new_n613), .C1(new_n615), .C2(new_n612), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n579), .A2(new_n592), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n601), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n616), .A2(new_n619), .A3(KEYINPUT40), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n622), .A2(new_n602), .A3(new_n567), .A4(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n562), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT37), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n551), .B2(new_n554), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n551), .A2(new_n626), .A3(new_n554), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT88), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n551), .A2(KEYINPUT88), .A3(new_n626), .A4(new_n554), .ZN(new_n631));
  AOI211_X1 g430(.A(new_n561), .B(new_n627), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n625), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n605), .A2(new_n607), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT89), .B1(new_n632), .B2(new_n633), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT89), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n630), .A2(new_n631), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n559), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n637), .B(KEYINPUT38), .C1(new_n639), .C2(new_n627), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n538), .B(new_n624), .C1(new_n635), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n605), .A2(new_n607), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n566), .ZN(new_n644));
  INV_X1    g443(.A(new_n538), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n451), .A2(new_n543), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT71), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT36), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n539), .A2(new_n542), .A3(new_n541), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n541), .B1(new_n539), .B2(new_n542), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT36), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n642), .A2(new_n646), .A3(new_n649), .A4(new_n654), .ZN(new_n655));
  AOI211_X1 g454(.A(new_n275), .B(new_n365), .C1(new_n611), .C2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n643), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g458(.A1(new_n656), .A2(new_n567), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT16), .B(G8gat), .Z(new_n661));
  OAI211_X1 g460(.A(new_n660), .B(new_n661), .C1(KEYINPUT107), .C2(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n664), .B(new_n665), .C1(new_n229), .C2(new_n660), .ZN(G1325gat));
  INV_X1    g465(.A(new_n647), .ZN(new_n667));
  AOI21_X1  g466(.A(G15gat), .B1(new_n656), .B2(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT108), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT108), .ZN(new_n670));
  INV_X1    g469(.A(new_n654), .ZN(new_n671));
  INV_X1    g470(.A(new_n649), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n669), .A2(new_n670), .B1(new_n656), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n645), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n453), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  AND4_X1   g479(.A1(new_n646), .A2(new_n642), .A3(new_n649), .A4(new_n654), .ZN(new_n681));
  INV_X1    g480(.A(new_n610), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n544), .A2(KEYINPUT35), .A3(new_n608), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n339), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n340), .B1(new_n611), .B2(new_n655), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n304), .A2(new_n363), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n273), .A2(new_n274), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n264), .A2(new_n269), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n692), .B2(new_n693), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n690), .A2(new_n657), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n690), .A2(KEYINPUT111), .A3(new_n657), .A4(new_n698), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(G29gat), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n611), .A2(new_n655), .ZN(new_n704));
  INV_X1    g503(.A(new_n275), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n339), .A4(new_n691), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n207), .A3(new_n657), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n703), .A2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n208), .A3(new_n567), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(KEYINPUT46), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(KEYINPUT112), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT46), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n690), .A2(new_n567), .A3(new_n698), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n715), .B(new_n716), .C1(new_n208), .C2(new_n717), .ZN(G1329gat));
  NOR3_X1   g517(.A1(new_n706), .A2(G43gat), .A3(new_n647), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n687), .A2(new_n674), .A3(new_n689), .A4(new_n698), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(G43gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n538), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n687), .A2(new_n689), .A3(new_n698), .A4(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n706), .B2(new_n538), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n725), .A2(KEYINPUT114), .A3(new_n727), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(KEYINPUT48), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n731), .B1(new_n732), .B2(new_n734), .ZN(G1331gat));
  NAND2_X1  g534(.A1(new_n304), .A2(new_n340), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n611), .B2(new_n655), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n697), .A2(new_n364), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n643), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n278), .ZN(G1332gat));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n566), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n739), .B2(new_n673), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n739), .A2(G71gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n647), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g549(.A1(new_n739), .A2(new_n538), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(G78gat), .Z(G1335gat));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n697), .A2(new_n304), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n688), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n688), .B2(new_n754), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n757), .A2(new_n309), .A3(new_n657), .A4(new_n363), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n697), .A2(new_n304), .A3(new_n364), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n687), .A2(new_n657), .A3(new_n689), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G85gat), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n759), .B1(new_n758), .B2(new_n762), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(G1336gat));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n687), .A2(new_n567), .A3(new_n689), .A4(new_n760), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n768), .B2(KEYINPUT116), .ZN(new_n769));
  INV_X1    g568(.A(new_n756), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n688), .A2(new_n753), .A3(new_n754), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n770), .A2(new_n310), .A3(new_n363), .A4(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n772), .B2(new_n566), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  OAI221_X1 g573(.A(new_n768), .B1(KEYINPUT116), .B2(new_n766), .C1(new_n772), .C2(new_n566), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1337gat));
  NAND4_X1  g575(.A1(new_n757), .A2(new_n312), .A3(new_n363), .A4(new_n667), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n687), .A2(new_n674), .A3(new_n689), .A4(new_n760), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G99gat), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n778), .B1(new_n777), .B2(new_n780), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(G1338gat));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n687), .A2(new_n645), .A3(new_n689), .A4(new_n760), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G106gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(KEYINPUT118), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n313), .A3(new_n363), .A4(new_n771), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n788), .B2(new_n538), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  OAI221_X1 g589(.A(new_n786), .B1(KEYINPUT118), .B2(new_n784), .C1(new_n788), .C2(new_n538), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(new_n304), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n346), .A2(new_n347), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT106), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT10), .ZN(new_n796));
  INV_X1    g595(.A(new_n349), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n354), .B1(new_n798), .B2(new_n351), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n361), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n351), .A3(new_n354), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n353), .A2(new_n802), .A3(KEYINPUT54), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n801), .A2(new_n803), .A3(KEYINPUT55), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n806), .A2(new_n362), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n695), .B2(new_n696), .ZN(new_n809));
  INV_X1    g608(.A(new_n250), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n256), .A2(new_n257), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n259), .A2(new_n236), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n693), .A2(new_n363), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n339), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n693), .A2(new_n813), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n808), .A2(new_n339), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n793), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n365), .A2(new_n697), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n544), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n643), .A2(new_n567), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n412), .A3(new_n697), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT119), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(KEYINPUT119), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n275), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n826), .B1(new_n830), .B2(new_n412), .ZN(G1340gat));
  OR3_X1    g630(.A1(new_n827), .A2(new_n411), .A3(new_n364), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n364), .B1(new_n828), .B2(new_n829), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n409), .ZN(G1341gat));
  NAND3_X1  g633(.A1(new_n825), .A2(KEYINPUT120), .A3(new_n304), .ZN(new_n835));
  INV_X1    g634(.A(G127gat), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n827), .B2(new_n793), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n793), .B1(new_n828), .B2(new_n829), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(G127gat), .B2(new_n840), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n842), .A3(new_n339), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n340), .B1(new_n828), .B2(new_n829), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n842), .ZN(G1343gat));
  AOI21_X1  g646(.A(new_n538), .B1(new_n819), .B2(new_n821), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n673), .A2(new_n824), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n806), .A2(new_n362), .A3(new_n807), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n814), .B1(new_n852), .B2(new_n275), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n340), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n304), .B1(new_n854), .B2(new_n817), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n645), .B1(new_n855), .B2(new_n820), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n851), .B1(new_n856), .B2(KEYINPUT57), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n461), .B1(new_n859), .B2(new_n697), .ZN(new_n860));
  INV_X1    g659(.A(new_n851), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n848), .A2(new_n861), .A3(new_n461), .A4(new_n705), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT58), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n862), .B(KEYINPUT121), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n857), .A3(new_n705), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(G141gat), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n865), .A2(KEYINPUT123), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT123), .B1(new_n865), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n864), .B1(new_n869), .B2(new_n870), .ZN(G1344gat));
  AOI211_X1 g670(.A(KEYINPUT59), .B(new_n459), .C1(new_n859), .C2(new_n363), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n365), .A2(new_n705), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n849), .B(new_n645), .C1(new_n855), .C2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n848), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n363), .A3(new_n861), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n873), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n848), .A2(new_n861), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n363), .A2(new_n459), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n872), .A2(new_n880), .B1(new_n881), .B2(new_n882), .ZN(G1345gat));
  NOR3_X1   g682(.A1(new_n858), .A2(new_n487), .A3(new_n793), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n848), .A2(new_n304), .A3(new_n861), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n487), .B2(new_n885), .ZN(G1346gat));
  NOR3_X1   g685(.A1(new_n858), .A2(new_n488), .A3(new_n340), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n848), .A2(new_n339), .A3(new_n861), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n488), .B2(new_n888), .ZN(G1347gat));
  NAND2_X1  g688(.A1(new_n643), .A2(new_n567), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n823), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n275), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n697), .A2(new_n369), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(G1348gat));
  NOR2_X1   g694(.A1(new_n892), .A2(new_n364), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(new_n370), .ZN(G1349gat));
  INV_X1    g696(.A(new_n892), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n304), .A3(new_n394), .ZN(new_n899));
  OAI21_X1  g698(.A(G183gat), .B1(new_n892), .B2(new_n793), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(KEYINPUT124), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT60), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n899), .A2(KEYINPUT124), .A3(new_n900), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n898), .A2(new_n395), .A3(new_n339), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(KEYINPUT125), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(KEYINPUT125), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n898), .A2(new_n339), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(G190gat), .ZN(new_n911));
  AOI211_X1 g710(.A(KEYINPUT61), .B(new_n395), .C1(new_n898), .C2(new_n339), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n907), .A2(new_n908), .B1(new_n911), .B2(new_n912), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n674), .A2(new_n890), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n914), .B(new_n875), .C1(new_n848), .C2(new_n849), .ZN(new_n915));
  OAI21_X1  g714(.A(G197gat), .B1(new_n915), .B2(new_n275), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n848), .A2(new_n914), .ZN(new_n917));
  INV_X1    g716(.A(G197gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n697), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1352gat));
  XNOR2_X1  g719(.A(KEYINPUT126), .B(G204gat), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n363), .A3(new_n922), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n878), .A2(new_n363), .A3(new_n914), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n924), .B(new_n925), .C1(new_n922), .C2(new_n926), .ZN(G1353gat));
  OAI21_X1  g726(.A(G211gat), .B1(new_n915), .B2(new_n793), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT63), .Z(new_n929));
  NAND3_X1  g728(.A1(new_n917), .A2(new_n501), .A3(new_n304), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1354gat));
  OAI21_X1  g730(.A(G218gat), .B1(new_n915), .B2(new_n340), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n502), .A3(new_n339), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1355gat));
endmodule


