//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(G250), .B1(G257), .B2(G264), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(new_n213), .B2(new_n214), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n209), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n222), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n215), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n207), .A2(G1), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(KEYINPUT67), .A3(G50), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(new_n255), .B2(new_n201), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n254), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G50), .B2(new_n250), .ZN(new_n261));
  INV_X1    g0061(.A(new_n253), .ZN(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT8), .B(G58), .Z(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(new_n265), .B1(G150), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1698), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G222), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G223), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(G1698), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n274), .B1(new_n224), .B2(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  AND2_X1   g0081(.A1(G1), .A2(G13), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT65), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT65), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n206), .C1(G41), .C2(G45), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n284), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n282), .A2(new_n283), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n291), .A2(new_n285), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT66), .B(G226), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n280), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n270), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G179), .B2(new_n295), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n270), .B(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n295), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G190), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n301), .A2(new_n303), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT10), .B1(new_n310), .B2(new_n307), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n299), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n254), .A2(G68), .A3(new_n256), .ZN(new_n313));
  XOR2_X1   g0113(.A(new_n313), .B(KEYINPUT70), .Z(new_n314));
  AOI22_X1  g0114(.A1(new_n265), .A2(G77), .B1(G20), .B2(new_n217), .ZN(new_n315));
  INV_X1    g0115(.A(new_n266), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n201), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n317), .A2(new_n253), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n318), .A2(KEYINPUT11), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n251), .A2(new_n217), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT12), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(KEYINPUT11), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n314), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G97), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT69), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G33), .A3(G97), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n273), .B2(G226), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  OAI211_X1 g0131(.A(G232), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n291), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n291), .A2(G238), .A3(new_n285), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n289), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT13), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n289), .A2(new_n334), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n325), .A2(new_n327), .ZN(new_n338));
  INV_X1    g0138(.A(G1698), .ZN(new_n339));
  OAI211_X1 g0139(.A(G226), .B(new_n339), .C1(new_n330), .C2(new_n331), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n279), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT13), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n323), .B1(new_n346), .B2(G190), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n306), .B2(new_n346), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n337), .A2(new_n342), .A3(new_n343), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n337), .B2(new_n342), .ZN(new_n350));
  OAI21_X1  g0150(.A(G169), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n336), .A2(G179), .A3(new_n344), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT14), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(G169), .C1(new_n349), .C2(new_n350), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n323), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n254), .A2(G77), .A3(new_n256), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G77), .B2(new_n250), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(new_n263), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n316), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n360), .B1(new_n365), .B2(new_n253), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n330), .A2(new_n331), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n273), .A2(G232), .B1(new_n367), .B2(G107), .ZN(new_n368));
  INV_X1    g0168(.A(G238), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n277), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n279), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n290), .B1(G244), .B2(new_n292), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n366), .B1(new_n373), .B2(new_n296), .ZN(new_n374));
  INV_X1    g0174(.A(G179), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n373), .A2(G200), .ZN(new_n378));
  INV_X1    g0178(.A(G190), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n378), .B(new_n366), .C1(new_n379), .C2(new_n373), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n380), .A3(KEYINPUT68), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n377), .A2(new_n380), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(KEYINPUT68), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n312), .A2(new_n358), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n364), .A2(new_n255), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n254), .B1(new_n251), .B2(new_n364), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n367), .B2(new_n207), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NOR4_X1   g0189(.A1(new_n330), .A2(new_n331), .A3(new_n389), .A4(G20), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G159), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n392), .A2(G20), .A3(G33), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(G58), .A3(G68), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n397), .A3(new_n218), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(G20), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n262), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(new_n393), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT72), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT72), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n406), .B(new_n393), .C1(new_n398), .C2(G20), .ZN(new_n407));
  OAI211_X1 g0207(.A(KEYINPUT16), .B(new_n391), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n387), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n276), .A2(new_n339), .ZN(new_n411));
  INV_X1    g0211(.A(G226), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n411), .B(new_n413), .C1(new_n330), .C2(new_n331), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n279), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n291), .A2(G232), .A3(new_n285), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n417), .A2(G179), .A3(new_n289), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n289), .A2(new_n418), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n291), .B1(new_n414), .B2(new_n415), .ZN(new_n421));
  OAI21_X1  g0221(.A(G169), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n409), .A2(new_n410), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n389), .B1(new_n275), .B2(G20), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n367), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n217), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n399), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n401), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n408), .A2(new_n253), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n423), .B1(new_n430), .B2(new_n386), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT73), .B1(new_n431), .B2(KEYINPUT18), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT73), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n410), .C1(new_n409), .C2(new_n423), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n424), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n417), .A2(G190), .A3(new_n289), .A4(new_n418), .ZN(new_n436));
  OAI21_X1  g0236(.A(G200), .B1(new_n420), .B2(new_n421), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n430), .A2(new_n386), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n384), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n250), .A2(G107), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT25), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n206), .A2(G33), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n250), .A2(new_n448), .A3(new_n215), .A4(new_n252), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G107), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G116), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G20), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT23), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n207), .B2(G107), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n207), .B(G87), .C1(new_n330), .C2(new_n331), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(KEYINPUT22), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT24), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n452), .B1(new_n466), .B2(new_n253), .ZN(new_n467));
  OAI211_X1 g0267(.A(G257), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT77), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT77), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n275), .A2(new_n470), .A3(G257), .A4(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G294), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n275), .A2(G250), .A3(new_n339), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n279), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n480), .A2(G264), .A3(new_n291), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT78), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT78), .ZN(new_n484));
  AOI211_X1 g0284(.A(new_n484), .B(new_n481), .C1(new_n474), .C2(new_n279), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n284), .A2(new_n477), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(G200), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n475), .A2(new_n482), .ZN(new_n490));
  INV_X1    g0290(.A(new_n488), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n490), .A2(G190), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n467), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n484), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n481), .B1(new_n474), .B2(new_n279), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT78), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n494), .A2(G179), .A3(new_n488), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n296), .B1(new_n495), .B2(new_n488), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n467), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT74), .ZN(new_n504));
  AND2_X1   g0304(.A1(KEYINPUT4), .A2(G244), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n339), .B(new_n505), .C1(new_n330), .C2(new_n331), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n225), .B1(new_n271), .B2(new_n272), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(KEYINPUT4), .ZN(new_n509));
  OAI21_X1  g0309(.A(G250), .B1(new_n330), .B2(new_n331), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n339), .B1(new_n510), .B2(KEYINPUT4), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n279), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n279), .B1(new_n477), .B2(new_n487), .ZN(new_n513));
  INV_X1    g0313(.A(new_n480), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n513), .A2(G257), .B1(new_n514), .B2(new_n284), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n504), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n504), .A3(new_n515), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(G190), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT6), .ZN(new_n520));
  INV_X1    g0320(.A(G97), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n520), .A2(new_n521), .A3(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n524), .A2(new_n207), .B1(new_n224), .B2(new_n316), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n226), .B1(new_n425), .B2(new_n426), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n253), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n250), .A2(G97), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n450), .B2(G97), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n306), .B1(new_n512), .B2(new_n515), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n512), .A2(new_n504), .A3(new_n515), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n296), .B1(new_n533), .B2(new_n516), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n512), .A2(new_n515), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n375), .B1(new_n527), .B2(new_n529), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n519), .A2(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G87), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n521), .A3(new_n226), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n325), .B2(new_n327), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(G20), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n207), .B(G68), .C1(new_n330), .C2(new_n331), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n540), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n262), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n362), .A2(new_n250), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n449), .A2(new_n538), .ZN(new_n549));
  OR3_X1    g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n369), .A2(new_n339), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n225), .A2(G1698), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(new_n330), .C2(new_n331), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n291), .B1(new_n553), .B2(new_n453), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n477), .A2(new_n281), .ZN(new_n555));
  INV_X1    g0355(.A(G250), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n476), .B2(G1), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n291), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G190), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n306), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n550), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n548), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n449), .A2(new_n361), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n542), .A2(new_n546), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n564), .B(new_n566), .C1(new_n567), .C2(new_n262), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n547), .A2(new_n548), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT76), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n566), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n553), .A2(new_n453), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n375), .B(new_n558), .C1(new_n574), .C2(new_n291), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT75), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n560), .A2(KEYINPUT75), .A3(new_n375), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n558), .B1(new_n574), .B2(new_n291), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n577), .A2(new_n578), .B1(new_n296), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n563), .B1(new_n573), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n513), .A2(G270), .B1(new_n514), .B2(new_n284), .ZN(new_n582));
  OAI211_X1 g0382(.A(G257), .B(new_n339), .C1(new_n330), .C2(new_n331), .ZN(new_n583));
  OAI211_X1 g0383(.A(G264), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n584));
  INV_X1    g0384(.A(G303), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n275), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n279), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n450), .A2(G116), .ZN(new_n589));
  INV_X1    g0389(.A(G116), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n251), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n252), .A2(new_n215), .B1(G20), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n507), .B(new_n207), .C1(G33), .C2(new_n521), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT20), .B1(new_n592), .B2(new_n593), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n589), .B(new_n591), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n588), .A2(new_n596), .A3(KEYINPUT21), .A4(G169), .ZN(new_n597));
  INV_X1    g0397(.A(new_n596), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n582), .A2(new_n587), .A3(G190), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n582), .A2(new_n587), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n306), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n588), .A2(new_n596), .A3(G169), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n600), .A2(G179), .A3(new_n596), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n597), .A2(new_n601), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n537), .A2(new_n581), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n503), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n445), .A2(new_n608), .ZN(G372));
  NAND3_X1  g0409(.A1(new_n604), .A2(new_n605), .A3(new_n597), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n502), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n519), .A2(new_n532), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n534), .A2(new_n536), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n554), .A2(KEYINPUT79), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT79), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n616), .B(new_n291), .C1(new_n553), .C2(new_n453), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n558), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n296), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n568), .A3(new_n575), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(G200), .ZN(new_n621));
  INV_X1    g0421(.A(new_n549), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n621), .A2(new_n570), .A3(new_n622), .A4(new_n561), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n613), .A2(new_n614), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n612), .A2(new_n624), .A3(new_n493), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n534), .A2(new_n536), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n581), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT26), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n627), .A2(new_n630), .A3(new_n620), .A4(new_n623), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n620), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n445), .B1(new_n626), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n410), .B1(new_n409), .B2(new_n423), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n430), .A2(new_n386), .ZN(new_n635));
  INV_X1    g0435(.A(new_n423), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(KEYINPUT18), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n348), .A2(new_n376), .A3(new_n374), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(new_n357), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n640), .B2(new_n443), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT80), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n305), .B1(new_n304), .B2(new_n308), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n310), .A2(KEYINPUT10), .A3(new_n307), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n309), .A2(KEYINPUT80), .A3(new_n311), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n299), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n633), .A2(new_n648), .ZN(G369));
  NAND3_X1  g0449(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT81), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT82), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n655), .A2(G213), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g0457(.A(KEYINPUT83), .B(G343), .Z(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n501), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n493), .A2(new_n502), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT84), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT84), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n493), .A2(new_n663), .A3(new_n502), .A4(new_n660), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n659), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n502), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n659), .A2(new_n596), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n606), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n611), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n611), .A2(new_n659), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n662), .A2(new_n664), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n467), .B1(new_n497), .B2(new_n499), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n666), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n673), .A2(new_n678), .ZN(G399));
  NOR2_X1   g0479(.A1(new_n211), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n539), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n219), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n537), .A2(new_n581), .A3(new_n606), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n502), .A3(new_n493), .A4(new_n666), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n588), .A2(new_n579), .A3(new_n375), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n494), .A2(new_n689), .A3(new_n496), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n517), .A2(new_n518), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n533), .A2(new_n516), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n486), .A2(new_n693), .A3(KEYINPUT30), .A4(new_n689), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n618), .A2(new_n375), .A3(new_n588), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n535), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n494), .A2(new_n488), .A3(new_n496), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n692), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n659), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n687), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT85), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n483), .A2(new_n485), .A3(new_n491), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n498), .B1(new_n708), .B2(G179), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n707), .B(new_n611), .C1(new_n709), .C2(new_n467), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT85), .B1(new_n676), .B2(new_n610), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(new_n493), .A4(new_n624), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n571), .B1(new_n570), .B2(new_n566), .ZN(new_n713));
  NOR4_X1   g0513(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n548), .A4(new_n565), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n580), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n563), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n627), .A2(new_n630), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n623), .A2(new_n620), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT26), .B1(new_n718), .B2(new_n614), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n717), .A2(new_n719), .A3(new_n620), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n666), .B1(new_n626), .B2(new_n632), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n706), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n685), .B1(new_n726), .B2(G1), .ZN(G364));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n215), .B1(G20), .B2(new_n296), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n211), .A2(new_n275), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G45), .B2(new_n219), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(G45), .B2(new_n245), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n210), .A2(new_n275), .ZN(new_n736));
  INV_X1    g0536(.A(G355), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n736), .A2(new_n737), .B1(G116), .B2(new_n210), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n732), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n207), .A2(G13), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n206), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n680), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n207), .A2(G179), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n379), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n275), .B1(new_n747), .B2(G283), .ZN(new_n748));
  INV_X1    g0548(.A(G294), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n379), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n207), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n379), .A3(new_n306), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT92), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G329), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n748), .B1(new_n749), .B2(new_n751), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n745), .A2(G190), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT91), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(G20), .A2(G179), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT86), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n763), .A2(G303), .B1(G326), .B2(new_n767), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n765), .A2(new_n379), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(KEYINPUT33), .B(G317), .Z(new_n771));
  OAI21_X1  g0571(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT87), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n765), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n765), .A2(new_n773), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n775), .A2(G190), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n757), .B(new_n772), .C1(G322), .C2(new_n778), .ZN(new_n779));
  AND3_X1   g0579(.A1(new_n775), .A2(new_n379), .A3(new_n776), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT88), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT88), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n777), .A2(new_n202), .B1(new_n201), .B2(new_n766), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n783), .B2(G77), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT89), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n763), .A2(G87), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT90), .B(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n752), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n751), .A2(new_n521), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n746), .A2(new_n226), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n794), .A2(new_n795), .A3(new_n367), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n769), .A2(G68), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n790), .A2(new_n793), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n786), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n744), .B1(new_n799), .B2(new_n731), .ZN(new_n800));
  INV_X1    g0600(.A(new_n730), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n671), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n672), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n743), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(G330), .B2(new_n671), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  NAND3_X1  g0607(.A1(new_n666), .A2(new_n376), .A3(new_n374), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n380), .B1(new_n666), .B2(new_n366), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n377), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n723), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n666), .B(new_n811), .C1(new_n626), .C2(new_n632), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n706), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  INV_X1    g0616(.A(new_n743), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n813), .A2(new_n814), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n816), .B(new_n817), .C1(new_n706), .C2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n731), .A2(new_n728), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n743), .B1(G77), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT93), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n784), .A2(new_n590), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n367), .B1(new_n762), .B2(new_n226), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT94), .Z(new_n826));
  NOR2_X1   g0626(.A1(new_n777), .A2(new_n749), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n746), .A2(new_n538), .ZN(new_n828));
  INV_X1    g0628(.A(new_n755), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n794), .B(new_n828), .C1(new_n829), .C2(G311), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n831), .B2(new_n770), .C1(new_n585), .C2(new_n766), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n824), .A2(new_n826), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G137), .A2(new_n767), .B1(new_n769), .B2(G150), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT95), .B(G143), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n777), .B2(new_n835), .C1(new_n784), .C2(new_n791), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n275), .B1(new_n746), .B2(new_n217), .ZN(new_n839));
  INV_X1    g0639(.A(new_n751), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(G58), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n762), .B2(new_n201), .C1(new_n842), .C2(new_n755), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n836), .B2(new_n837), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n833), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n731), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n823), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(KEYINPUT96), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(KEYINPUT96), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(new_n729), .C2(new_n811), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n819), .A2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(new_n524), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n852), .A2(KEYINPUT35), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(KEYINPUT35), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n853), .A2(G116), .A3(new_n216), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT36), .Z(new_n856));
  NAND4_X1  g0656(.A1(new_n220), .A2(G77), .A3(new_n397), .A4(new_n395), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n857), .A2(KEYINPUT98), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n857), .A2(KEYINPUT98), .B1(new_n201), .B2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n206), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT101), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n408), .A2(new_n253), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n391), .B1(new_n405), .B2(new_n407), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n401), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n387), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n657), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n435), .B2(new_n443), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n439), .B1(new_n866), .B2(new_n657), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n866), .A2(new_n423), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n430), .A2(new_n386), .A3(new_n438), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n409), .A2(new_n657), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n431), .A2(KEYINPUT100), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT100), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n409), .A2(new_n877), .A3(new_n423), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n873), .B(new_n875), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n868), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n868), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n862), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n868), .A2(new_n880), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n868), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(KEYINPUT101), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n355), .A2(new_n353), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n354), .B1(new_n345), .B2(G169), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n323), .B(new_n659), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT99), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n356), .A2(KEYINPUT99), .A3(new_n323), .A4(new_n659), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n659), .A2(new_n323), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n348), .A2(new_n357), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n811), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n486), .A2(new_n693), .A3(new_n689), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n901), .A2(new_n688), .B1(new_n697), .B2(new_n696), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n666), .B1(new_n902), .B2(new_n694), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n608), .A2(new_n666), .B1(KEYINPUT31), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n700), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n699), .A2(KEYINPUT104), .A3(new_n659), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n701), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n900), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT40), .B1(new_n889), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT17), .B1(new_n409), .B2(new_n438), .ZN(new_n912));
  AND4_X1   g0712(.A1(KEYINPUT17), .A2(new_n430), .A3(new_n386), .A4(new_n438), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n875), .B1(new_n914), .B2(new_n638), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n439), .B(new_n916), .C1(new_n409), .C2(new_n657), .ZN(new_n917));
  INV_X1    g0717(.A(new_n431), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n877), .ZN(new_n919));
  INV_X1    g0719(.A(new_n878), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n872), .A2(new_n431), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n916), .B1(new_n922), .B2(new_n875), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n915), .A2(KEYINPUT103), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n925), .B(new_n875), .C1(new_n914), .C2(new_n638), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n885), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n911), .B1(new_n927), .B2(new_n887), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n910), .B1(new_n909), .B2(new_n928), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n444), .B(new_n384), .C1(new_n904), .C2(new_n908), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(G330), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n929), .A2(new_n930), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n634), .A2(new_n637), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n874), .B1(new_n937), .B2(new_n443), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n918), .A2(new_n439), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT37), .B1(new_n939), .B2(new_n874), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n938), .A2(new_n925), .B1(new_n879), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n926), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n936), .B1(new_n943), .B2(new_n881), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n356), .A2(new_n323), .A3(new_n666), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT102), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n896), .A2(new_n898), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n814), .B2(new_n808), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n881), .A2(new_n882), .A3(new_n862), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT101), .B1(new_n886), .B2(new_n887), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n937), .A2(new_n657), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n725), .A2(new_n445), .A3(new_n722), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n648), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n935), .A2(new_n959), .B1(new_n206), .B2(new_n740), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n935), .A2(new_n959), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n861), .B1(new_n960), .B2(new_n961), .ZN(G367));
  NAND2_X1  g0762(.A1(new_n659), .A2(new_n550), .ZN(new_n963));
  MUX2_X1   g0763(.A(new_n620), .B(new_n718), .S(new_n963), .Z(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT105), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n659), .A2(new_n530), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n537), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n627), .A2(new_n659), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n662), .A2(new_n664), .A3(new_n674), .A4(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT42), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n614), .B1(new_n968), .B2(new_n502), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n971), .A2(KEYINPUT42), .B1(new_n666), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT106), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n972), .B2(new_n974), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n966), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n972), .A2(new_n974), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT106), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n981), .B(new_n976), .C1(KEYINPUT43), .C2(new_n965), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n673), .A2(new_n970), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n983), .B1(new_n979), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n680), .B(KEYINPUT41), .Z(new_n987));
  NAND3_X1  g0787(.A1(new_n675), .A2(new_n677), .A3(new_n970), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n675), .A2(KEYINPUT45), .A3(new_n677), .A4(new_n970), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n970), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT44), .B1(new_n678), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n995), .B(new_n970), .C1(new_n675), .C2(new_n677), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n990), .A2(new_n992), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n673), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n678), .A2(new_n993), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n995), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n678), .A2(KEYINPUT44), .A3(new_n993), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n673), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n988), .A2(new_n989), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n991), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n665), .A2(new_n667), .A3(new_n674), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n672), .A3(new_n675), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n675), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n803), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n998), .A2(new_n1006), .A3(new_n726), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n987), .B1(new_n1013), .B2(new_n726), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n986), .B1(new_n1014), .B2(new_n742), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n770), .A2(new_n791), .B1(new_n766), .B2(new_n835), .ZN(new_n1016));
  INV_X1    g0816(.A(G137), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n275), .B1(new_n752), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G68), .B2(new_n840), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n224), .B2(new_n746), .C1(new_n202), .C2(new_n762), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1016), .B(new_n1020), .C1(G150), .C2(new_n778), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n784), .B2(new_n201), .ZN(new_n1022));
  AOI21_X1  g0822(.A(KEYINPUT46), .B1(new_n763), .B2(G116), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(KEYINPUT107), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1023), .A2(KEYINPUT107), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G303), .C2(new_n778), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1027));
  INV_X1    g0827(.A(G317), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n367), .B1(new_n752), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G107), .B2(new_n840), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n521), .B2(new_n746), .C1(new_n770), .C2(new_n749), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G311), .B2(new_n767), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1026), .A2(new_n1027), .A3(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n784), .A2(new_n831), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1022), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n731), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n732), .B1(new_n210), .B2(new_n361), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n733), .B2(new_n241), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n817), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(new_n801), .C2(new_n965), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1015), .A2(new_n1041), .ZN(G387));
  AOI22_X1  g0842(.A1(new_n763), .A2(G294), .B1(G283), .B2(new_n840), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G322), .A2(new_n767), .B1(new_n769), .B2(G311), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n777), .B2(new_n1028), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n783), .B2(G303), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n1046), .B2(KEYINPUT48), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT48), .B2(new_n1046), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT49), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n752), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n275), .B1(new_n1050), .B2(G326), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n590), .B2(new_n746), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n778), .A2(G50), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n767), .A2(G159), .ZN(new_n1055));
  INV_X1    g0855(.A(G150), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n275), .B1(new_n752), .B2(new_n1056), .C1(new_n521), .C2(new_n746), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n362), .B2(new_n840), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n763), .A2(G77), .B1(new_n263), .B2(new_n769), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n783), .B2(G68), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n731), .B1(new_n1053), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n238), .A2(new_n476), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n263), .A2(new_n201), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n682), .B(new_n476), .C1(new_n217), .C2(new_n224), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n733), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1063), .B1(KEYINPUT108), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(KEYINPUT108), .B2(new_n1067), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(G107), .B2(new_n210), .C1(new_n682), .C2(new_n736), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n817), .B1(new_n1070), .B2(new_n732), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1062), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n668), .B2(new_n730), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n742), .B2(new_n1012), .ZN(new_n1074));
  OR3_X1    g0874(.A1(new_n1012), .A2(KEYINPUT109), .A3(new_n726), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1012), .A2(new_n726), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT109), .B1(new_n1012), .B2(new_n726), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1075), .A2(new_n680), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1074), .A2(new_n1078), .ZN(G393));
  NOR2_X1   g0879(.A1(new_n997), .A2(new_n673), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1076), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n680), .A3(new_n1013), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n998), .A2(new_n742), .A3(new_n1006), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT111), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n275), .B1(new_n752), .B2(new_n835), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n828), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n840), .A2(G77), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n201), .B2(new_n770), .C1(new_n217), .C2(new_n762), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n777), .A2(new_n392), .B1(new_n1056), .B2(new_n766), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT51), .Z(new_n1092));
  AOI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(new_n263), .C2(new_n783), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(KEYINPUT110), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n777), .A2(new_n785), .B1(new_n1028), .B2(new_n766), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  INV_X1    g0897(.A(G322), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n367), .B1(new_n752), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n795), .B(new_n1099), .C1(G116), .C2(new_n840), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n585), .B2(new_n770), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G283), .B2(new_n763), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1097), .B(new_n1102), .C1(new_n784), .C2(new_n749), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT110), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1103), .B1(new_n1093), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n731), .B1(new_n1095), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n733), .A2(new_n248), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n730), .B(new_n731), .C1(new_n211), .C2(G97), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n817), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(new_n801), .C2(new_n970), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1084), .A2(new_n1085), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1085), .B1(new_n1084), .B2(new_n1110), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1083), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT112), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(KEYINPUT112), .B(new_n1083), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(G390));
  NAND3_X1  g0917(.A1(new_n704), .A2(G330), .A3(new_n811), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1118), .A2(new_n950), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT39), .B1(new_n927), .B2(new_n887), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n881), .A2(new_n882), .A3(new_n936), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1120), .A2(new_n1121), .B1(new_n951), .B2(new_n947), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n810), .A2(new_n377), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n659), .B(new_n1123), .C1(new_n712), .C2(new_n720), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n899), .B1(new_n1124), .B2(new_n809), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n947), .B1(new_n927), .B2(new_n887), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT113), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1119), .B(new_n1122), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n946), .B1(new_n943), .B2(new_n881), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n810), .A2(new_n377), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n721), .A2(new_n666), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n950), .B1(new_n1133), .B2(new_n808), .ZN(new_n1134));
  OAI21_X1  g0934(.A(KEYINPUT113), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n951), .A2(new_n947), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n944), .A2(new_n948), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1135), .A2(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n900), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n906), .A2(new_n701), .A3(new_n907), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n687), .A2(new_n703), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(G330), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1130), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n814), .A2(new_n808), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1118), .A2(KEYINPUT114), .A3(new_n950), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1143), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT114), .B1(new_n1118), .B2(new_n950), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(G330), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n950), .B1(new_n1150), .B2(new_n812), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1151), .A2(new_n1119), .A3(new_n808), .A4(new_n1133), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n445), .B(G330), .C1(new_n1142), .C2(new_n1141), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n957), .A3(new_n648), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1144), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1122), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1143), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1155), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n1162), .A3(new_n1130), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n680), .A3(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1130), .B(new_n742), .C1(new_n1139), .C2(new_n1143), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT115), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT115), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1161), .A2(new_n1167), .A3(new_n742), .A4(new_n1130), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT54), .B(G143), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n784), .A2(new_n1170), .B1(new_n1017), .B2(new_n770), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1171), .A2(KEYINPUT116), .B1(G159), .B2(new_n840), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(KEYINPUT116), .B2(new_n1171), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT117), .Z(new_n1174));
  NOR2_X1   g0974(.A1(new_n762), .A2(new_n1056), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT53), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n275), .B1(new_n746), .B2(new_n201), .ZN(new_n1177));
  INV_X1    g0977(.A(G128), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n766), .A2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(new_n829), .C2(G125), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1176), .B(new_n1180), .C1(new_n842), .C2(new_n777), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT118), .B1(new_n1174), .B2(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n755), .A2(new_n749), .B1(new_n217), .B2(new_n746), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT119), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n790), .A2(new_n367), .A3(new_n1088), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n770), .A2(new_n226), .B1(new_n831), .B2(new_n766), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n590), .B2(new_n777), .C1(new_n784), .C2(new_n521), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1174), .A2(KEYINPUT118), .A3(new_n1181), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n731), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1138), .A2(new_n728), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n817), .B1(new_n364), .B2(new_n820), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1164), .A2(new_n1169), .A3(new_n1194), .ZN(G378));
  NAND3_X1  g0995(.A1(new_n645), .A2(new_n298), .A3(new_n646), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n657), .A2(new_n270), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1197), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n645), .A2(new_n298), .A3(new_n646), .A4(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n927), .A2(new_n887), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n909), .A3(KEYINPUT40), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(G330), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1204), .B1(new_n910), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1201), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n933), .B1(new_n928), .B2(new_n909), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n883), .B2(new_n888), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1213), .B(new_n1214), .C1(new_n1216), .C2(KEYINPUT40), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1208), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n956), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1208), .A2(new_n956), .A3(new_n1217), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1204), .A2(new_n728), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n743), .B1(G50), .B2(new_n821), .ZN(new_n1224));
  INV_X1    g1024(.A(G41), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n367), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n840), .B2(G68), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n202), .B2(new_n746), .C1(new_n755), .C2(new_n831), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n770), .A2(new_n521), .B1(new_n762), .B2(new_n224), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G116), .C2(new_n767), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n226), .B2(new_n777), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n362), .B2(new_n783), .ZN(new_n1232));
  XOR2_X1   g1032(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1233));
  AOI21_X1  g1033(.A(G50), .B1(new_n264), .B2(new_n1225), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1232), .A2(new_n1233), .B1(new_n1226), .B2(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G33), .B(G41), .C1(new_n1050), .C2(G124), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n791), .B2(new_n746), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT121), .Z(new_n1238));
  NOR2_X1   g1038(.A1(new_n777), .A2(new_n1178), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1170), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n763), .A2(new_n1240), .B1(G125), .B2(new_n767), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n842), .B2(new_n770), .C1(new_n1056), .C2(new_n751), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1239), .B(new_n1242), .C1(new_n783), .C2(G137), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT59), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1238), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1243), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1235), .B1(new_n1233), .B2(new_n1232), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1224), .B1(new_n1248), .B2(new_n731), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1222), .A2(new_n742), .B1(new_n1223), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1130), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1143), .B1(new_n1252), .B2(new_n1122), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1155), .B1(new_n1254), .B2(new_n1153), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1208), .A2(new_n956), .A3(new_n1217), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n956), .B1(new_n1208), .B2(new_n1217), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT57), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n680), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1163), .A2(new_n1156), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT57), .B1(new_n1260), .B2(new_n1222), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1250), .B1(new_n1259), .B2(new_n1261), .ZN(G375));
  OAI21_X1  g1062(.A(new_n743), .B1(G68), .B2(new_n821), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n899), .A2(new_n729), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n275), .B1(new_n747), .B2(G77), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n361), .B2(new_n751), .C1(new_n755), .C2(new_n585), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n763), .A2(G97), .B1(G116), .B2(new_n769), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n749), .B2(new_n766), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1266), .B(new_n1268), .C1(G283), .C2(new_n778), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n784), .B2(new_n226), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n275), .B1(new_n746), .B2(new_n202), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G50), .B2(new_n840), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1272), .B1(new_n762), .B2(new_n392), .C1(new_n1178), .C2(new_n755), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n783), .B2(G150), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT122), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(G132), .A2(new_n767), .B1(new_n769), .B2(new_n1240), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n777), .B2(new_n1017), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1270), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1263), .B(new_n1264), .C1(new_n731), .C2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1153), .B2(new_n742), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n987), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1157), .A2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1280), .B1(new_n1282), .B2(new_n1283), .ZN(G381));
  NAND3_X1  g1084(.A1(new_n1074), .A2(new_n806), .A3(new_n1078), .ZN(new_n1285));
  OR3_X1    g1085(.A1(new_n1285), .A2(G381), .A3(G384), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1286), .A2(G390), .A3(G387), .ZN(new_n1287));
  XOR2_X1   g1087(.A(new_n1287), .B(KEYINPUT123), .Z(new_n1288));
  NOR2_X1   g1088(.A1(G375), .A2(G378), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G407));
  NAND2_X1  g1090(.A1(new_n658), .A2(G213), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT124), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(G407), .A2(G213), .A3(new_n1293), .ZN(G409));
  NAND3_X1  g1094(.A1(new_n1260), .A2(new_n1222), .A3(new_n1281), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1250), .A2(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1164), .A2(new_n1169), .A3(new_n1194), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1292), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G375), .A2(G378), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1149), .A2(new_n1152), .A3(KEYINPUT60), .A4(new_n1155), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(new_n1157), .A3(new_n680), .A4(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1303), .A2(G384), .A3(new_n1280), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G384), .B1(new_n1303), .B2(new_n1280), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1298), .A2(new_n1299), .B1(KEYINPUT125), .B2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G2897), .B(new_n1292), .C1(new_n1306), .C2(KEYINPUT125), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1292), .A2(G2897), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1309), .B(new_n1310), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G393), .A2(G396), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1285), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G387), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1041), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1013), .A2(new_n726), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1281), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n741), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1319), .B1(new_n1322), .B2(new_n986), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1084), .A2(new_n1110), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT111), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1084), .A2(new_n1085), .A3(new_n1110), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT112), .B1(new_n1327), .B2(new_n1083), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1116), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1323), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(G387), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1318), .A2(new_n1332), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1330), .A2(new_n1317), .A3(new_n1331), .A4(new_n1315), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1336), .B1(new_n1337), .B2(new_n1306), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1306), .ZN(new_n1340));
  NOR3_X1   g1140(.A1(new_n1339), .A2(KEYINPUT63), .A3(new_n1340), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1313), .B(new_n1335), .C1(new_n1338), .C2(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(KEYINPUT62), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1337), .A2(new_n1344), .A3(new_n1306), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1313), .A2(new_n1343), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1342), .B1(new_n1346), .B2(new_n1335), .ZN(G405));
  NAND3_X1  g1147(.A1(new_n1260), .A2(new_n1222), .A3(KEYINPUT57), .ZN(new_n1348));
  AOI22_X1  g1148(.A1(new_n1156), .A2(new_n1163), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1348), .B(new_n680), .C1(KEYINPUT57), .C2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1350), .A2(new_n1297), .A3(new_n1250), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1299), .A2(KEYINPUT127), .A3(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(KEYINPUT127), .B1(new_n1299), .B2(new_n1351), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1334), .B(new_n1333), .C1(new_n1352), .C2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1299), .A2(KEYINPUT127), .A3(new_n1351), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT127), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1297), .B1(new_n1350), .B2(new_n1250), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1356), .B1(new_n1289), .B2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1330), .A2(KEYINPUT126), .ZN(new_n1359));
  AOI22_X1  g1159(.A1(new_n1359), .A2(new_n1315), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1334), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1355), .B(new_n1358), .C1(new_n1360), .C2(new_n1361), .ZN(new_n1362));
  AND3_X1   g1162(.A1(new_n1354), .A2(new_n1362), .A3(new_n1306), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1306), .B1(new_n1354), .B2(new_n1362), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1363), .A2(new_n1364), .ZN(G402));
endmodule


