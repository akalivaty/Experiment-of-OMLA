//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G107), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR4_X1   g0023(.A1(new_n214), .A2(new_n217), .A3(new_n220), .A4(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT65), .B(G77), .Z(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G244), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n208), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  INV_X1    g0029(.A(G250), .ZN(new_n230));
  INV_X1    g0030(.A(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n208), .A2(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n230), .B(new_n232), .C1(new_n211), .C2(new_n213), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n202), .A2(G50), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n235), .A2(new_n207), .A3(new_n236), .ZN(new_n237));
  NOR3_X1   g0037(.A1(new_n229), .A2(new_n234), .A3(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n216), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  INV_X1    g0043(.A(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT66), .B(G264), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT67), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G68), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G50), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n252), .B(new_n255), .Z(G351));
  AOI21_X1  g0056(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT77), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(KEYINPUT3), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(new_n260), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT76), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(KEYINPUT76), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n259), .B(G33), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n222), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G244), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n269), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G116), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n260), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n258), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n206), .A2(G45), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n258), .A2(G250), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT84), .ZN(new_n283));
  INV_X1    g0083(.A(new_n279), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G274), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n282), .A2(new_n283), .A3(G190), .A4(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n263), .A2(new_n268), .B1(new_n272), .B2(G1698), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n276), .B1(new_n287), .B2(new_n271), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n285), .B(new_n280), .C1(new_n288), .C2(new_n258), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT84), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(G200), .ZN(new_n293));
  XOR2_X1   g0093(.A(KEYINPUT15), .B(G87), .Z(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n206), .A2(G20), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n231), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT82), .ZN(new_n299));
  AOI211_X1 g0099(.A(G20), .B(new_n221), .C1(new_n263), .C2(new_n268), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G97), .A2(G107), .ZN(new_n301));
  INV_X1    g0101(.A(G87), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT19), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n304), .A2(new_n260), .A3(new_n210), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n305), .B2(G20), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n260), .A2(G20), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G97), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n304), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n299), .B1(new_n300), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n236), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n269), .A2(new_n207), .A3(G68), .ZN(new_n314));
  INV_X1    g0114(.A(new_n310), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(KEYINPUT82), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n311), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  AOI211_X1 g0117(.A(new_n313), .B(new_n297), .C1(new_n206), .C2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G87), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n293), .A2(new_n298), .A3(new_n317), .A4(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n292), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n289), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n294), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n317), .A2(new_n324), .A3(new_n298), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT83), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT83), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n317), .A2(new_n327), .A3(new_n324), .A4(new_n298), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n323), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n321), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n333));
  INV_X1    g0133(.A(G274), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n258), .A2(new_n333), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n266), .A2(G33), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n226), .A2(new_n341), .ZN(new_n342));
  MUX2_X1   g0142(.A(G222), .B(G223), .S(G1698), .Z(new_n343));
  OAI21_X1  g0143(.A(new_n257), .B1(new_n343), .B2(new_n340), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n336), .B1(new_n337), .B2(new_n219), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  XOR2_X1   g0145(.A(new_n345), .B(KEYINPUT68), .Z(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G190), .ZN(new_n347));
  INV_X1    g0147(.A(G200), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n346), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT8), .B(G58), .Z(new_n350));
  NAND3_X1  g0150(.A1(new_n207), .A2(new_n260), .A3(KEYINPUT69), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT69), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(G20), .B2(G33), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n307), .A2(new_n350), .B1(new_n354), .B2(G150), .ZN(new_n355));
  XOR2_X1   g0155(.A(new_n355), .B(KEYINPUT70), .Z(new_n356));
  AOI21_X1  g0156(.A(new_n207), .B1(new_n201), .B2(new_n218), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT71), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n313), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n297), .A2(new_n218), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT72), .ZN(new_n361));
  INV_X1    g0161(.A(new_n296), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(new_n218), .ZN(new_n363));
  INV_X1    g0163(.A(new_n297), .ZN(new_n364));
  INV_X1    g0164(.A(new_n313), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n296), .A2(KEYINPUT72), .A3(G50), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n363), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n359), .A2(new_n360), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT9), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n349), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n372), .B(new_n373), .C1(new_n371), .C2(new_n370), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT10), .B1(new_n370), .B2(new_n349), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n375), .A2(new_n376), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n346), .A2(new_n330), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n368), .C1(G169), .C2(new_n346), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n202), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n354), .A2(G159), .B1(new_n384), .B2(G20), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n263), .A2(new_n207), .A3(new_n268), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n221), .B1(new_n387), .B2(KEYINPUT7), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n263), .A2(new_n389), .A3(new_n268), .A4(new_n207), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n386), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n340), .B2(new_n207), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n266), .A2(KEYINPUT76), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT78), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .A4(new_n260), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n395), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT78), .B(new_n339), .C1(new_n399), .C2(G33), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n393), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n385), .B1(new_n401), .B2(new_n221), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n392), .A2(new_n404), .A3(new_n313), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n350), .A2(new_n297), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n362), .A2(new_n313), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n408), .B2(new_n350), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(G223), .A2(G1698), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n270), .A2(G226), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n269), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT79), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n260), .C2(new_n302), .ZN(new_n418));
  AOI211_X1 g0218(.A(new_n412), .B(new_n414), .C1(new_n263), .C2(new_n268), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n260), .A2(new_n302), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT79), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n421), .A3(new_n257), .ZN(new_n422));
  INV_X1    g0222(.A(new_n337), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n335), .B1(new_n423), .B2(G232), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(G179), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G169), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n422), .B2(new_n424), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n411), .B(KEYINPUT18), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n422), .A2(new_n424), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G169), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT18), .B1(new_n433), .B2(new_n411), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(G200), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n365), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n409), .B1(new_n437), .B2(new_n404), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n422), .A2(G190), .A3(new_n424), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT17), .A4(new_n439), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n435), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n216), .A2(G1698), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(G226), .B2(G1698), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n447), .A2(new_n340), .B1(new_n260), .B2(new_n210), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n335), .B1(new_n448), .B2(new_n257), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n222), .B2(new_n337), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT13), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G169), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(KEYINPUT14), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n451), .A2(new_n330), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT14), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n451), .B2(G169), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n297), .A2(new_n221), .ZN(new_n458));
  XOR2_X1   g0258(.A(new_n458), .B(KEYINPUT12), .Z(new_n459));
  INV_X1    g0259(.A(new_n354), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n218), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n307), .A2(G77), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n207), .B2(G68), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n313), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  XOR2_X1   g0264(.A(new_n464), .B(KEYINPUT11), .Z(new_n465));
  AOI211_X1 g0265(.A(new_n459), .B(new_n465), .C1(G68), .C2(new_n407), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n451), .A2(G200), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n466), .B(new_n468), .C1(new_n290), .C2(new_n451), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n225), .A2(new_n297), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT73), .ZN(new_n473));
  INV_X1    g0273(.A(G77), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n226), .A2(G20), .B1(new_n294), .B2(new_n307), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n350), .A2(new_n354), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI221_X1 g0277(.A(new_n473), .B1(new_n474), .B2(new_n408), .C1(new_n477), .C2(new_n365), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n222), .A2(G1698), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(G232), .B2(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n258), .B1(new_n341), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G107), .B2(new_n341), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(new_n336), .C1(new_n272), .C2(new_n337), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n427), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n478), .B(new_n484), .C1(G179), .C2(new_n483), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n445), .A2(new_n471), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n478), .B1(G200), .B2(new_n483), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n290), .B2(new_n483), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n382), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n364), .A2(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n354), .A2(G77), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n212), .A2(KEYINPUT6), .A3(G97), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n210), .A2(new_n212), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n301), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G20), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n492), .B(new_n497), .C1(new_n401), .C2(new_n212), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n491), .B1(new_n498), .B2(new_n313), .ZN(new_n499));
  INV_X1    g0299(.A(new_n318), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n210), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n270), .A2(G244), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n269), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT80), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT4), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n502), .A2(new_n506), .B1(new_n230), .B2(new_n270), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n341), .A2(new_n508), .B1(G33), .B2(G283), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n263), .B2(new_n268), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT80), .B1(new_n510), .B2(KEYINPUT4), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n257), .ZN(new_n513));
  XOR2_X1   g0313(.A(KEYINPUT5), .B(G41), .Z(new_n514));
  OAI21_X1  g0314(.A(new_n258), .B1(new_n514), .B2(new_n279), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n211), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n285), .A2(new_n514), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n513), .A2(new_n330), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n516), .B(new_n518), .C1(new_n512), .C2(new_n257), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n501), .B(new_n520), .C1(new_n521), .C2(G169), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n513), .A2(G190), .A3(new_n517), .A4(new_n519), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n500), .A2(new_n210), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n491), .B(new_n525), .C1(new_n498), .C2(new_n313), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n526), .C1(new_n521), .C2(new_n348), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT81), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n516), .B1(new_n512), .B2(new_n257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n519), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G200), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(KEYINPUT81), .A3(new_n526), .A4(new_n524), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n523), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n276), .A2(new_n207), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n207), .A2(G107), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n536), .B(KEYINPUT23), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT22), .A2(G87), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n338), .A2(KEYINPUT77), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n399), .B2(G33), .ZN(new_n541));
  AOI211_X1 g0341(.A(KEYINPUT77), .B(new_n260), .C1(new_n394), .C2(new_n395), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n207), .B(new_n539), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT86), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n341), .A2(new_n207), .A3(G87), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT22), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n543), .B2(new_n547), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n535), .B(new_n537), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT24), .ZN(new_n551));
  AOI211_X1 g0351(.A(G20), .B(new_n538), .C1(new_n263), .C2(new_n268), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n545), .A2(new_n546), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT86), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(new_n535), .A4(new_n537), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n313), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT25), .B1(new_n297), .B2(new_n212), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n212), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n318), .A2(G107), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n230), .A2(new_n270), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n211), .A2(G1698), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n269), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G294), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n258), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n515), .A2(new_n213), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n569), .A2(new_n518), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G190), .ZN(new_n572));
  INV_X1    g0372(.A(new_n570), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n567), .A2(new_n568), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n519), .B(new_n573), .C1(new_n574), .C2(new_n258), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G200), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n560), .A2(new_n564), .A3(new_n572), .A4(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT87), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n571), .B2(new_n427), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(KEYINPUT87), .A3(G169), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n571), .A2(G179), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n365), .B1(new_n551), .B2(new_n558), .ZN(new_n583));
  INV_X1    g0383(.A(new_n564), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G283), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n586), .B(new_n207), .C1(G33), .C2(new_n210), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n275), .A2(G20), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n313), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(KEYINPUT85), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n318), .A2(G116), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n589), .A2(new_n595), .A3(new_n590), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n297), .A2(new_n275), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n211), .A2(new_n270), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n213), .A2(G1698), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n269), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n340), .A2(G303), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n258), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n519), .B1(new_n515), .B2(new_n244), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n598), .B(G169), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n603), .A2(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G190), .ZN(new_n609));
  INV_X1    g0409(.A(new_n598), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n609), .B(new_n610), .C1(new_n348), .C2(new_n608), .ZN(new_n611));
  INV_X1    g0411(.A(new_n608), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(KEYINPUT21), .A3(G169), .A4(new_n598), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n608), .A2(G179), .A3(new_n598), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n607), .A2(new_n611), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n577), .A2(new_n585), .A3(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n332), .A2(new_n490), .A3(new_n534), .A4(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n529), .A2(new_n533), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n332), .A2(new_n618), .A3(new_n522), .A4(new_n577), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n613), .A2(new_n607), .A3(new_n614), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n585), .A2(KEYINPUT88), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT88), .B1(new_n585), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n326), .A2(new_n328), .ZN(new_n626));
  INV_X1    g0426(.A(new_n323), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n331), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n292), .A2(new_n320), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n523), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n332), .A2(KEYINPUT26), .A3(new_n523), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT89), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n329), .A2(KEYINPUT89), .A3(new_n331), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n632), .A2(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n490), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n467), .ZN(new_n640));
  AOI211_X1 g0440(.A(new_n444), .B(new_n470), .C1(new_n640), .C2(new_n485), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n379), .B1(new_n641), .B2(new_n435), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n381), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n644), .ZN(G369));
  NAND2_X1  g0445(.A1(new_n560), .A2(new_n564), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n207), .A2(G13), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .A3(G1), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT27), .B1(new_n647), .B2(G1), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g0450(.A(KEYINPUT90), .B(G343), .Z(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n585), .A3(new_n577), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n646), .A2(new_n582), .A3(new_n653), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n655), .B(new_n656), .C1(new_n621), .C2(new_n653), .ZN(new_n657));
  INV_X1    g0457(.A(new_n653), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n610), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n620), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n621), .A2(new_n611), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n659), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n621), .A2(new_n653), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n585), .A3(new_n577), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n646), .A2(new_n582), .A3(new_n658), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(G399));
  NOR2_X1   g0469(.A1(new_n303), .A2(G116), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT91), .Z(new_n671));
  NOR2_X1   g0471(.A1(new_n232), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n235), .B2(new_n673), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT93), .ZN(new_n676));
  XNOR2_X1  g0476(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT95), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n530), .A2(new_n571), .ZN(new_n681));
  NAND2_X1  g0481(.A1(KEYINPUT94), .A2(KEYINPUT30), .ZN(new_n682));
  NOR2_X1   g0482(.A1(KEYINPUT94), .A2(KEYINPUT30), .ZN(new_n683));
  NOR4_X1   g0483(.A1(new_n603), .A2(new_n330), .A3(new_n604), .A4(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n681), .A2(new_n322), .A3(new_n682), .A4(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n530), .A2(new_n684), .A3(new_n322), .A4(new_n571), .ZN(new_n686));
  INV_X1    g0486(.A(new_n682), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n571), .B1(new_n530), .B2(new_n519), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n330), .A3(new_n289), .A4(new_n612), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n680), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n686), .A2(new_n687), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n686), .A2(new_n687), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n680), .B(new_n691), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n653), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n618), .A2(new_n332), .A3(new_n522), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n577), .A2(new_n585), .A3(new_n615), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n698), .A2(new_n699), .A3(new_n653), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n689), .A2(new_n691), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n679), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT96), .ZN(new_n706));
  AND4_X1   g0506(.A1(KEYINPUT89), .A2(new_n626), .A3(new_n627), .A4(new_n331), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT89), .B1(new_n329), .B2(new_n331), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n635), .A2(KEYINPUT96), .A3(new_n636), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n632), .A2(new_n633), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n585), .A2(new_n621), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n534), .A2(new_n332), .A3(new_n577), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT97), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n715), .A2(new_n716), .A3(new_n658), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n715), .B2(new_n658), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT29), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n653), .B1(new_n625), .B2(new_n637), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n705), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n678), .B1(new_n723), .B2(G1), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT98), .ZN(G364));
  XNOR2_X1  g0525(.A(new_n647), .B(KEYINPUT99), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G45), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n727), .A2(KEYINPUT100), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(KEYINPUT100), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n672), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n663), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G330), .B2(new_n662), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n236), .B1(G20), .B2(new_n427), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n330), .A2(new_n348), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n207), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n341), .B1(new_n738), .B2(new_n221), .ZN(new_n739));
  NAND2_X1  g0539(.A1(G20), .A2(G190), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n330), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n741), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G50), .A2(new_n743), .B1(new_n746), .B2(G58), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n348), .A2(G179), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n741), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n302), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n737), .A2(new_n748), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n739), .B(new_n750), .C1(G107), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n330), .A2(new_n348), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT103), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n737), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G159), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT104), .B(KEYINPUT32), .Z(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n207), .B1(new_n756), .B2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G97), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n737), .A2(new_n744), .A3(KEYINPUT102), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT102), .B1(new_n737), .B2(new_n744), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n759), .A2(new_n760), .B1(new_n226), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n753), .A2(new_n761), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G294), .ZN(new_n771));
  INV_X1    g0571(.A(G303), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n762), .A2(new_n771), .B1(new_n772), .B2(new_n749), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(G329), .B2(new_n758), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n752), .A2(G283), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n768), .A2(G311), .ZN(new_n776));
  INV_X1    g0576(.A(new_n738), .ZN(new_n777));
  INV_X1    g0577(.A(G317), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(KEYINPUT105), .B(G326), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n743), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n341), .B(new_n784), .C1(G322), .C2(new_n746), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n735), .B1(new_n770), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n734), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n255), .A2(G45), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT101), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n269), .A2(new_n232), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(G45), .C2(new_n235), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n232), .A2(new_n340), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G355), .A2(new_n797), .B1(new_n275), .B2(new_n232), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n792), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n731), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n787), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n790), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n662), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n733), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n485), .A2(new_n653), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n478), .A2(new_n653), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n488), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(new_n808), .B2(new_n485), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n720), .B(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(new_n705), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n800), .ZN(new_n812));
  INV_X1    g0612(.A(new_n269), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G150), .A2(new_n777), .B1(new_n746), .B2(G143), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n815), .B2(new_n742), .C1(new_n767), .C2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT34), .Z(new_n818));
  AOI211_X1 g0618(.A(new_n813), .B(new_n818), .C1(G132), .C2(new_n758), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n819), .B1(new_n218), .B2(new_n749), .C1(new_n221), .C2(new_n751), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n762), .A2(new_n215), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n764), .B1(new_n822), .B2(new_n738), .C1(new_n823), .C2(new_n757), .ZN(new_n824));
  INV_X1    g0624(.A(new_n749), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(G107), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n752), .A2(G87), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(new_n275), .C2(new_n767), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n340), .B1(new_n745), .B2(new_n771), .C1(new_n772), .C2(new_n742), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n820), .A2(new_n821), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n734), .ZN(new_n831));
  INV_X1    g0631(.A(new_n809), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n800), .B1(new_n832), .B2(new_n788), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n734), .A2(new_n788), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n831), .B(new_n833), .C1(G77), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n812), .A2(new_n836), .ZN(G384));
  NOR2_X1   g0637(.A1(new_n726), .A2(new_n206), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT39), .ZN(new_n839));
  INV_X1    g0639(.A(new_n650), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n411), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n445), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n433), .A2(new_n411), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n843), .A2(new_n440), .A3(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT37), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n846), .A3(new_n440), .A4(new_n841), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT38), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n437), .B1(KEYINPUT16), .B2(new_n391), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n410), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n840), .B(new_n851), .C1(new_n435), .C2(new_n444), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n433), .B2(new_n840), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(new_n440), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n847), .B1(new_n854), .B2(new_n846), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n852), .A2(new_n855), .A3(KEYINPUT38), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n839), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n852), .A2(new_n855), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n856), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n858), .B1(new_n839), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n640), .A2(new_n653), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n435), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n466), .A2(new_n658), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n471), .A2(new_n869), .B1(new_n467), .B2(new_n653), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n618), .A2(new_n332), .A3(new_n522), .A4(new_n577), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n871), .A2(new_n623), .A3(new_n622), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT26), .B1(new_n332), .B2(new_n523), .ZN(new_n873));
  AND4_X1   g0673(.A1(KEYINPUT26), .A2(new_n628), .A3(new_n629), .A4(new_n523), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n873), .A2(new_n874), .B1(new_n708), .B2(new_n707), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n658), .B(new_n809), .C1(new_n872), .C2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n806), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n862), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n866), .B1(new_n867), .B2(new_n840), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n719), .A2(new_n490), .A3(new_n722), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT106), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n719), .A2(KEYINPUT106), .A3(new_n722), .A4(new_n490), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n643), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n881), .B(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n870), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n616), .A2(new_n332), .A3(new_n534), .A4(new_n658), .ZN(new_n889));
  INV_X1    g0689(.A(new_n696), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n692), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n889), .A2(KEYINPUT31), .B1(new_n891), .B2(new_n653), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n697), .A2(new_n701), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n809), .B(new_n888), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT107), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n891), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n702), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n898), .A2(KEYINPUT107), .A3(new_n809), .A4(new_n888), .ZN(new_n899));
  INV_X1    g0699(.A(new_n849), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n856), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n896), .A2(new_n899), .A3(KEYINPUT40), .A4(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n898), .A2(new_n862), .A3(new_n809), .A4(new_n888), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n679), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n490), .A2(G330), .A3(new_n898), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n903), .A2(new_n904), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n902), .A2(new_n490), .A3(new_n898), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT108), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n838), .B1(new_n887), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT109), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n913), .B2(new_n887), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n275), .B1(new_n496), .B2(KEYINPUT35), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n236), .A2(new_n207), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n917), .B(new_n918), .C1(KEYINPUT35), .C2(new_n496), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n202), .A2(G50), .A3(new_n383), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n921), .A2(new_n225), .B1(G50), .B2(new_n221), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n231), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n916), .A2(new_n920), .A3(new_n923), .ZN(G367));
  INV_X1    g0724(.A(new_n534), .ZN(new_n925));
  OR3_X1    g0725(.A1(new_n925), .A2(new_n666), .A3(KEYINPUT42), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT42), .B1(new_n925), .B2(new_n666), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n501), .A2(new_n653), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n534), .A2(new_n646), .A3(new_n582), .A4(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n653), .B1(new_n930), .B2(new_n522), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n928), .A2(KEYINPUT110), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n317), .A2(new_n298), .A3(new_n319), .ZN(new_n933));
  OR4_X1    g0733(.A1(new_n933), .A2(new_n707), .A3(new_n708), .A4(new_n658), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n332), .B1(new_n933), .B2(new_n658), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT43), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT110), .B1(new_n928), .B2(new_n931), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n932), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n534), .A2(new_n929), .B1(new_n523), .B2(new_n653), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n932), .A2(new_n938), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n939), .B1(new_n664), .B2(new_n940), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n664), .ZN(new_n944));
  INV_X1    g0744(.A(new_n940), .ZN(new_n945));
  INV_X1    g0745(.A(new_n939), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(new_n932), .B2(new_n938), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n672), .B(KEYINPUT41), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n666), .A2(new_n668), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n945), .A2(new_n953), .A3(KEYINPUT45), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT45), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n940), .B2(new_n952), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g0758(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT112), .Z(new_n960));
  NAND4_X1  g0760(.A1(new_n940), .A2(new_n952), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n940), .A2(new_n952), .A3(new_n958), .ZN(new_n962));
  INV_X1    g0762(.A(new_n960), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n957), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT113), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n664), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT114), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n957), .A2(new_n961), .A3(new_n964), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n968), .A2(new_n969), .B1(new_n970), .B2(new_n664), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(new_n967), .A3(KEYINPUT114), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n657), .A2(new_n663), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n667), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n971), .A2(new_n723), .A3(new_n972), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n951), .B1(new_n976), .B2(new_n723), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n949), .B1(new_n977), .B2(new_n730), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n763), .A2(G68), .B1(new_n226), .B2(new_n752), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n815), .B2(new_n757), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n340), .B(new_n980), .C1(G150), .C2(new_n746), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n777), .A2(G159), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n768), .A2(G50), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G143), .A2(new_n743), .B1(new_n825), .B2(G58), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT46), .B1(new_n825), .B2(G116), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n813), .B1(new_n210), .B2(new_n751), .C1(new_n757), .C2(new_n778), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT115), .Z(new_n988));
  AOI22_X1  g0788(.A1(G311), .A2(new_n743), .B1(new_n746), .B2(G303), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n825), .A2(KEYINPUT46), .A3(G116), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n771), .B2(new_n738), .C1(new_n767), .C2(new_n822), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G107), .B2(new_n763), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n985), .B1(new_n986), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT47), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n734), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n934), .A2(new_n790), .A3(new_n935), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n294), .A2(new_n232), .ZN(new_n998));
  INV_X1    g0798(.A(new_n795), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n791), .B(new_n998), .C1(new_n247), .C2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n731), .A3(new_n997), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n978), .A2(new_n1001), .ZN(G387));
  NAND2_X1  g0802(.A1(new_n715), .A2(new_n658), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT97), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n715), .A2(new_n716), .A3(new_n658), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n721), .B1(new_n1006), .B2(KEYINPUT29), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n974), .B1(new_n1007), .B2(new_n705), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n723), .A2(new_n975), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n1009), .A3(new_n672), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n743), .A2(G322), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n823), .B2(new_n738), .C1(new_n778), .C2(new_n745), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n768), .B2(G303), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT48), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n822), .B2(new_n762), .C1(new_n771), .C2(new_n749), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT49), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n269), .B1(new_n758), .B2(new_n782), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n275), .C2(new_n751), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n763), .A2(new_n294), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n218), .B2(new_n745), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT116), .Z(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(new_n813), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n758), .A2(G150), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n768), .A2(G68), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n225), .A2(new_n749), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n742), .A2(new_n816), .B1(new_n751), .B2(new_n210), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n350), .C2(new_n777), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n735), .B1(new_n1018), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(G45), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n795), .B1(new_n242), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n797), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n671), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n671), .B(new_n1030), .C1(new_n221), .C2(new_n474), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n350), .A2(new_n218), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT50), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1033), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n232), .A2(new_n212), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n792), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1029), .A2(new_n800), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n655), .A2(new_n656), .A3(new_n790), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n975), .A2(new_n730), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1010), .A2(new_n1042), .ZN(G393));
  XNOR2_X1  g0843(.A(new_n965), .B(new_n944), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1009), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n976), .A2(new_n1045), .A3(new_n672), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n730), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n940), .A2(new_n790), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n791), .B1(new_n252), .B2(new_n999), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G97), .B2(new_n232), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n738), .A2(new_n772), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G317), .A2(new_n743), .B1(new_n746), .B2(G311), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n762), .B2(new_n275), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1052), .B(new_n1055), .C1(G322), .C2(new_n758), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1053), .A2(KEYINPUT52), .B1(new_n767), .B2(new_n771), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n341), .B(new_n1057), .C1(G283), .C2(new_n825), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(new_n212), .C2(new_n751), .ZN(new_n1059));
  INV_X1    g0859(.A(G150), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n742), .A2(new_n1060), .B1(new_n745), .B2(new_n816), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n763), .A2(G77), .B1(new_n758), .B2(G143), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n269), .B1(new_n218), .B2(new_n738), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n827), .B1(new_n221), .B2(new_n749), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n768), .B2(new_n350), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1059), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n800), .B(new_n1051), .C1(new_n1070), .C2(new_n734), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1049), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1048), .A2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1046), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  NAND2_X1  g0875(.A1(new_n863), .A2(new_n788), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n341), .B1(new_n751), .B2(new_n218), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n758), .B2(G125), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT120), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT54), .B(G143), .Z(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n767), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n825), .A2(G150), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT53), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(G159), .C2(new_n763), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n746), .A2(G132), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n777), .A2(G137), .B1(new_n743), .B2(G128), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1080), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n762), .A2(new_n474), .B1(new_n757), .B2(new_n771), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G97), .B2(new_n768), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n746), .A2(G116), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n752), .A2(G68), .B1(new_n825), .B2(G87), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n742), .A2(new_n822), .B1(new_n738), .B2(new_n212), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n341), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n735), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1077), .A2(new_n800), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n350), .B2(new_n835), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT118), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n878), .B2(new_n864), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n806), .B1(new_n720), .B2(new_n809), .ZN(new_n1102));
  OAI211_X1 g0902(.A(KEYINPUT118), .B(new_n865), .C1(new_n1102), .C2(new_n870), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1103), .A3(new_n863), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1004), .A2(new_n1005), .A3(new_n877), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n808), .A2(new_n485), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n888), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n864), .B1(new_n900), .B2(new_n856), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n704), .ZN(new_n1110));
  OAI211_X1 g0910(.A(G330), .B(new_n809), .C1(new_n892), .C2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1111), .A2(new_n870), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1104), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT119), .B1(new_n894), .B2(new_n679), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n832), .B1(new_n702), .B2(new_n897), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT119), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1115), .A2(new_n1116), .A3(G330), .A4(new_n888), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1099), .B1(new_n1120), .B2(new_n1047), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1111), .A2(new_n870), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1114), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1102), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1115), .A2(G330), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n870), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n870), .C2(new_n1111), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1130), .A2(new_n886), .A3(new_n908), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1104), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n1118), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n673), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1120), .A2(new_n1131), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1121), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT106), .B1(new_n1007), .B2(new_n490), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n885), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n644), .B(new_n908), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT122), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n886), .A2(KEYINPUT122), .A3(new_n908), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n1120), .C2(new_n1131), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n866), .B1(new_n867), .B2(new_n840), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n879), .A2(new_n880), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n368), .A2(new_n840), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n382), .B(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT121), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n906), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n902), .A2(new_n905), .A3(KEYINPUT121), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1155), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT121), .B1(new_n902), .B2(new_n905), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1151), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1158), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1160), .B1(new_n1164), .B2(new_n1161), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1157), .A2(new_n1155), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n881), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1140), .B1(new_n1148), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1147), .A2(KEYINPUT57), .A3(new_n1163), .A4(new_n1167), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n672), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1163), .A2(new_n1167), .A3(new_n730), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n800), .B1(new_n1160), .B2(new_n788), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n763), .A2(G150), .B1(G128), .B2(new_n746), .ZN(new_n1174));
  INV_X1    g0974(.A(G132), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1082), .A2(new_n749), .B1(new_n1175), .B2(new_n738), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G125), .B2(new_n743), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1174), .B(new_n1177), .C1(new_n815), .C2(new_n767), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT59), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n752), .C2(G159), .ZN(new_n1180));
  INV_X1    g0980(.A(G124), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n757), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G33), .A2(G41), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n218), .B1(new_n269), .B2(G41), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1179), .A2(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G116), .A2(new_n743), .B1(new_n746), .B2(G107), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n210), .B2(new_n738), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1025), .B(new_n1187), .C1(G283), .C2(new_n758), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G41), .B(new_n269), .C1(new_n763), .C2(G68), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n768), .A2(new_n294), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n752), .A2(G58), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT58), .Z(new_n1193));
  OAI21_X1  g0993(.A(new_n734), .B1(new_n1185), .B2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1173), .B(new_n1194), .C1(G50), .C2(new_n835), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1172), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1171), .A2(new_n1197), .ZN(G375));
  INV_X1    g0998(.A(G128), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1191), .B1(new_n757), .B2(new_n1199), .C1(new_n762), .C2(new_n218), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n813), .B(new_n1200), .C1(G137), .C2(new_n746), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n777), .A2(new_n1081), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n768), .A2(G150), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G132), .A2(new_n743), .B1(new_n825), .B2(G159), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1019), .B1(new_n210), .B2(new_n749), .C1(new_n772), .C2(new_n757), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n341), .B(new_n1206), .C1(G294), .C2(new_n743), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G116), .A2(new_n777), .B1(new_n752), .B2(G77), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n212), .C2(new_n767), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n745), .A2(new_n822), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1205), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n734), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n731), .B(new_n1212), .C1(new_n888), .C2(new_n789), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n221), .B2(new_n834), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1130), .B2(new_n730), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n643), .B(new_n907), .C1(new_n884), .C2(new_n885), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n950), .B1(new_n1216), .B2(new_n1130), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1217), .B2(new_n1132), .ZN(G381));
  NOR2_X1   g1018(.A1(G375), .A2(G378), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n978), .A2(new_n1074), .A3(new_n1001), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1010), .A2(new_n804), .A3(new_n1042), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G381), .A2(G384), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT123), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1224), .B(new_n1225), .ZN(G407));
  NAND2_X1  g1026(.A1(new_n1219), .A2(new_n652), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(G407), .A2(G213), .A3(new_n1227), .ZN(G409));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1147), .A2(new_n950), .A3(new_n1163), .A4(new_n1167), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1138), .A2(new_n1230), .A3(new_n1172), .A4(new_n1195), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n652), .A2(G213), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G375), .B2(G378), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT60), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1216), .B2(new_n1130), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1112), .B1(new_n1106), .B2(new_n1105), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1127), .A2(new_n1237), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1143), .A2(KEYINPUT60), .A3(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n672), .A3(new_n1239), .A4(new_n1131), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1240), .A2(G384), .A3(new_n1215), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G384), .B1(new_n1240), .B2(new_n1215), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n652), .A2(G213), .A3(G2897), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1239), .A2(new_n672), .A3(new_n1131), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT60), .B1(new_n1143), .B2(new_n1238), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1215), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G384), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1240), .A2(G384), .A3(new_n1215), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1243), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1245), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1229), .B1(new_n1234), .B2(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1245), .A2(new_n1252), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1138), .B1(new_n1171), .B2(new_n1197), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(KEYINPUT125), .C1(new_n1256), .C2(new_n1233), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1256), .A2(new_n1260), .A3(new_n1233), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n804), .B1(new_n1010), .B2(new_n1042), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1221), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n978), .A2(new_n1074), .A3(new_n1001), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1074), .B1(new_n978), .B2(new_n1001), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(G390), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1221), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1263), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1265), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1273), .A3(new_n1220), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1268), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1262), .B1(new_n1276), .B2(KEYINPUT61), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(KEYINPUT127), .A3(new_n1278), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1261), .A2(KEYINPUT63), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT124), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1261), .B2(KEYINPUT63), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1147), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n673), .B1(new_n1284), .B2(new_n1140), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1196), .B1(new_n1285), .B2(new_n1170), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1283), .B(new_n1259), .C1(new_n1138), .C2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(KEYINPUT124), .A3(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1258), .A2(new_n1280), .A3(new_n1282), .A4(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1278), .B1(new_n1261), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1255), .B1(new_n1256), .B2(new_n1233), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT62), .B1(new_n1293), .B2(new_n1287), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1276), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(G405));
  OAI21_X1  g1096(.A(new_n1259), .B1(new_n1219), .B2(new_n1256), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1256), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1286), .A2(new_n1138), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1260), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1275), .ZN(G402));
endmodule


