//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT10), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G146), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(new_n195), .ZN(new_n199));
  AOI21_X1  g013(.A(G146), .B1(new_n190), .B2(new_n192), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  OAI21_X1  g015(.A(G128), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(G107), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G104), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n213), .A3(new_n214), .A4(new_n206), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n203), .A2(new_n204), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n202), .A2(new_n199), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n216), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT80), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n188), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n194), .A2(G143), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n201), .B1(G143), .B2(new_n194), .ZN(new_n225));
  OAI22_X1  g039(.A1(new_n200), .A2(new_n224), .B1(new_n196), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n219), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n221), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n191), .A2(G143), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n194), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n224), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n193), .A2(new_n230), .A3(new_n195), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n229), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n193), .A2(new_n230), .A3(new_n195), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n190), .A2(new_n192), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n224), .B1(new_n241), .B2(new_n194), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n240), .B(KEYINPUT67), .C1(new_n242), .C2(new_n232), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n210), .A2(new_n213), .A3(new_n206), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G101), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n248), .A3(G101), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n228), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G137), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(G134), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT11), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI211_X1 g075(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n253), .C2(G134), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n257), .B(new_n265), .C1(new_n261), .C2(new_n262), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n223), .A2(new_n252), .A3(new_n268), .ZN(new_n269));
  OAI22_X1  g083(.A1(new_n217), .A2(new_n222), .B1(new_n227), .B2(new_n221), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT12), .B1(new_n270), .B2(new_n267), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n227), .A2(new_n221), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n204), .B1(new_n203), .B2(new_n216), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n220), .A2(KEYINPUT80), .A3(new_n221), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT12), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n275), .A2(new_n276), .A3(new_n268), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n269), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(G110), .B(G140), .ZN(new_n279));
  INV_X1    g093(.A(G953), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n280), .A2(G227), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT10), .B1(new_n273), .B2(new_n274), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n284), .A2(new_n267), .A3(new_n251), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n282), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n267), .B1(new_n284), .B2(new_n251), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G469), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n278), .A2(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT81), .B(G469), .C1(new_n292), .C2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n269), .A2(new_n287), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n282), .ZN(new_n295));
  INV_X1    g109(.A(new_n282), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n269), .A2(KEYINPUT82), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n270), .A2(KEYINPUT12), .A3(new_n267), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n276), .B1(new_n275), .B2(new_n268), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT82), .B1(new_n269), .B2(new_n296), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT73), .B(G902), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n290), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n291), .A2(new_n293), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  XNOR2_X1  g123(.A(G110), .B(G122), .ZN(new_n310));
  XOR2_X1   g124(.A(G116), .B(G119), .Z(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT2), .B(G113), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n312), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n247), .A3(new_n249), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT5), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G116), .ZN(new_n319));
  OAI211_X1 g133(.A(G113), .B(new_n319), .C1(new_n311), .C2(new_n317), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n221), .A2(new_n313), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n310), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT6), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT6), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n316), .A2(new_n310), .A3(new_n321), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n316), .A2(new_n321), .A3(KEYINPUT83), .A4(new_n310), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n323), .B1(new_n329), .B2(new_n322), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT85), .B(G224), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n280), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT86), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT84), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n240), .B1(new_n242), .B2(new_n232), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(G125), .B2(new_n227), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n334), .B(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(KEYINPUT7), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n337), .A2(new_n340), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n310), .B(KEYINPUT8), .Z(new_n343));
  NAND2_X1  g157(.A1(new_n320), .A2(new_n313), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n216), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n345), .B2(new_n321), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n341), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n327), .A2(new_n328), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n309), .B1(new_n339), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n339), .A2(new_n309), .A3(new_n349), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n308), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT9), .B(G234), .ZN(new_n354));
  OAI21_X1  g168(.A(G221), .B1(new_n354), .B2(G902), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n355), .B(KEYINPUT79), .Z(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n306), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G902), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT93), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n280), .A3(G214), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT87), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT64), .B(G143), .ZN(new_n365));
  NOR2_X1   g179(.A1(G237), .A2(G953), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT87), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G214), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(G143), .A3(G214), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n364), .A2(KEYINPUT88), .A3(new_n365), .A4(new_n368), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G131), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n371), .A2(new_n265), .A3(new_n372), .A4(new_n373), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n361), .B1(new_n377), .B2(KEYINPUT17), .ZN(new_n378));
  INV_X1    g192(.A(new_n375), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT16), .ZN(new_n382));
  INV_X1    g196(.A(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G125), .ZN(new_n384));
  INV_X1    g198(.A(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G140), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT76), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n382), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G146), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n382), .B(new_n194), .C1(new_n387), .C2(new_n388), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(KEYINPUT77), .A3(G146), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n379), .A2(KEYINPUT17), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT17), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n375), .A2(KEYINPUT93), .A3(new_n396), .A4(new_n376), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n378), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G113), .B(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n205), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT18), .A2(G131), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n367), .B1(new_n366), .B2(G214), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n241), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT88), .B1(new_n404), .B2(new_n368), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n373), .A2(new_n372), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n371), .A2(new_n401), .A3(new_n372), .A4(new_n373), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n384), .A2(new_n386), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G146), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n380), .A2(new_n194), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n374), .A2(new_n402), .B1(new_n411), .B2(new_n410), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT89), .A3(new_n408), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n398), .A2(new_n400), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n400), .B1(new_n398), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n360), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G475), .ZN(new_n422));
  NOR2_X1   g236(.A1(G475), .A2(G902), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n409), .B1(new_n424), .B2(KEYINPUT19), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n409), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(G146), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(G146), .B2(new_n389), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n377), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT89), .B1(new_n416), .B2(new_n408), .ZN(new_n431));
  AND4_X1   g245(.A1(KEYINPUT89), .A2(new_n407), .A3(new_n408), .A4(new_n412), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT91), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n436));
  INV_X1    g250(.A(new_n400), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT91), .B(new_n430), .C1(new_n431), .C2(new_n432), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n398), .A2(new_n400), .A3(new_n418), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n415), .A2(new_n417), .B1(new_n377), .B2(new_n429), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n400), .B1(new_n442), .B2(KEYINPUT91), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n436), .B1(new_n443), .B2(new_n435), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n423), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT94), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT20), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(KEYINPUT20), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n438), .A2(new_n437), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT91), .B1(new_n418), .B2(new_n430), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT92), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n440), .A3(new_n439), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n454), .A2(new_n446), .A3(KEYINPUT20), .A4(new_n423), .ZN(new_n455));
  INV_X1    g269(.A(G952), .ZN(new_n456));
  AOI211_X1 g270(.A(G953), .B(new_n456), .C1(G234), .C2(G237), .ZN(new_n457));
  AOI211_X1 g271(.A(new_n280), .B(new_n304), .C1(G234), .C2(G237), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(G898), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AND4_X1   g275(.A1(new_n422), .A2(new_n450), .A3(new_n455), .A4(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(KEYINPUT95), .A2(G122), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT95), .A2(G122), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G116), .ZN(new_n466));
  INV_X1    g280(.A(G122), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G116), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n466), .A2(new_n212), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G116), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n463), .B2(new_n464), .ZN(new_n472));
  OAI21_X1  g286(.A(G107), .B1(new_n472), .B2(new_n468), .ZN(new_n473));
  AND2_X1   g287(.A1(KEYINPUT14), .A2(G107), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n470), .A2(new_n473), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  AND4_X1   g289(.A1(KEYINPUT14), .A2(new_n466), .A3(G107), .A4(new_n469), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT96), .B1(new_n241), .B2(new_n196), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT96), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n365), .A2(new_n479), .A3(G128), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n196), .A2(G143), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n481), .A2(new_n255), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n255), .B1(new_n481), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT97), .B1(new_n477), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n475), .A2(new_n476), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT97), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n487), .B(new_n488), .C1(new_n483), .C2(new_n484), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n255), .A3(new_n482), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n470), .A2(new_n473), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT13), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n481), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n478), .A2(KEYINPUT13), .A3(new_n480), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n494), .A2(new_n482), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n491), .B(new_n492), .C1(new_n496), .C2(new_n255), .ZN(new_n497));
  INV_X1    g311(.A(G217), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n354), .A2(new_n498), .A3(G953), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n490), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n490), .B2(new_n497), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n304), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G478), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n490), .A2(new_n497), .ZN(new_n506));
  INV_X1    g320(.A(new_n499), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n490), .A2(new_n497), .A3(new_n499), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n504), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n304), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT98), .B1(new_n462), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n450), .A2(new_n422), .A3(new_n455), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT98), .ZN(new_n517));
  NOR4_X1   g331(.A1(new_n516), .A2(new_n517), .A3(new_n513), .A4(new_n460), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n359), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT99), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(KEYINPUT99), .B(new_n359), .C1(new_n515), .C2(new_n518), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n280), .A2(G221), .A3(G234), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n196), .A2(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n318), .A2(G128), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT24), .B(G110), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n531));
  OAI211_X1 g345(.A(G119), .B(new_n196), .C1(new_n531), .C2(KEYINPUT23), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(KEYINPUT74), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n318), .B2(G128), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n536), .A2(KEYINPUT75), .ZN(new_n537));
  INV_X1    g351(.A(G110), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n536), .B2(KEYINPUT75), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n530), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n393), .A2(new_n540), .A3(new_n394), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n528), .A2(new_n529), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n536), .B2(G110), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n390), .A2(new_n411), .A3(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n541), .A2(KEYINPUT78), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT78), .B1(new_n541), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n525), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n525), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n541), .A2(new_n544), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT78), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n498), .B1(new_n304), .B2(G234), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n557));
  INV_X1    g371(.A(new_n304), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n547), .A2(KEYINPUT25), .A3(new_n304), .A4(new_n551), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n556), .B1(new_n561), .B2(new_n553), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n366), .A2(G210), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT27), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT26), .B(G101), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n255), .A2(G137), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n253), .A2(G134), .ZN(new_n569));
  OAI21_X1  g383(.A(G131), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT66), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(KEYINPUT66), .B(G131), .C1(new_n568), .C2(new_n569), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n226), .A2(new_n219), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n266), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n268), .B2(new_n335), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(KEYINPUT71), .A3(new_n315), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT69), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n315), .B(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n267), .A2(new_n239), .A3(new_n243), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n575), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT71), .B1(new_n576), .B2(new_n315), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT28), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(new_n575), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n315), .B(KEYINPUT69), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT28), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n567), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(KEYINPUT30), .A3(new_n575), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT30), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n572), .A2(new_n573), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n227), .A2(new_n593), .A3(new_n266), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n335), .B1(new_n264), .B2(new_n266), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT68), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n591), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n580), .A2(KEYINPUT68), .A3(KEYINPUT30), .A4(new_n575), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n315), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT70), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n567), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n581), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT31), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n587), .B1(new_n600), .B2(new_n315), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(KEYINPUT31), .A3(new_n604), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n590), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(G472), .A2(G902), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT32), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n584), .A2(new_n589), .ZN(new_n614));
  INV_X1    g428(.A(new_n567), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT31), .B1(new_n608), .B2(new_n604), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n598), .A2(new_n599), .B1(new_n313), .B2(new_n314), .ZN(new_n618));
  NOR4_X1   g432(.A1(new_n618), .A2(new_n606), .A3(new_n587), .A4(new_n603), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT32), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n621), .A3(new_n611), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n614), .A2(new_n567), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n608), .A2(new_n615), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT29), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT72), .B1(new_n585), .B2(new_n586), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n581), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT28), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n589), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n567), .A2(KEYINPUT29), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n304), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(G472), .B1(new_n626), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n563), .B1(new_n623), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n521), .A2(new_n522), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND2_X1  g450(.A1(new_n607), .A2(new_n609), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n558), .B1(new_n637), .B2(new_n616), .ZN(new_n638));
  INV_X1    g452(.A(G472), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n610), .A2(new_n612), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND4_X1   g456(.A1(new_n357), .A2(new_n642), .A3(new_n306), .A4(new_n562), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n558), .A2(new_n503), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n510), .A2(KEYINPUT33), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n508), .B2(new_n509), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n502), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT100), .B(G478), .Z(new_n650));
  OAI21_X1  g464(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n516), .A2(new_n461), .A3(new_n353), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n643), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NAND2_X1  g470(.A1(new_n353), .A2(new_n513), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n516), .A2(new_n460), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n643), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT35), .B(G107), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT101), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(G9));
  NAND2_X1  g476(.A1(new_n561), .A2(new_n553), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n549), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n554), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n642), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n521), .A2(new_n522), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  INV_X1    g487(.A(new_n667), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n623), .B2(new_n633), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n457), .B1(new_n458), .B2(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n516), .A2(new_n514), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n678), .A3(new_n359), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XOR2_X1   g494(.A(new_n677), .B(KEYINPUT39), .Z(new_n681));
  NAND3_X1  g495(.A1(new_n306), .A2(new_n357), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT40), .Z(new_n683));
  OAI21_X1  g497(.A(new_n567), .B1(new_n618), .B2(new_n587), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AOI211_X1 g499(.A(G902), .B(new_n685), .C1(new_n615), .C2(new_n628), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n623), .B1(new_n639), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n352), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n350), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT38), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n690), .A2(new_n514), .A3(new_n308), .A4(new_n667), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n683), .A2(new_n516), .A3(new_n687), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n241), .ZN(G45));
  INV_X1    g507(.A(new_n677), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n516), .A2(new_n651), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n675), .A3(new_n359), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  AND3_X1   g511(.A1(new_n620), .A2(new_n621), .A3(new_n611), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n621), .B1(new_n620), .B2(new_n611), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n633), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n305), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n290), .B1(new_n303), .B2(new_n304), .ZN(new_n702));
  INV_X1    g516(.A(new_n355), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n562), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n652), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT41), .B(G113), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  INV_X1    g522(.A(new_n449), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n447), .B(new_n709), .C1(new_n454), .C2(new_n423), .ZN(new_n710));
  INV_X1    g524(.A(new_n455), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n307), .B1(new_n688), .B2(new_n350), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n514), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n712), .A2(new_n422), .A3(new_n461), .A4(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT103), .B1(new_n705), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n658), .A2(new_n634), .A3(new_n717), .A4(new_n704), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  INV_X1    g534(.A(new_n702), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(new_n353), .A3(new_n355), .A4(new_n305), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n675), .B(new_n723), .C1(new_n515), .C2(new_n518), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NAND2_X1  g539(.A1(new_n620), .A2(new_n304), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n627), .B(new_n587), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n588), .B1(new_n727), .B2(KEYINPUT28), .ZN(new_n728));
  OAI22_X1  g542(.A1(new_n617), .A2(new_n619), .B1(new_n728), .B2(new_n567), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n726), .A2(G472), .B1(new_n611), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n704), .A3(new_n461), .A4(new_n562), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n516), .A2(new_n714), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n467), .ZN(G24));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n611), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n667), .B(new_n735), .C1(new_n638), .C2(new_n639), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n695), .A2(new_n723), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT104), .B(G125), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G27));
  NOR3_X1   g554(.A1(new_n688), .A2(new_n308), .A3(new_n350), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n289), .A2(new_n290), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n355), .B(new_n741), .C1(new_n701), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n695), .A2(new_n634), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(KEYINPUT42), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n695), .A2(new_n634), .A3(new_n744), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND3_X1  g568(.A1(new_n678), .A2(new_n634), .A3(new_n744), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n283), .A2(new_n288), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n290), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  OAI22_X1  g575(.A1(new_n760), .A2(new_n761), .B1(new_n759), .B2(new_n758), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n290), .A2(new_n360), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n757), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI221_X1 g580(.A(KEYINPUT46), .B1(new_n290), .B2(new_n360), .C1(new_n762), .C2(new_n763), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n305), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n355), .A3(new_n681), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n516), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n651), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n649), .A2(new_n650), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n645), .A2(new_n647), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n776), .B1(new_n777), .B2(new_n644), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n779));
  OAI22_X1  g593(.A1(new_n516), .A2(new_n778), .B1(KEYINPUT108), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n667), .B1(new_n640), .B2(new_n641), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT44), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n771), .A2(new_n741), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  NAND2_X1  g601(.A1(new_n768), .A2(new_n355), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n768), .A2(KEYINPUT47), .A3(new_n355), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n516), .A2(new_n651), .A3(new_n694), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n351), .A2(new_n307), .A3(new_n352), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n793), .A2(new_n700), .A3(new_n562), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n792), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  OR2_X1    g615(.A1(new_n687), .A2(new_n563), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n690), .A2(new_n307), .A3(new_n357), .A4(new_n651), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n721), .A2(new_n305), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT49), .ZN(new_n805));
  OR4_X1    g619(.A1(new_n516), .A2(new_n802), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  INV_X1    g621(.A(new_n457), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n775), .B2(new_n780), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n741), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n807), .B1(new_n811), .B2(new_n704), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n721), .A2(new_n355), .A3(new_n305), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n810), .A2(KEYINPUT112), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n737), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n704), .A2(new_n457), .A3(new_n741), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n802), .A2(new_n516), .A3(new_n651), .A4(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n735), .B(new_n562), .C1(new_n638), .C2(new_n639), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n813), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n809), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n690), .A2(new_n308), .ZN(new_n822));
  OR3_X1    g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n820), .B2(new_n822), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n817), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n815), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n815), .A2(new_n825), .A3(KEYINPUT113), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n790), .B(new_n791), .C1(new_n357), .C2(new_n804), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n810), .A2(new_n818), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n802), .A2(new_n816), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n772), .A2(new_n778), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n456), .B(G953), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n713), .B2(new_n820), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n634), .B1(new_n812), .B2(new_n814), .ZN(new_n839));
  NOR2_X1   g653(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n839), .B2(new_n841), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n838), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n817), .B1(new_n831), .B2(new_n832), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n823), .A2(KEYINPUT111), .A3(new_n824), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT111), .B1(new_n823), .B2(new_n824), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n846), .B(new_n815), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n830), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n834), .A2(new_n845), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n834), .A2(new_n845), .A3(new_n850), .A4(KEYINPUT115), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT110), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n705), .A2(new_n652), .B1(new_n731), .B2(new_n732), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n718), .B2(new_n716), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n857), .B2(new_n724), .ZN(new_n858));
  INV_X1    g672(.A(new_n856), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n855), .A2(new_n719), .A3(new_n859), .A4(new_n724), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n643), .B1(new_n653), .B2(new_n658), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n635), .A2(new_n671), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n732), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n355), .B1(new_n701), .B2(new_n742), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n667), .A3(new_n677), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n687), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n696), .A2(new_n679), .A3(new_n738), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT52), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n359), .B(new_n675), .C1(new_n695), .C2(new_n678), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n738), .A4(new_n867), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n736), .A2(new_n743), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n695), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n422), .A2(new_n505), .A3(new_n512), .A4(new_n694), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n794), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n877), .A2(new_n306), .A3(new_n357), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n675), .A2(new_n878), .A3(new_n712), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n755), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n753), .A2(KEYINPUT53), .A3(new_n875), .A4(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n861), .A2(new_n863), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n719), .A2(new_n859), .A3(new_n724), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n755), .A2(new_n879), .A3(new_n875), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n748), .B2(new_n752), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n887), .A3(new_n869), .A4(new_n872), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n635), .A2(new_n671), .A3(new_n862), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n883), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n888), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n863), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n884), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n893), .B1(new_n896), .B2(KEYINPUT54), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n853), .A2(new_n854), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n806), .B1(new_n898), .B2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n280), .A2(G952), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT118), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n304), .B(new_n309), .C1(new_n883), .C2(new_n890), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n330), .B(new_n338), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n902), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n903), .B2(KEYINPUT116), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n883), .A2(new_n890), .ZN(new_n910));
  INV_X1    g724(.A(new_n309), .ZN(new_n911));
  AND4_X1   g725(.A1(KEYINPUT116), .A2(new_n910), .A3(new_n558), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n905), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(KEYINPUT117), .B(new_n905), .C1(new_n909), .C2(new_n912), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(G51));
  XOR2_X1   g731(.A(new_n764), .B(KEYINPUT119), .Z(new_n918));
  AOI211_X1 g732(.A(new_n304), .B(new_n918), .C1(new_n883), .C2(new_n890), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n765), .B(KEYINPUT57), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n891), .B1(new_n883), .B2(new_n890), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n893), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n922), .B2(new_n303), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT120), .B1(new_n923), .B2(new_n901), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  INV_X1    g739(.A(new_n901), .ZN(new_n926));
  INV_X1    g740(.A(new_n303), .ZN(new_n927));
  INV_X1    g741(.A(new_n921), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n892), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n929), .B2(new_n920), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n925), .B(new_n926), .C1(new_n930), .C2(new_n919), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n931), .ZN(G54));
  AND4_X1   g746(.A1(KEYINPUT58), .A2(new_n910), .A3(G475), .A4(new_n558), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n926), .B1(new_n933), .B2(new_n454), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n454), .B2(new_n933), .ZN(G60));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n777), .B(KEYINPUT121), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n936), .B(new_n937), .C1(new_n897), .C2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n895), .A2(new_n884), .ZN(new_n942));
  INV_X1    g756(.A(new_n890), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT54), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n940), .B1(new_n944), .B2(new_n892), .ZN(new_n945));
  INV_X1    g759(.A(new_n937), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT123), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n902), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n937), .A2(new_n940), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n929), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n941), .A2(new_n947), .A3(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT60), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n910), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n948), .B1(new_n954), .B2(new_n552), .ZN(new_n955));
  INV_X1    g769(.A(new_n954), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT124), .B1(new_n956), .B2(new_n665), .ZN(new_n957));
  AND4_X1   g771(.A1(KEYINPUT124), .A2(new_n910), .A3(new_n665), .A4(new_n953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(KEYINPUT61), .B(new_n955), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G66));
  INV_X1    g777(.A(new_n459), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n280), .B1(new_n964), .B2(new_n331), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n863), .A2(new_n885), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n280), .ZN(new_n967));
  INV_X1    g781(.A(new_n330), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(G898), .B2(new_n280), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n967), .B(new_n969), .Z(G69));
  AND2_X1   g784(.A1(new_n870), .A2(new_n738), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n692), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  INV_X1    g787(.A(new_n634), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n974), .A2(new_n682), .A3(new_n794), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n516), .A2(new_n514), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n836), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT125), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n973), .A2(new_n800), .A3(new_n786), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n280), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n600), .B(new_n427), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n981), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n280), .A2(G900), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n971), .A2(new_n753), .A3(new_n755), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n974), .A2(new_n732), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n771), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n800), .A2(new_n987), .A3(new_n786), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n984), .B1(new_n988), .B2(new_n280), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n983), .B1(new_n989), .B2(KEYINPUT126), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n991), .B(new_n984), .C1(new_n988), .C2(new_n280), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n982), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n280), .B1(G227), .B2(G900), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n994), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n982), .B(new_n996), .C1(new_n990), .C2(new_n992), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n979), .B2(new_n966), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n901), .B1(new_n1001), .B2(new_n685), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n896), .A2(new_n625), .A3(new_n684), .A4(new_n1000), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1000), .B1(new_n988), .B2(new_n966), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n625), .B(KEYINPUT127), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1002), .A2(new_n1003), .A3(new_n1006), .ZN(G57));
endmodule


