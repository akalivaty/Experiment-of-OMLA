

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XNOR2_X1 U324 ( .A(n482), .B(KEYINPUT37), .ZN(n535) );
  XNOR2_X1 U325 ( .A(n461), .B(KEYINPUT121), .ZN(n570) );
  XOR2_X1 U326 ( .A(n350), .B(n349), .Z(n585) );
  XOR2_X1 U327 ( .A(KEYINPUT13), .B(KEYINPUT73), .Z(n292) );
  XOR2_X1 U328 ( .A(n448), .B(n447), .Z(n293) );
  AND2_X1 U329 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U330 ( .A(n442), .B(KEYINPUT55), .Z(n295) );
  INV_X1 U331 ( .A(G183GAT), .ZN(n451) );
  XNOR2_X1 U332 ( .A(n452), .B(n451), .ZN(n453) );
  AND2_X1 U333 ( .A1(n574), .A2(n441), .ZN(n442) );
  XNOR2_X1 U334 ( .A(n300), .B(n294), .ZN(n301) );
  XNOR2_X1 U335 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U336 ( .A(n302), .B(n301), .ZN(n303) );
  INV_X1 U337 ( .A(n459), .ZN(n460) );
  XNOR2_X1 U338 ( .A(n309), .B(n308), .ZN(n310) );
  AND2_X1 U339 ( .A1(n481), .A2(n495), .ZN(n482) );
  NAND2_X1 U340 ( .A1(n295), .A2(n460), .ZN(n461) );
  XNOR2_X1 U341 ( .A(n311), .B(n310), .ZN(n374) );
  INV_X1 U342 ( .A(G190GAT), .ZN(n491) );
  INV_X1 U343 ( .A(G50GAT), .ZN(n488) );
  XNOR2_X1 U344 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U345 ( .A(n488), .B(KEYINPUT112), .ZN(n489) );
  XNOR2_X1 U346 ( .A(n494), .B(n493), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n490), .B(n489), .ZN(G1331GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT76), .B(G92GAT), .Z(n297) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G71GAT), .Z(n448) );
  XOR2_X1 U350 ( .A(G176GAT), .B(G64GAT), .Z(n388) );
  XNOR2_X1 U351 ( .A(n448), .B(n388), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U353 ( .A(KEYINPUT32), .B(KEYINPUT79), .Z(n299) );
  XNOR2_X1 U354 ( .A(KEYINPUT33), .B(KEYINPUT77), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n303), .B(KEYINPUT31), .ZN(n311) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(G85GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(KEYINPUT75), .ZN(n312) );
  XOR2_X1 U359 ( .A(n312), .B(KEYINPUT78), .Z(n309) );
  XOR2_X1 U360 ( .A(G78GAT), .B(G148GAT), .Z(n306) );
  XNOR2_X1 U361 ( .A(G106GAT), .B(G204GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n401) );
  XNOR2_X1 U363 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n292), .B(n307), .ZN(n342) );
  XNOR2_X1 U365 ( .A(n401), .B(n342), .ZN(n308) );
  XOR2_X1 U366 ( .A(G134GAT), .B(KEYINPUT83), .Z(n421) );
  XOR2_X1 U367 ( .A(n312), .B(n421), .Z(n314) );
  NAND2_X1 U368 ( .A1(G232GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n316) );
  XNOR2_X1 U371 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U373 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n318) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U376 ( .A(n320), .B(n319), .Z(n324) );
  XNOR2_X1 U377 ( .A(G50GAT), .B(KEYINPUT80), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n321), .B(G162GAT), .ZN(n404) );
  XNOR2_X1 U379 ( .A(G36GAT), .B(G190GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n322), .B(G92GAT), .ZN(n385) );
  XNOR2_X1 U381 ( .A(n404), .B(n385), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U384 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n328) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G29GAT), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U387 ( .A(KEYINPUT7), .B(n329), .Z(n370) );
  XNOR2_X1 U388 ( .A(n330), .B(n370), .ZN(n496) );
  XOR2_X1 U389 ( .A(KEYINPUT36), .B(n496), .Z(n590) );
  XOR2_X1 U390 ( .A(KEYINPUT89), .B(KEYINPUT14), .Z(n332) );
  XNOR2_X1 U391 ( .A(KEYINPUT12), .B(KEYINPUT84), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n350) );
  XOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .Z(n384) );
  XOR2_X1 U394 ( .A(n384), .B(G211GAT), .Z(n334) );
  XOR2_X1 U395 ( .A(G22GAT), .B(G155GAT), .Z(n410) );
  XNOR2_X1 U396 ( .A(n410), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n346) );
  XOR2_X1 U398 ( .A(KEYINPUT86), .B(G64GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G127GAT), .B(G71GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U401 ( .A(KEYINPUT15), .B(KEYINPUT88), .Z(n338) );
  XNOR2_X1 U402 ( .A(KEYINPUT85), .B(KEYINPUT87), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U404 ( .A(n340), .B(n339), .Z(n344) );
  XNOR2_X1 U405 ( .A(G15GAT), .B(G1GAT), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n341), .B(KEYINPUT71), .ZN(n365) );
  XNOR2_X1 U407 ( .A(n365), .B(n342), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U409 ( .A(n346), .B(n345), .Z(n348) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  INV_X1 U412 ( .A(n585), .ZN(n495) );
  NOR2_X1 U413 ( .A1(n590), .A2(n495), .ZN(n351) );
  XOR2_X1 U414 ( .A(KEYINPUT45), .B(n351), .Z(n352) );
  NOR2_X1 U415 ( .A1(n374), .A2(n352), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n353), .B(KEYINPUT117), .ZN(n373) );
  XOR2_X1 U417 ( .A(G8GAT), .B(G113GAT), .Z(n355) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(G197GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U420 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n357) );
  XNOR2_X1 U421 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U423 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U424 ( .A(KEYINPUT68), .B(KEYINPUT72), .Z(n361) );
  NAND2_X1 U425 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U427 ( .A(KEYINPUT69), .B(n362), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U429 ( .A(G36GAT), .B(G50GAT), .Z(n367) );
  XNOR2_X1 U430 ( .A(G141GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U432 ( .A(n369), .B(n368), .Z(n372) );
  XNOR2_X1 U433 ( .A(n370), .B(G22GAT), .ZN(n371) );
  XOR2_X1 U434 ( .A(n372), .B(n371), .Z(n521) );
  INV_X1 U435 ( .A(n521), .ZN(n577) );
  NOR2_X1 U436 ( .A1(n373), .A2(n577), .ZN(n382) );
  INV_X1 U437 ( .A(KEYINPUT41), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n561) );
  NAND2_X1 U439 ( .A1(n577), .A2(n561), .ZN(n377) );
  INV_X1 U440 ( .A(KEYINPUT46), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n379) );
  INV_X1 U442 ( .A(n496), .ZN(n552) );
  NAND2_X1 U443 ( .A1(n495), .A2(n552), .ZN(n378) );
  NOR2_X1 U444 ( .A1(n379), .A2(n378), .ZN(n380) );
  XOR2_X1 U445 ( .A(n380), .B(KEYINPUT47), .Z(n381) );
  NOR2_X1 U446 ( .A1(n382), .A2(n381), .ZN(n383) );
  XOR2_X1 U447 ( .A(KEYINPUT48), .B(n383), .Z(n557) );
  XOR2_X1 U448 ( .A(n385), .B(n384), .Z(n390) );
  XOR2_X1 U449 ( .A(G211GAT), .B(KEYINPUT21), .Z(n387) );
  XNOR2_X1 U450 ( .A(G197GAT), .B(G218GAT), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n402) );
  XNOR2_X1 U452 ( .A(n402), .B(n388), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U454 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n392) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U457 ( .A(n394), .B(n393), .Z(n398) );
  XOR2_X1 U458 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n396) );
  XNOR2_X1 U459 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n450) );
  XNOR2_X1 U461 ( .A(n450), .B(G204GAT), .ZN(n397) );
  XOR2_X1 U462 ( .A(n398), .B(n397), .Z(n515) );
  INV_X1 U463 ( .A(n515), .ZN(n538) );
  NAND2_X1 U464 ( .A1(n557), .A2(n538), .ZN(n400) );
  XOR2_X1 U465 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n399) );
  XNOR2_X1 U466 ( .A(n400), .B(n399), .ZN(n574) );
  XOR2_X1 U467 ( .A(n402), .B(n401), .Z(n406) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n403) );
  XNOR2_X1 U469 ( .A(n403), .B(KEYINPUT2), .ZN(n422) );
  XNOR2_X1 U470 ( .A(n404), .B(n422), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n414) );
  XOR2_X1 U472 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n408) );
  XNOR2_X1 U473 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U475 ( .A(n410), .B(n409), .Z(n412) );
  NAND2_X1 U476 ( .A1(G228GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n470) );
  XOR2_X1 U479 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n416) );
  XNOR2_X1 U480 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U482 ( .A(KEYINPUT1), .B(n417), .Z(n419) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U485 ( .A(n420), .B(KEYINPUT97), .Z(n427) );
  XOR2_X1 U486 ( .A(n421), .B(G85GAT), .Z(n424) );
  XNOR2_X1 U487 ( .A(G162GAT), .B(n422), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(n425), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U491 ( .A(G148GAT), .B(G155GAT), .Z(n429) );
  XNOR2_X1 U492 ( .A(G29GAT), .B(G120GAT), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U494 ( .A(n431), .B(n430), .Z(n440) );
  XOR2_X1 U495 ( .A(KEYINPUT91), .B(KEYINPUT0), .Z(n433) );
  XNOR2_X1 U496 ( .A(KEYINPUT90), .B(G127GAT), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U498 ( .A(G113GAT), .B(n434), .Z(n458) );
  INV_X1 U499 ( .A(n458), .ZN(n438) );
  XOR2_X1 U500 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n436) );
  XNOR2_X1 U501 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n435) );
  XNOR2_X1 U502 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U503 ( .A(n438), .B(n437), .Z(n439) );
  XOR2_X1 U504 ( .A(n440), .B(n439), .Z(n536) );
  NOR2_X1 U505 ( .A1(n470), .A2(n536), .ZN(n441) );
  XOR2_X1 U506 ( .A(KEYINPUT92), .B(G176GAT), .Z(n444) );
  XNOR2_X1 U507 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n443) );
  XNOR2_X1 U508 ( .A(n444), .B(n443), .ZN(n456) );
  XOR2_X1 U509 ( .A(G134GAT), .B(G99GAT), .Z(n446) );
  XNOR2_X1 U510 ( .A(G43GAT), .B(G190GAT), .ZN(n445) );
  XNOR2_X1 U511 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U512 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n293), .B(n449), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n450), .B(KEYINPUT93), .ZN(n452) );
  XOR2_X1 U515 ( .A(n456), .B(n455), .Z(n457) );
  XOR2_X1 U516 ( .A(n458), .B(n457), .Z(n459) );
  NAND2_X1 U517 ( .A1(n570), .A2(n561), .ZN(n465) );
  XOR2_X1 U518 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n463) );
  XNOR2_X1 U519 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  XNOR2_X1 U522 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n466) );
  XOR2_X1 U523 ( .A(n466), .B(n470), .Z(n541) );
  INV_X1 U524 ( .A(n541), .ZN(n487) );
  INV_X1 U525 ( .A(KEYINPUT38), .ZN(n485) );
  NOR2_X1 U526 ( .A1(n459), .A2(n515), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n470), .A2(n467), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT25), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n469), .B(KEYINPUT105), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT104), .B(KEYINPUT26), .Z(n472) );
  NAND2_X1 U531 ( .A1(n459), .A2(n470), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n473), .B(KEYINPUT103), .ZN(n575) );
  XNOR2_X1 U534 ( .A(n515), .B(KEYINPUT27), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n575), .A2(n477), .ZN(n474) );
  NOR2_X1 U536 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U537 ( .A1(n536), .A2(n476), .ZN(n480) );
  INV_X1 U538 ( .A(n536), .ZN(n573) );
  NOR2_X1 U539 ( .A1(n477), .A2(n573), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n478), .B(KEYINPUT102), .ZN(n556) );
  NAND2_X1 U541 ( .A1(n556), .A2(n487), .ZN(n546) );
  NOR2_X1 U542 ( .A1(n546), .A2(n460), .ZN(n479) );
  NOR2_X1 U543 ( .A1(n480), .A2(n479), .ZN(n498) );
  NOR2_X1 U544 ( .A1(n590), .A2(n498), .ZN(n481) );
  INV_X1 U545 ( .A(n374), .ZN(n483) );
  NAND2_X1 U546 ( .A1(n577), .A2(n483), .ZN(n501) );
  NOR2_X1 U547 ( .A1(n535), .A2(n501), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U549 ( .A(KEYINPUT110), .B(n486), .ZN(n517) );
  NOR2_X1 U550 ( .A1(n487), .A2(n517), .ZN(n490) );
  NAND2_X1 U551 ( .A1(n570), .A2(n496), .ZN(n494) );
  XOR2_X1 U552 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT107), .B(KEYINPUT34), .Z(n504) );
  NOR2_X1 U554 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(KEYINPUT16), .ZN(n500) );
  INV_X1 U556 ( .A(n498), .ZN(n499) );
  NAND2_X1 U557 ( .A1(n500), .A2(n499), .ZN(n522) );
  NOR2_X1 U558 ( .A1(n501), .A2(n522), .ZN(n502) );
  XNOR2_X1 U559 ( .A(KEYINPUT106), .B(n502), .ZN(n511) );
  NAND2_X1 U560 ( .A1(n511), .A2(n536), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U562 ( .A(G1GAT), .B(n505), .ZN(G1324GAT) );
  NAND2_X1 U563 ( .A1(n511), .A2(n538), .ZN(n506) );
  XNOR2_X1 U564 ( .A(n506), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT35), .B(KEYINPUT109), .Z(n508) );
  NAND2_X1 U566 ( .A1(n511), .A2(n460), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n508), .B(n507), .ZN(n510) );
  XOR2_X1 U568 ( .A(G15GAT), .B(KEYINPUT108), .Z(n509) );
  XNOR2_X1 U569 ( .A(n510), .B(n509), .ZN(G1326GAT) );
  NAND2_X1 U570 ( .A1(n511), .A2(n541), .ZN(n512) );
  XNOR2_X1 U571 ( .A(n512), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U572 ( .A1(n573), .A2(n517), .ZN(n513) );
  XNOR2_X1 U573 ( .A(n513), .B(KEYINPUT39), .ZN(n514) );
  XNOR2_X1 U574 ( .A(G29GAT), .B(n514), .ZN(G1328GAT) );
  NOR2_X1 U575 ( .A1(n515), .A2(n517), .ZN(n516) );
  XOR2_X1 U576 ( .A(G36GAT), .B(n516), .Z(G1329GAT) );
  NOR2_X1 U577 ( .A1(n517), .A2(n459), .ZN(n519) );
  XNOR2_X1 U578 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n518) );
  XNOR2_X1 U579 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U580 ( .A(G43GAT), .B(n520), .ZN(G1330GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n525) );
  NAND2_X1 U582 ( .A1(n561), .A2(n521), .ZN(n534) );
  NOR2_X1 U583 ( .A1(n522), .A2(n534), .ZN(n523) );
  XOR2_X1 U584 ( .A(KEYINPUT113), .B(n523), .Z(n531) );
  NAND2_X1 U585 ( .A1(n531), .A2(n536), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U587 ( .A(G57GAT), .B(n526), .Z(G1332GAT) );
  XOR2_X1 U588 ( .A(G64GAT), .B(KEYINPUT115), .Z(n528) );
  NAND2_X1 U589 ( .A1(n531), .A2(n538), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n528), .B(n527), .ZN(G1333GAT) );
  NAND2_X1 U591 ( .A1(n460), .A2(n531), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n529), .B(KEYINPUT116), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G71GAT), .B(n530), .ZN(G1334GAT) );
  XOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT43), .Z(n533) );
  NAND2_X1 U595 ( .A1(n531), .A2(n541), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1335GAT) );
  NOR2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n542), .A2(n536), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n537), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n542), .A2(n538), .ZN(n539) );
  XNOR2_X1 U601 ( .A(n539), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n460), .A2(n542), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(KEYINPUT44), .ZN(n544) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(n544), .ZN(G1339GAT) );
  NAND2_X1 U607 ( .A1(n557), .A2(n460), .ZN(n545) );
  NOR2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n553), .A2(n577), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U612 ( .A1(n553), .A2(n561), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  NAND2_X1 U614 ( .A1(n553), .A2(n585), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(KEYINPUT50), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U618 ( .A1(n553), .A2(n496), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U621 ( .A1(n575), .A2(n558), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n567), .A2(n577), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n559), .B(KEYINPUT118), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n563) );
  NAND2_X1 U626 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT119), .Z(n564) );
  XNOR2_X1 U629 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n567), .A2(n585), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n496), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n570), .A2(n577), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(G183GAT), .B(KEYINPUT123), .Z(n572) );
  NAND2_X1 U637 ( .A1(n570), .A2(n585), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n588) );
  NAND2_X1 U642 ( .A1(n588), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n581) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n583) );
  NAND2_X1 U647 ( .A1(n588), .A2(n374), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  INV_X1 U653 ( .A(n588), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

