

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724;

  NOR2_X1 U373 ( .A1(n661), .A2(n548), .ZN(n534) );
  INV_X1 U374 ( .A(G953), .ZN(n714) );
  INV_X2 U375 ( .A(n490), .ZN(n487) );
  NOR2_X2 U376 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X2 U377 ( .A(n537), .B(KEYINPUT1), .ZN(n659) );
  XNOR2_X1 U378 ( .A(n431), .B(n430), .ZN(n528) );
  NOR2_X1 U379 ( .A1(n723), .A2(n720), .ZN(n542) );
  OR2_X2 U380 ( .A1(n528), .A2(n433), .ZN(n547) );
  XNOR2_X1 U381 ( .A(n408), .B(G472), .ZN(n525) );
  NAND2_X1 U382 ( .A1(n588), .A2(n712), .ZN(n649) );
  XNOR2_X2 U383 ( .A(n410), .B(KEYINPUT33), .ZN(n688) );
  XNOR2_X2 U384 ( .A(n443), .B(KEYINPUT0), .ZN(n490) );
  AND2_X1 U385 ( .A1(n559), .A2(n558), .ZN(n571) );
  XNOR2_X1 U386 ( .A(n357), .B(G131), .ZN(n358) );
  XNOR2_X1 U387 ( .A(G134), .B(G137), .ZN(n357) );
  XNOR2_X1 U388 ( .A(n707), .B(G146), .ZN(n402) );
  XNOR2_X1 U389 ( .A(n530), .B(KEYINPUT39), .ZN(n584) );
  XNOR2_X1 U390 ( .A(n456), .B(n351), .ZN(n457) );
  OR2_X1 U391 ( .A1(n607), .A2(G902), .ZN(n456) );
  AND2_X1 U392 ( .A1(n594), .A2(G953), .ZN(n705) );
  XNOR2_X1 U393 ( .A(n397), .B(n396), .ZN(n412) );
  XNOR2_X1 U394 ( .A(G140), .B(KEYINPUT10), .ZN(n371) );
  XNOR2_X1 U395 ( .A(n508), .B(KEYINPUT45), .ZN(n588) );
  XNOR2_X1 U396 ( .A(n387), .B(KEYINPUT25), .ZN(n388) );
  XNOR2_X1 U397 ( .A(n386), .B(KEYINPUT77), .ZN(n387) );
  INV_X1 U398 ( .A(KEYINPUT69), .ZN(n367) );
  XNOR2_X1 U399 ( .A(n402), .B(n401), .ZN(n407) );
  XNOR2_X1 U400 ( .A(n381), .B(n380), .ZN(n466) );
  XNOR2_X1 U401 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U402 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n377) );
  BUF_X1 U403 ( .A(n478), .Z(n664) );
  XNOR2_X1 U404 ( .A(n532), .B(n531), .ZN(n723) );
  INV_X1 U405 ( .A(KEYINPUT40), .ZN(n531) );
  NOR2_X1 U406 ( .A1(n545), .A2(n544), .ZN(n638) );
  XNOR2_X1 U407 ( .A(n593), .B(n592), .ZN(n595) );
  XOR2_X1 U408 ( .A(n451), .B(n706), .Z(n350) );
  XOR2_X1 U409 ( .A(KEYINPUT96), .B(KEYINPUT13), .Z(n351) );
  AND2_X1 U410 ( .A1(n539), .A2(n475), .ZN(n352) );
  AND2_X1 U411 ( .A1(n638), .A2(n546), .ZN(n353) );
  INV_X1 U412 ( .A(KEYINPUT70), .ZN(n395) );
  XNOR2_X1 U413 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U414 ( .A(n412), .B(n398), .ZN(n400) );
  XNOR2_X1 U415 ( .A(n400), .B(n399), .ZN(n401) );
  INV_X1 U416 ( .A(KEYINPUT68), .ZN(n378) );
  INV_X1 U417 ( .A(KEYINPUT34), .ZN(n444) );
  NOR2_X1 U418 ( .A1(n495), .A2(n493), .ZN(n539) );
  XNOR2_X1 U419 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U420 ( .A(n367), .B(G469), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n424), .B(n358), .ZN(n707) );
  BUF_X1 U422 ( .A(n588), .Z(n651) );
  BUF_X1 U423 ( .A(n528), .Z(n581) );
  XNOR2_X1 U424 ( .A(n591), .B(KEYINPUT118), .ZN(n592) );
  OR2_X2 U425 ( .A1(n483), .A2(n477), .ZN(n500) );
  XNOR2_X1 U426 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U427 ( .A(n519), .B(n518), .ZN(G69) );
  NAND2_X1 U428 ( .A1(G953), .A2(G224), .ZN(n354) );
  XNOR2_X1 U429 ( .A(KEYINPUT61), .B(n354), .ZN(n355) );
  NAND2_X1 U430 ( .A1(n355), .A2(G898), .ZN(n356) );
  XNOR2_X1 U431 ( .A(KEYINPUT119), .B(n356), .ZN(n511) );
  XNOR2_X2 U432 ( .A(G143), .B(G128), .ZN(n461) );
  XNOR2_X1 U433 ( .A(n461), .B(KEYINPUT4), .ZN(n424) );
  XNOR2_X1 U434 ( .A(G140), .B(KEYINPUT89), .ZN(n365) );
  XOR2_X1 U435 ( .A(KEYINPUT78), .B(G107), .Z(n360) );
  XNOR2_X1 U436 ( .A(G101), .B(G104), .ZN(n359) );
  XNOR2_X1 U437 ( .A(n360), .B(n359), .ZN(n363) );
  XNOR2_X1 U438 ( .A(KEYINPUT75), .B(G110), .ZN(n414) );
  NAND2_X1 U439 ( .A1(G227), .A2(n714), .ZN(n361) );
  XNOR2_X1 U440 ( .A(n414), .B(n361), .ZN(n362) );
  XNOR2_X1 U441 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U442 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U443 ( .A(n402), .B(n366), .ZN(n695) );
  NOR2_X1 U444 ( .A1(G902), .A2(n695), .ZN(n369) );
  XNOR2_X2 U445 ( .A(n369), .B(n368), .ZN(n537) );
  INV_X2 U446 ( .A(G146), .ZN(n370) );
  XNOR2_X2 U447 ( .A(n370), .B(G125), .ZN(n421) );
  XNOR2_X2 U448 ( .A(n421), .B(n371), .ZN(n706) );
  XNOR2_X1 U449 ( .A(n706), .B(KEYINPUT23), .ZN(n376) );
  XOR2_X1 U450 ( .A(G110), .B(G119), .Z(n373) );
  XNOR2_X1 U451 ( .A(G128), .B(G137), .ZN(n372) );
  XNOR2_X1 U452 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U453 ( .A(n374), .B(KEYINPUT24), .Z(n375) );
  XNOR2_X1 U454 ( .A(n376), .B(n375), .ZN(n383) );
  XNOR2_X1 U455 ( .A(n377), .B(KEYINPUT81), .ZN(n381) );
  NAND2_X1 U456 ( .A1(G234), .A2(n714), .ZN(n379) );
  AND2_X1 U457 ( .A1(n466), .A2(G221), .ZN(n382) );
  XNOR2_X1 U458 ( .A(n383), .B(n382), .ZN(n703) );
  NOR2_X1 U459 ( .A1(G902), .A2(n703), .ZN(n389) );
  XNOR2_X1 U460 ( .A(KEYINPUT15), .B(G902), .ZN(n589) );
  NAND2_X1 U461 ( .A1(n589), .A2(G234), .ZN(n385) );
  XNOR2_X1 U462 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n384) );
  XNOR2_X1 U463 ( .A(n385), .B(n384), .ZN(n390) );
  NAND2_X1 U464 ( .A1(G217), .A2(n390), .ZN(n386) );
  XNOR2_X1 U465 ( .A(n389), .B(n388), .ZN(n478) );
  AND2_X1 U466 ( .A1(n390), .A2(G221), .ZN(n392) );
  INV_X1 U467 ( .A(KEYINPUT21), .ZN(n391) );
  XNOR2_X1 U468 ( .A(n392), .B(n391), .ZN(n663) );
  NOR2_X1 U469 ( .A1(n478), .A2(n663), .ZN(n393) );
  XNOR2_X1 U470 ( .A(n393), .B(KEYINPUT65), .ZN(n658) );
  NOR2_X1 U471 ( .A1(n659), .A2(n658), .ZN(n394) );
  XNOR2_X1 U472 ( .A(n394), .B(KEYINPUT72), .ZN(n486) );
  XNOR2_X1 U473 ( .A(n395), .B(KEYINPUT3), .ZN(n397) );
  XNOR2_X1 U474 ( .A(G119), .B(G101), .ZN(n396) );
  XOR2_X1 U475 ( .A(KEYINPUT5), .B(KEYINPUT73), .Z(n398) );
  INV_X1 U476 ( .A(KEYINPUT74), .ZN(n399) );
  NOR2_X1 U477 ( .A1(G237), .A2(G953), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n403), .B(KEYINPUT76), .ZN(n452) );
  AND2_X1 U479 ( .A1(n452), .A2(G210), .ZN(n405) );
  XNOR2_X1 U480 ( .A(G113), .B(G116), .ZN(n404) );
  XNOR2_X1 U481 ( .A(n407), .B(n406), .ZN(n599) );
  INV_X1 U482 ( .A(G902), .ZN(n429) );
  NAND2_X1 U483 ( .A1(n599), .A2(n429), .ZN(n408) );
  XNOR2_X1 U484 ( .A(KEYINPUT101), .B(KEYINPUT6), .ZN(n409) );
  XNOR2_X1 U485 ( .A(n525), .B(n409), .ZN(n477) );
  AND2_X2 U486 ( .A1(n486), .A2(n477), .ZN(n410) );
  XNOR2_X1 U487 ( .A(G122), .B(G113), .ZN(n411) );
  XNOR2_X1 U488 ( .A(n411), .B(G104), .ZN(n451) );
  XNOR2_X1 U489 ( .A(n412), .B(n451), .ZN(n418) );
  XNOR2_X1 U490 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n413) );
  XNOR2_X1 U491 ( .A(n414), .B(n413), .ZN(n416) );
  INV_X1 U492 ( .A(G116), .ZN(n415) );
  XNOR2_X1 U493 ( .A(n415), .B(G107), .ZN(n460) );
  XNOR2_X1 U494 ( .A(n416), .B(n460), .ZN(n417) );
  XNOR2_X1 U495 ( .A(n418), .B(n417), .ZN(n512) );
  NAND2_X1 U496 ( .A1(n714), .A2(G224), .ZN(n419) );
  XNOR2_X1 U497 ( .A(n419), .B(KEYINPUT85), .ZN(n423) );
  XNOR2_X1 U498 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n420) );
  XNOR2_X1 U499 ( .A(n423), .B(n422), .ZN(n425) );
  XNOR2_X1 U500 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U501 ( .A(n512), .B(n426), .ZN(n613) );
  INV_X1 U502 ( .A(n589), .ZN(n427) );
  OR2_X2 U503 ( .A1(n613), .A2(n427), .ZN(n431) );
  INV_X1 U504 ( .A(G237), .ZN(n428) );
  NAND2_X1 U505 ( .A1(n429), .A2(n428), .ZN(n432) );
  NAND2_X1 U506 ( .A1(n432), .A2(G210), .ZN(n430) );
  NAND2_X1 U507 ( .A1(n432), .A2(G214), .ZN(n672) );
  INV_X1 U508 ( .A(n672), .ZN(n433) );
  XNOR2_X2 U509 ( .A(n547), .B(KEYINPUT19), .ZN(n543) );
  NAND2_X1 U510 ( .A1(G234), .A2(G237), .ZN(n434) );
  XNOR2_X1 U511 ( .A(n434), .B(KEYINPUT86), .ZN(n435) );
  XNOR2_X1 U512 ( .A(KEYINPUT14), .B(n435), .ZN(n438) );
  AND2_X1 U513 ( .A1(n438), .A2(G953), .ZN(n436) );
  NAND2_X1 U514 ( .A1(G902), .A2(n436), .ZN(n521) );
  NOR2_X1 U515 ( .A1(G898), .A2(n521), .ZN(n437) );
  XOR2_X1 U516 ( .A(KEYINPUT87), .B(n437), .Z(n439) );
  NAND2_X1 U517 ( .A1(G952), .A2(n438), .ZN(n686) );
  NOR2_X1 U518 ( .A1(G953), .A2(n686), .ZN(n523) );
  NOR2_X1 U519 ( .A1(n439), .A2(n523), .ZN(n441) );
  INV_X1 U520 ( .A(KEYINPUT88), .ZN(n440) );
  XNOR2_X1 U521 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U522 ( .A1(n543), .A2(n442), .ZN(n443) );
  NOR2_X1 U523 ( .A1(n688), .A2(n490), .ZN(n445) );
  XNOR2_X1 U524 ( .A(n445), .B(n444), .ZN(n473) );
  XOR2_X1 U525 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n447) );
  XNOR2_X1 U526 ( .A(KEYINPUT95), .B(KEYINPUT12), .ZN(n446) );
  XNOR2_X1 U527 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U528 ( .A(n448), .B(KEYINPUT11), .Z(n450) );
  XNOR2_X1 U529 ( .A(G131), .B(G143), .ZN(n449) );
  XNOR2_X1 U530 ( .A(n450), .B(n449), .ZN(n455) );
  NAND2_X1 U531 ( .A1(G214), .A2(n452), .ZN(n453) );
  XNOR2_X1 U532 ( .A(n350), .B(n453), .ZN(n454) );
  XOR2_X1 U533 ( .A(n455), .B(n454), .Z(n607) );
  XNOR2_X1 U534 ( .A(n457), .B(G475), .ZN(n495) );
  XOR2_X1 U535 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n459) );
  XNOR2_X1 U536 ( .A(G134), .B(G122), .ZN(n458) );
  XNOR2_X1 U537 ( .A(n459), .B(n458), .ZN(n465) );
  XOR2_X1 U538 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n463) );
  XNOR2_X1 U539 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U540 ( .A(n463), .B(n462), .Z(n464) );
  XOR2_X1 U541 ( .A(n465), .B(n464), .Z(n468) );
  NAND2_X1 U542 ( .A1(G217), .A2(n466), .ZN(n467) );
  XNOR2_X1 U543 ( .A(n468), .B(n467), .ZN(n591) );
  NOR2_X1 U544 ( .A1(G902), .A2(n591), .ZN(n470) );
  XNOR2_X1 U545 ( .A(KEYINPUT99), .B(G478), .ZN(n469) );
  XNOR2_X1 U546 ( .A(n470), .B(n469), .ZN(n493) );
  NAND2_X1 U547 ( .A1(n495), .A2(n493), .ZN(n471) );
  XNOR2_X1 U548 ( .A(n471), .B(KEYINPUT102), .ZN(n562) );
  XOR2_X1 U549 ( .A(n562), .B(KEYINPUT79), .Z(n472) );
  XNOR2_X1 U550 ( .A(n474), .B(KEYINPUT35), .ZN(n721) );
  INV_X1 U551 ( .A(n663), .ZN(n475) );
  NAND2_X1 U552 ( .A1(n487), .A2(n352), .ZN(n476) );
  XNOR2_X1 U553 ( .A(n476), .B(KEYINPUT22), .ZN(n483) );
  INV_X1 U554 ( .A(n659), .ZN(n482) );
  NAND2_X1 U555 ( .A1(n482), .A2(n664), .ZN(n479) );
  NOR2_X2 U556 ( .A1(n500), .A2(n479), .ZN(n481) );
  XNOR2_X1 U557 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n480) );
  XNOR2_X1 U558 ( .A(n481), .B(n480), .ZN(n598) );
  INV_X1 U559 ( .A(n664), .ZN(n498) );
  NOR2_X1 U560 ( .A1(n482), .A2(n498), .ZN(n578) );
  INV_X1 U561 ( .A(n525), .ZN(n661) );
  NAND2_X1 U562 ( .A1(n578), .A2(n661), .ZN(n484) );
  NOR2_X1 U563 ( .A1(n484), .A2(n483), .ZN(n596) );
  NOR2_X1 U564 ( .A1(n598), .A2(n596), .ZN(n485) );
  NAND2_X1 U565 ( .A1(n721), .A2(n485), .ZN(n505) );
  NAND2_X1 U566 ( .A1(n505), .A2(KEYINPUT44), .ZN(n503) );
  AND2_X1 U567 ( .A1(n486), .A2(n525), .ZN(n669) );
  NAND2_X1 U568 ( .A1(n669), .A2(n487), .ZN(n488) );
  XOR2_X1 U569 ( .A(KEYINPUT31), .B(n488), .Z(n643) );
  NOR2_X1 U570 ( .A1(n658), .A2(n537), .ZN(n489) );
  XNOR2_X1 U571 ( .A(n489), .B(KEYINPUT91), .ZN(n520) );
  NOR2_X1 U572 ( .A1(n520), .A2(n490), .ZN(n491) );
  XNOR2_X1 U573 ( .A(n491), .B(KEYINPUT92), .ZN(n492) );
  NAND2_X1 U574 ( .A1(n492), .A2(n661), .ZN(n626) );
  NAND2_X1 U575 ( .A1(n643), .A2(n626), .ZN(n497) );
  INV_X1 U576 ( .A(n493), .ZN(n494) );
  OR2_X1 U577 ( .A1(n495), .A2(n494), .ZN(n644) );
  AND2_X1 U578 ( .A1(n495), .A2(n494), .ZN(n637) );
  INV_X1 U579 ( .A(n637), .ZN(n640) );
  NAND2_X1 U580 ( .A1(n644), .A2(n640), .ZN(n496) );
  XNOR2_X1 U581 ( .A(KEYINPUT100), .B(n496), .ZN(n553) );
  AND2_X1 U582 ( .A1(n497), .A2(n553), .ZN(n501) );
  NAND2_X1 U583 ( .A1(n659), .A2(n498), .ZN(n499) );
  NOR2_X1 U584 ( .A1(n500), .A2(n499), .ZN(n621) );
  NOR2_X1 U585 ( .A1(n501), .A2(n621), .ZN(n502) );
  NAND2_X1 U586 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U587 ( .A(n504), .B(KEYINPUT83), .ZN(n507) );
  OR2_X1 U588 ( .A1(n505), .A2(KEYINPUT44), .ZN(n506) );
  NAND2_X1 U589 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U590 ( .A1(n651), .A2(n714), .ZN(n509) );
  XOR2_X1 U591 ( .A(KEYINPUT120), .B(n509), .Z(n510) );
  NOR2_X1 U592 ( .A1(n511), .A2(n510), .ZN(n519) );
  INV_X1 U593 ( .A(n512), .ZN(n514) );
  OR2_X1 U594 ( .A1(G898), .A2(n714), .ZN(n513) );
  NAND2_X1 U595 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U596 ( .A(n515), .B(KEYINPUT121), .ZN(n517) );
  INV_X1 U597 ( .A(KEYINPUT122), .ZN(n516) );
  XNOR2_X1 U598 ( .A(n520), .B(KEYINPUT104), .ZN(n524) );
  NOR2_X1 U599 ( .A1(G900), .A2(n521), .ZN(n522) );
  NOR2_X1 U600 ( .A1(n523), .A2(n522), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n524), .A2(n533), .ZN(n561) );
  INV_X1 U602 ( .A(KEYINPUT30), .ZN(n527) );
  NAND2_X1 U603 ( .A1(n525), .A2(n672), .ZN(n526) );
  XNOR2_X1 U604 ( .A(n527), .B(n526), .ZN(n560) );
  XNOR2_X1 U605 ( .A(n581), .B(KEYINPUT38), .ZN(n673) );
  AND2_X1 U606 ( .A1(n560), .A2(n673), .ZN(n529) );
  NAND2_X1 U607 ( .A1(n561), .A2(n529), .ZN(n530) );
  NAND2_X1 U608 ( .A1(n584), .A2(n637), .ZN(n532) );
  INV_X1 U609 ( .A(KEYINPUT28), .ZN(n535) );
  NOR2_X1 U610 ( .A1(n663), .A2(n533), .ZN(n575) );
  NAND2_X1 U611 ( .A1(n664), .A2(n575), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n535), .B(n534), .ZN(n536) );
  NOR2_X1 U613 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U614 ( .A(KEYINPUT105), .B(n538), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n673), .A2(n672), .ZN(n677) );
  INV_X1 U616 ( .A(n539), .ZN(n675) );
  NOR2_X1 U617 ( .A1(n677), .A2(n675), .ZN(n540) );
  XNOR2_X1 U618 ( .A(KEYINPUT41), .B(n540), .ZN(n687) );
  NOR2_X1 U619 ( .A1(n545), .A2(n687), .ZN(n541) );
  XNOR2_X1 U620 ( .A(n541), .B(KEYINPUT42), .ZN(n720) );
  XNOR2_X1 U621 ( .A(n542), .B(KEYINPUT46), .ZN(n573) );
  INV_X1 U622 ( .A(n543), .ZN(n544) );
  NAND2_X1 U623 ( .A1(n553), .A2(KEYINPUT66), .ZN(n555) );
  NOR2_X1 U624 ( .A1(KEYINPUT47), .A2(n555), .ZN(n546) );
  NAND2_X1 U625 ( .A1(n477), .A2(n637), .ZN(n577) );
  INV_X1 U626 ( .A(n577), .ZN(n550) );
  NOR2_X1 U627 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U628 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U629 ( .A(KEYINPUT36), .B(n551), .ZN(n552) );
  NOR2_X1 U630 ( .A1(n659), .A2(n552), .ZN(n646) );
  NOR2_X1 U631 ( .A1(n353), .A2(n646), .ZN(n559) );
  INV_X1 U632 ( .A(KEYINPUT80), .ZN(n566) );
  INV_X1 U633 ( .A(n553), .ZN(n676) );
  NAND2_X1 U634 ( .A1(n566), .A2(n676), .ZN(n554) );
  NAND2_X1 U635 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U636 ( .A1(n638), .A2(n556), .ZN(n557) );
  NAND2_X1 U637 ( .A1(n557), .A2(KEYINPUT47), .ZN(n558) );
  NAND2_X1 U638 ( .A1(n676), .A2(KEYINPUT47), .ZN(n565) );
  AND2_X1 U639 ( .A1(n561), .A2(n560), .ZN(n564) );
  NOR2_X1 U640 ( .A1(n562), .A2(n581), .ZN(n563) );
  NAND2_X1 U641 ( .A1(n564), .A2(n563), .ZN(n636) );
  NAND2_X1 U642 ( .A1(n565), .A2(n636), .ZN(n567) );
  NAND2_X1 U643 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U644 ( .A1(n636), .A2(KEYINPUT80), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n569), .A2(n568), .ZN(n570) );
  AND2_X1 U646 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U647 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U648 ( .A(KEYINPUT48), .B(n574), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n575), .A2(n672), .ZN(n576) );
  NOR2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U652 ( .A(n580), .B(KEYINPUT43), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U654 ( .A(KEYINPUT103), .B(n583), .Z(n718) );
  INV_X1 U655 ( .A(n644), .ZN(n631) );
  AND2_X1 U656 ( .A1(n584), .A2(n631), .ZN(n648) );
  INV_X1 U657 ( .A(n648), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n718), .A2(n585), .ZN(n586) );
  NOR2_X2 U659 ( .A1(n587), .A2(n586), .ZN(n712) );
  XNOR2_X1 U660 ( .A(n649), .B(KEYINPUT2), .ZN(n590) );
  AND2_X2 U661 ( .A1(n590), .A2(n427), .ZN(n701) );
  NAND2_X1 U662 ( .A1(n701), .A2(G478), .ZN(n593) );
  INV_X1 U663 ( .A(G952), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n705), .ZN(G63) );
  XOR2_X1 U665 ( .A(G110), .B(n596), .Z(G12) );
  XNOR2_X1 U666 ( .A(G119), .B(KEYINPUT125), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n598), .B(n597), .ZN(G21) );
  NAND2_X1 U668 ( .A1(n701), .A2(G472), .ZN(n601) );
  XNOR2_X1 U669 ( .A(n599), .B(KEYINPUT62), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n601), .B(n600), .ZN(n602) );
  INV_X1 U671 ( .A(n705), .ZN(n617) );
  NAND2_X1 U672 ( .A1(n602), .A2(n617), .ZN(n604) );
  XNOR2_X1 U673 ( .A(KEYINPUT84), .B(KEYINPUT63), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n604), .B(n603), .ZN(G57) );
  NAND2_X1 U675 ( .A1(n701), .A2(G475), .ZN(n609) );
  XNOR2_X1 U676 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n605) );
  XOR2_X1 U677 ( .A(n605), .B(KEYINPUT59), .Z(n606) );
  XNOR2_X1 U678 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n610), .A2(n617), .ZN(n612) );
  INV_X1 U681 ( .A(KEYINPUT60), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n612), .B(n611), .ZN(G60) );
  NAND2_X1 U683 ( .A1(n701), .A2(G210), .ZN(n616) );
  XNOR2_X1 U684 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n613), .B(n614), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n620) );
  INV_X1 U688 ( .A(KEYINPUT56), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n620), .B(n619), .ZN(G51) );
  XOR2_X1 U690 ( .A(G101), .B(n621), .Z(G3) );
  NOR2_X1 U691 ( .A1(n640), .A2(n626), .ZN(n622) );
  XOR2_X1 U692 ( .A(KEYINPUT106), .B(n622), .Z(n623) );
  XNOR2_X1 U693 ( .A(G104), .B(n623), .ZN(G6) );
  XOR2_X1 U694 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n625) );
  XNOR2_X1 U695 ( .A(KEYINPUT107), .B(KEYINPUT27), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n630) );
  NOR2_X1 U697 ( .A1(n644), .A2(n626), .ZN(n628) );
  XNOR2_X1 U698 ( .A(G107), .B(KEYINPUT26), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(n629) );
  XOR2_X1 U700 ( .A(n630), .B(n629), .Z(G9) );
  XOR2_X1 U701 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n633) );
  NAND2_X1 U702 ( .A1(n638), .A2(n631), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U704 ( .A(G128), .B(n634), .ZN(G30) );
  XOR2_X1 U705 ( .A(G143), .B(KEYINPUT111), .Z(n635) );
  XNOR2_X1 U706 ( .A(n636), .B(n635), .ZN(G45) );
  NAND2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U708 ( .A(n639), .B(G146), .ZN(G48) );
  NOR2_X1 U709 ( .A1(n640), .A2(n643), .ZN(n641) );
  XOR2_X1 U710 ( .A(KEYINPUT112), .B(n641), .Z(n642) );
  XNOR2_X1 U711 ( .A(G113), .B(n642), .ZN(G15) );
  NOR2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U713 ( .A(G116), .B(n645), .Z(G18) );
  XNOR2_X1 U714 ( .A(G125), .B(n646), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U716 ( .A(G134), .B(n648), .Z(G36) );
  NAND2_X1 U717 ( .A1(n649), .A2(KEYINPUT2), .ZN(n653) );
  INV_X1 U718 ( .A(KEYINPUT2), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n656) );
  NOR2_X1 U721 ( .A1(n712), .A2(KEYINPUT2), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT82), .ZN(n655) );
  OR2_X1 U723 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n657), .A2(n714), .ZN(n693) );
  NAND2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U726 ( .A(n660), .B(KEYINPUT50), .ZN(n662) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n667) );
  NAND2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U729 ( .A(KEYINPUT49), .B(n665), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U731 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U732 ( .A(KEYINPUT51), .B(n670), .Z(n671) );
  NOR2_X1 U733 ( .A1(n687), .A2(n671), .ZN(n682) );
  NOR2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U735 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U736 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U737 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U738 ( .A1(n680), .A2(n688), .ZN(n681) );
  NOR2_X1 U739 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U740 ( .A(n683), .B(KEYINPUT113), .Z(n684) );
  XNOR2_X1 U741 ( .A(KEYINPUT52), .B(n684), .ZN(n685) );
  NOR2_X1 U742 ( .A1(n686), .A2(n685), .ZN(n690) );
  NOR2_X1 U743 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U744 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U745 ( .A(KEYINPUT114), .B(n691), .Z(n692) );
  NOR2_X1 U746 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U747 ( .A(KEYINPUT53), .B(n694), .ZN(G75) );
  NAND2_X1 U748 ( .A1(n701), .A2(G469), .ZN(n699) );
  XNOR2_X1 U749 ( .A(KEYINPUT58), .B(KEYINPUT115), .ZN(n697) );
  XNOR2_X1 U750 ( .A(n695), .B(KEYINPUT57), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U753 ( .A1(n705), .A2(n700), .ZN(G54) );
  NAND2_X1 U754 ( .A1(n701), .A2(G217), .ZN(n702) );
  XNOR2_X1 U755 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U756 ( .A1(n705), .A2(n704), .ZN(G66) );
  XNOR2_X1 U757 ( .A(n706), .B(KEYINPUT89), .ZN(n708) );
  XNOR2_X1 U758 ( .A(n708), .B(n707), .ZN(n713) );
  XNOR2_X1 U759 ( .A(KEYINPUT123), .B(n713), .ZN(n709) );
  XNOR2_X1 U760 ( .A(G227), .B(n709), .ZN(n710) );
  NAND2_X1 U761 ( .A1(n710), .A2(G900), .ZN(n711) );
  NAND2_X1 U762 ( .A1(n711), .A2(G953), .ZN(n717) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U764 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U765 ( .A1(n717), .A2(n716), .ZN(G72) );
  XNOR2_X1 U766 ( .A(G140), .B(n718), .ZN(G42) );
  XOR2_X1 U767 ( .A(G137), .B(KEYINPUT126), .Z(n719) );
  XNOR2_X1 U768 ( .A(n720), .B(n719), .ZN(G39) );
  XNOR2_X1 U769 ( .A(G122), .B(KEYINPUT124), .ZN(n722) );
  XNOR2_X1 U770 ( .A(n722), .B(n721), .ZN(G24) );
  XNOR2_X1 U771 ( .A(G131), .B(KEYINPUT127), .ZN(n724) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(G33) );
endmodule

