//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT69), .Z(G261));
  AOI22_X1  g031(.A1(new_n451), .A2(G567), .B1(new_n454), .B2(G2106), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT70), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n460), .B1(new_n465), .B2(KEYINPUT71), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n462), .A2(new_n464), .A3(new_n468), .A4(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n459), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G2105), .B1(G101), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n470), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n466), .A2(new_n469), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n479), .A2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(G136), .B2(new_n485), .ZN(G162));
  XOR2_X1   g061(.A(KEYINPUT72), .B(KEYINPUT4), .Z(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR4_X1   g063(.A1(new_n487), .A2(new_n473), .A3(new_n488), .A4(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n465), .A2(KEYINPUT71), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n488), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n490), .A2(new_n469), .A3(new_n459), .A4(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n489), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n493), .A2(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT73), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(new_n510), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n509), .A2(new_n516), .ZN(G166));
  AND2_X1   g092(.A1(new_n506), .A2(new_n510), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G89), .B1(G51), .B2(new_n512), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT75), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n504), .A2(new_n524), .A3(new_n505), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n524), .B1(new_n504), .B2(new_n505), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n523), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n518), .A2(G90), .B1(G52), .B2(new_n512), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n508), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  NAND2_X1  g108(.A1(new_n512), .A2(G43), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n514), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(G68), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n504), .A2(new_n505), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n504), .A2(new_n524), .A3(new_n505), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n536), .B1(new_n543), .B2(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT76), .Z(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n518), .A2(G91), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OR3_X1    g127(.A1(new_n511), .A2(KEYINPUT9), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n511), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n551), .B(new_n555), .C1(new_n508), .C2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G168), .ZN(G286));
  INV_X1    g133(.A(G166), .ZN(G303));
  AOI22_X1  g134(.A1(new_n518), .A2(G87), .B1(G49), .B2(new_n512), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT77), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(new_n564), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G288));
  NAND3_X1  g142(.A1(new_n504), .A2(G61), .A3(new_n505), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n568), .A2(KEYINPUT78), .B1(G73), .B2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n508), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n512), .A2(G48), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n514), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  XNOR2_X1  g151(.A(KEYINPUT80), .B(G85), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n518), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(KEYINPUT79), .B(G47), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n512), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT81), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n578), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n508), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(KEYINPUT82), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT82), .B1(new_n585), .B2(new_n588), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G171), .A2(G868), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n506), .A2(G92), .A3(new_n510), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n538), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(new_n512), .B2(G54), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT83), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n594), .B1(new_n603), .B2(G868), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT84), .ZN(G284));
  XOR2_X1   g180(.A(new_n604), .B(KEYINPUT85), .Z(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(G168), .B2(new_n607), .ZN(G280));
  INV_X1    g185(.A(G860), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n603), .B1(G559), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT86), .Z(G148));
  INV_X1    g188(.A(new_n544), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n607), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n603), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g193(.A1(new_n476), .A2(new_n459), .A3(new_n472), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n485), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n480), .A2(G123), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n625), .A2(KEYINPUT87), .B1(new_n626), .B2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(KEYINPUT87), .B2(new_n625), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT88), .B(G2096), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n622), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT91), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT90), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT14), .ZN(new_n647));
  OAI21_X1  g222(.A(G14), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n641), .ZN(G401));
  XOR2_X1   g224(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n653), .B2(new_n650), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n656), .B(new_n658), .Z(new_n659));
  XNOR2_X1  g234(.A(G2096), .B(G2100), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  AOI211_X1 g246(.A(new_n668), .B(new_n671), .C1(new_n663), .C2(new_n667), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  NAND2_X1  g253(.A1(new_n592), .A2(G16), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G16), .B2(G24), .ZN(new_n680));
  INV_X1    g255(.A(G1986), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(G6), .A2(G16), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n575), .B2(G16), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G23), .ZN(new_n688));
  INV_X1    g263(.A(new_n562), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT33), .B(G1976), .Z(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(G22), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G166), .B2(new_n687), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n686), .A2(new_n692), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT34), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n680), .A2(new_n681), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n485), .A2(G131), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n480), .A2(G119), .ZN(new_n702));
  OR2_X1    g277(.A1(G95), .A2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n703), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT94), .B(G29), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G25), .B(new_n705), .S(new_n707), .Z(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT35), .B(G1991), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR4_X1   g285(.A1(new_n682), .A2(new_n699), .A3(new_n700), .A4(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT36), .Z(new_n712));
  NOR2_X1   g287(.A1(new_n629), .A2(new_n706), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT102), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT103), .B(G2078), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT104), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n707), .A2(G27), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G164), .B2(new_n707), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n714), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n687), .A2(G20), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT23), .ZN(new_n721));
  INV_X1    g296(.A(G299), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n687), .ZN(new_n723));
  INV_X1    g298(.A(G1956), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G11), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT30), .B(G28), .Z(new_n727));
  OAI211_X1 g302(.A(new_n725), .B(new_n726), .C1(G29), .C2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(G34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(G34), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n706), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G160), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n719), .B(new_n728), .C1(new_n729), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n687), .A2(G4), .ZN(new_n738));
  INV_X1    g313(.A(new_n603), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n687), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G1348), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n687), .A2(G19), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n544), .B2(new_n687), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1341), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n740), .B2(G1348), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n718), .A2(new_n716), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n687), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n687), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(new_n749), .B2(G1961), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT98), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G105), .B2(new_n476), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n485), .A2(G141), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n480), .A2(G129), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n735), .A2(G32), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT99), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n750), .B(new_n764), .C1(G1961), .C2(new_n749), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n737), .A2(new_n741), .A3(new_n746), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n706), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n485), .A2(G140), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT96), .Z(new_n770));
  OR2_X1    g345(.A1(new_n467), .A2(G116), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n480), .A2(G128), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(new_n735), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT97), .ZN(new_n778));
  INV_X1    g353(.A(G2067), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n736), .A2(new_n729), .ZN(new_n781));
  INV_X1    g356(.A(G2072), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n735), .A2(G33), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n485), .A2(G139), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT25), .Z(new_n786));
  INV_X1    g361(.A(G127), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n473), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n784), .B(new_n786), .C1(new_n467), .C2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(G29), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n781), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n782), .B2(new_n791), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n763), .B2(new_n760), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT100), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n707), .A2(G35), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G162), .B2(new_n707), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT29), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G2090), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n687), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n687), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT101), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1966), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n766), .A2(new_n780), .A3(new_n795), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n712), .A2(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n739), .A2(G559), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT38), .Z(new_n809));
  NAND3_X1  g384(.A1(new_n539), .A2(G67), .A3(new_n540), .ZN(new_n810));
  INV_X1    g385(.A(G80), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n499), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT105), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n810), .A2(KEYINPUT105), .A3(new_n813), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(new_n817), .A3(G651), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n506), .A2(G93), .A3(new_n510), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n512), .A2(G55), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT106), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n819), .A2(KEYINPUT106), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n818), .A2(new_n825), .A3(new_n544), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n544), .B1(new_n818), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n809), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n830));
  AOI21_X1  g405(.A(G860), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n810), .A2(KEYINPUT105), .A3(new_n813), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT105), .B1(new_n810), .B2(new_n813), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n833), .A2(new_n834), .A3(new_n508), .ZN(new_n835));
  INV_X1    g410(.A(new_n825), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(new_n611), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n832), .A2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n775), .B(G164), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n480), .A2(G130), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n467), .A2(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G142), .B2(new_n485), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n841), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT107), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n705), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n620), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n757), .B(new_n790), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n847), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n629), .B(G160), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  AOI21_X1  g430(.A(G37), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n853), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g433(.A(KEYINPUT82), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n578), .A2(new_n583), .A3(new_n580), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n583), .B1(new_n578), .B2(new_n580), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n859), .B1(new_n862), .B2(new_n587), .ZN(new_n863));
  AOI21_X1  g438(.A(G305), .B1(new_n863), .B2(new_n589), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n562), .B(G166), .Z(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(G305), .A3(new_n589), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n863), .A2(G305), .A3(new_n589), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(new_n864), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT42), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n616), .B(new_n828), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n595), .B(KEYINPUT10), .ZN(new_n875));
  INV_X1    g450(.A(new_n601), .ZN(new_n876));
  OAI21_X1  g451(.A(G299), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n556), .A2(new_n508), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n518), .A2(G91), .B1(new_n553), .B2(new_n554), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n597), .A2(new_n878), .A3(new_n879), .A4(new_n601), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n877), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n874), .A2(new_n884), .ZN(new_n885));
  NOR3_X1   g460(.A1(G299), .A2(new_n875), .A3(new_n876), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n597), .A2(new_n601), .B1(new_n878), .B2(new_n879), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT108), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n885), .B1(new_n874), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n873), .B1(new_n890), .B2(KEYINPUT109), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(KEYINPUT109), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G868), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g470(.A(new_n894), .B1(G868), .B2(new_n837), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n898));
  NAND2_X1  g473(.A1(G301), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n826), .B2(new_n827), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n614), .B1(new_n835), .B2(new_n836), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n818), .A2(new_n825), .A3(new_n544), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n903), .A3(new_n899), .ZN(new_n904));
  AOI21_X1  g479(.A(G286), .B1(G171), .B2(KEYINPUT111), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n901), .B2(new_n904), .ZN(new_n907));
  OAI22_X1  g482(.A1(new_n906), .A2(new_n907), .B1(new_n882), .B2(new_n883), .ZN(new_n908));
  INV_X1    g483(.A(new_n905), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n826), .A2(new_n827), .A3(new_n900), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n888), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n872), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n872), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n889), .A3(new_n913), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT41), .B1(new_n886), .B2(new_n887), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(KEYINPUT113), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT113), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n883), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(new_n912), .B2(new_n913), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n919), .B1(new_n926), .B2(KEYINPUT114), .ZN(new_n927));
  AOI211_X1 g502(.A(KEYINPUT113), .B(new_n881), .C1(new_n877), .C2(new_n880), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n884), .B2(KEYINPUT113), .ZN(new_n929));
  OAI211_X1 g504(.A(KEYINPUT114), .B(new_n929), .C1(new_n906), .C2(new_n907), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(KEYINPUT115), .B(new_n918), .C1(new_n927), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(new_n906), .B2(new_n907), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT114), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n930), .A3(new_n919), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT115), .B1(new_n937), .B2(new_n918), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n917), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n908), .A2(new_n914), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n941), .B(new_n916), .C1(new_n942), .C2(new_n872), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n872), .B1(new_n908), .B2(new_n914), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT112), .B1(new_n944), .B2(G37), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n943), .A2(new_n945), .A3(new_n915), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n897), .B1(new_n940), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n917), .B(new_n946), .C1(new_n933), .C2(new_n938), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n945), .A3(new_n915), .ZN(new_n950));
  INV_X1    g525(.A(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n949), .A2(new_n952), .A3(new_n897), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n948), .A2(new_n953), .ZN(G397));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n493), .B2(new_n497), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(KEYINPUT45), .B(new_n955), .C1(new_n493), .C2(new_n497), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n470), .A2(new_n477), .A3(G40), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT56), .B(G2072), .Z(new_n964));
  NOR3_X1   g539(.A1(new_n959), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n494), .A2(new_n496), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n967));
  INV_X1    g542(.A(new_n489), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n955), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT122), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n956), .A2(KEYINPUT50), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n962), .ZN(new_n975));
  AOI211_X1 g550(.A(KEYINPUT122), .B(new_n961), .C1(new_n956), .C2(KEYINPUT50), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n965), .B1(new_n977), .B2(new_n724), .ZN(new_n978));
  XNOR2_X1  g553(.A(G299), .B(KEYINPUT57), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT125), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT125), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n971), .B1(new_n970), .B2(new_n955), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT122), .B1(new_n983), .B2(new_n961), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n961), .B1(new_n956), .B2(KEYINPUT50), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n973), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G1956), .B1(new_n987), .B2(new_n972), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n982), .B(new_n979), .C1(new_n988), .C2(new_n965), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT61), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n978), .B2(new_n980), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n981), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n978), .A2(new_n980), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n979), .B(new_n965), .C1(new_n977), .C2(new_n724), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT60), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n985), .A2(new_n972), .ZN(new_n997));
  INV_X1    g572(.A(G1348), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n956), .A2(new_n961), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n999), .B(new_n602), .C1(G2067), .C2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(G2067), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1348), .B1(new_n985), .B2(new_n972), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n597), .B(new_n601), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n996), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT59), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n958), .A2(new_n1008), .A3(new_n962), .A4(new_n960), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT58), .B(G1341), .Z(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n956), .B2(new_n961), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1007), .B1(new_n1012), .B2(new_n544), .ZN(new_n1013));
  AOI211_X1 g588(.A(KEYINPUT59), .B(new_n614), .C1(new_n1009), .C2(new_n1011), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR4_X1   g590(.A1(new_n1003), .A2(new_n1004), .A3(KEYINPUT60), .A4(new_n602), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1006), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n992), .A2(new_n995), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n989), .A2(new_n981), .A3(new_n1005), .ZN(new_n1019));
  INV_X1    g594(.A(new_n994), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT126), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(KEYINPUT126), .A3(new_n1021), .ZN(new_n1025));
  INV_X1    g600(.A(G2078), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n958), .A2(new_n1026), .A3(new_n962), .A4(new_n960), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  INV_X1    g605(.A(G1961), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n997), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G171), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1032), .A2(new_n1030), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT45), .B1(new_n956), .B2(KEYINPUT116), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(KEYINPUT116), .B2(new_n956), .ZN(new_n1037));
  INV_X1    g612(.A(new_n963), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(KEYINPUT53), .A3(new_n1026), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(G301), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n959), .B2(new_n963), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n985), .A2(new_n729), .A3(new_n972), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1045), .A2(G286), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G286), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT51), .B(G8), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1045), .A2(G168), .A3(new_n1046), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1039), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G171), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(KEYINPUT54), .C1(G171), .C2(new_n1033), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1043), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT118), .B(G2090), .Z(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n972), .C1(new_n975), .C2(new_n976), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1971), .B1(new_n1038), .B2(new_n958), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1052), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT55), .B(G8), .C1(new_n509), .C2(new_n516), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT119), .ZN(new_n1066));
  OAI21_X1  g641(.A(G8), .B1(new_n509), .B2(new_n516), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OR3_X1    g647(.A1(new_n1063), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n985), .A2(new_n1059), .A3(new_n972), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1072), .B(G8), .C1(new_n1061), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n1076));
  INV_X1    g651(.A(G1976), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n563), .A2(new_n1077), .A3(new_n565), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n560), .A2(G1976), .A3(new_n561), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(G8), .C1(new_n956), .C2(new_n961), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1076), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1082), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(KEYINPUT121), .A3(new_n1079), .A4(new_n1078), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1981), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n575), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(G1981), .B1(new_n571), .B2(new_n574), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1088), .A2(KEYINPUT49), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT49), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1000), .A2(new_n1052), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1092), .A2(new_n1093), .B1(KEYINPUT52), .B2(new_n1082), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1075), .A2(new_n1086), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1064), .B1(new_n1063), .B2(new_n1072), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1073), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT127), .B1(new_n1058), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT54), .B1(new_n1033), .B2(G171), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1049), .B(new_n1053), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT54), .B1(new_n1034), .B2(new_n1040), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1073), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT127), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1024), .A2(new_n1025), .A3(new_n1098), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(new_n1075), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1077), .B(new_n566), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1052), .B(new_n1000), .C1(new_n1110), .C2(new_n1088), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1048), .A2(G8), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1073), .A2(new_n1095), .A3(new_n1096), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1075), .A2(new_n1086), .A3(new_n1094), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1113), .A2(KEYINPUT63), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1061), .A2(new_n1074), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1072), .B1(new_n1119), .B2(G8), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT124), .B(new_n1112), .C1(new_n1116), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1112), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1034), .B1(new_n1054), .B2(KEYINPUT62), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1104), .B(new_n1127), .C1(KEYINPUT62), .C2(new_n1054), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1107), .A2(new_n1122), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1037), .A2(new_n961), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1008), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n757), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1130), .B(KEYINPUT117), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n776), .A2(new_n779), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n775), .A2(G2067), .ZN(new_n1135));
  INV_X1    g710(.A(new_n757), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1134), .B(new_n1135), .C1(new_n1008), .C2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n705), .A2(new_n709), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n705), .A2(new_n709), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1133), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n592), .B(new_n681), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1130), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1129), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1133), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n1147), .B2(new_n1134), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1131), .B(KEYINPUT46), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1134), .A2(new_n1136), .A3(new_n1135), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT47), .Z(new_n1152));
  INV_X1    g727(.A(new_n1142), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n592), .A2(new_n681), .A3(new_n1130), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT48), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1148), .B(new_n1152), .C1(new_n1153), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1145), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g732(.A1(new_n949), .A2(new_n952), .ZN(new_n1159));
  INV_X1    g733(.A(G227), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1160), .A2(G319), .ZN(new_n1161));
  NOR3_X1   g735(.A1(G229), .A2(G401), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n857), .A3(new_n1162), .ZN(G225));
  INV_X1    g737(.A(G225), .ZN(G308));
endmodule


