//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT75), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n204), .B(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NOR4_X1   g013(.A1(KEYINPUT66), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n216), .B1(new_n214), .B2(new_n213), .ZN(new_n217));
  OAI221_X1 g016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT27), .B(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n221), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n223), .A3(new_n220), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n227), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n229), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n231), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n230), .A3(new_n212), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT64), .ZN(new_n241));
  INV_X1    g040(.A(new_n236), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT25), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n225), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(G226gat), .A2(G233gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(KEYINPUT29), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n237), .B1(new_n231), .B2(new_n236), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n241), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(new_n225), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n211), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G8gat), .B(G36gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT76), .ZN(new_n255));
  XNOR2_X1  g054(.A(G64gat), .B(G92gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  NOR3_X1   g056(.A1(new_n246), .A2(new_n251), .A3(new_n211), .ZN(new_n258));
  OR3_X1    g057(.A1(new_n253), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n258), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n252), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n257), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n262), .A3(KEYINPUT30), .ZN(new_n263));
  OR3_X1    g062(.A1(new_n261), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n267));
  INV_X1    g066(.A(G141gat), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(G148gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT81), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G155gat), .ZN(new_n273));
  INV_X1    g072(.A(G162gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT81), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT80), .B(G148gat), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n278), .B(new_n270), .C1(new_n279), .C2(new_n268), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT82), .B(G155gat), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT2), .B1(new_n281), .B2(new_n274), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n272), .A2(new_n277), .A3(new_n280), .A4(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT78), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n276), .A2(new_n284), .A3(KEYINPUT2), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G141gat), .B(G148gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n284), .B1(new_n276), .B2(KEYINPUT2), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT79), .ZN(new_n290));
  AND2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT77), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n294), .A3(new_n276), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n289), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n293), .A2(new_n295), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT78), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G141gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n270), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n285), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT79), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n283), .B1(new_n297), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n290), .B1(new_n289), .B2(new_n296), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n298), .A2(KEYINPUT79), .A3(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(new_n283), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n314));
  INV_X1    g113(.A(G113gat), .ZN(new_n315));
  INV_X1    g114(.A(G120gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318));
  NAND2_X1  g117(.A1(G113gat), .A2(G120gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G134gat), .ZN(new_n321));
  OR3_X1    g120(.A1(new_n321), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n314), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n324));
  NAND4_X1  g123(.A1(new_n324), .A2(new_n313), .A3(new_n317), .A4(new_n319), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n312), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(new_n306), .B2(new_n326), .ZN(new_n330));
  INV_X1    g129(.A(new_n326), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n310), .A2(KEYINPUT4), .A3(new_n283), .A4(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n327), .A2(new_n328), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT83), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n330), .A2(new_n332), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n339), .A2(new_n328), .A3(new_n327), .A4(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n306), .B(new_n331), .ZN(new_n342));
  INV_X1    g141(.A(new_n328), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT0), .ZN(new_n349));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n345), .B1(new_n338), .B2(new_n340), .ZN(new_n354));
  INV_X1    g153(.A(new_n351), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(KEYINPUT6), .A3(new_n355), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n265), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G22gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n211), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n312), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n306), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n203), .A2(KEYINPUT87), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(new_n210), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(KEYINPUT87), .B2(new_n203), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n367), .B2(new_n210), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT3), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n365), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n311), .B1(new_n211), .B2(KEYINPUT29), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n363), .B1(new_n306), .B2(new_n373), .ZN(new_n374));
  OAI221_X1 g173(.A(new_n360), .B1(new_n363), .B2(new_n372), .C1(new_n374), .C2(new_n365), .ZN(new_n375));
  INV_X1    g174(.A(new_n363), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n306), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n365), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n372), .A2(new_n363), .ZN(new_n379));
  OAI21_X1  g178(.A(G22gat), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT86), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n375), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n375), .A2(new_n380), .A3(KEYINPUT88), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(G50gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n382), .A2(new_n383), .A3(new_n389), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n244), .A2(new_n331), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n250), .A2(new_n326), .A3(new_n225), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G227gat), .ZN(new_n397));
  INV_X1    g196(.A(G233gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT34), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n399), .B2(new_n402), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n397), .A2(new_n398), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n394), .A2(new_n406), .A3(new_n395), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n407), .A2(KEYINPUT32), .ZN(new_n408));
  XNOR2_X1  g207(.A(G15gat), .B(G43gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n411), .A2(KEYINPUT72), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(KEYINPUT72), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n414));
  OR3_X1    g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n411), .B1(new_n407), .B2(KEYINPUT32), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT70), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n407), .A2(new_n419), .A3(new_n414), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n407), .B2(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT71), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n420), .A4(new_n418), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n417), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n405), .B1(new_n427), .B2(KEYINPUT74), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT74), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n429), .B(new_n417), .C1(new_n423), .C2(new_n426), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n423), .A2(new_n426), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n416), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n433), .A2(new_n405), .A3(new_n429), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n359), .B(new_n393), .C1(new_n431), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT35), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(KEYINPUT91), .A3(KEYINPUT35), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n431), .B2(new_n434), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n433), .A2(new_n429), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT74), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n405), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n430), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT90), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT35), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n359), .A2(new_n393), .A3(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n438), .A2(new_n439), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n339), .A2(new_n327), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n343), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT39), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n342), .B2(new_n328), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n454), .A3(new_n343), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n351), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n456), .A2(KEYINPUT40), .A3(new_n351), .A4(new_n457), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n263), .A2(new_n264), .ZN(new_n463));
  AOI211_X1 g262(.A(new_n351), .B(new_n345), .C1(new_n338), .C2(new_n340), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n462), .A2(new_n465), .B1(new_n391), .B2(new_n392), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(new_n464), .ZN(new_n468));
  INV_X1    g267(.A(new_n358), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT37), .B1(new_n253), .B2(new_n258), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n260), .A2(new_n252), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT38), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n471), .A2(new_n473), .A3(new_n474), .A4(new_n257), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n475), .A2(new_n259), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT89), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n357), .A2(KEYINPUT89), .A3(new_n358), .A4(new_n476), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n471), .A2(new_n473), .A3(new_n257), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT38), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n466), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n444), .A2(KEYINPUT36), .A3(new_n445), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n431), .B2(new_n434), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n359), .A2(new_n393), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n482), .A2(new_n483), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n202), .B1(new_n451), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n450), .A2(new_n441), .A3(new_n446), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n435), .A2(KEYINPUT91), .A3(KEYINPUT35), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT91), .B1(new_n435), .B2(KEYINPUT35), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT92), .A3(new_n487), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497));
  OR2_X1    g296(.A1(G43gat), .A2(G50gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(G43gat), .A2(G50gat), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(G29gat), .A2(G36gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT14), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT93), .B(G50gat), .Z(new_n506));
  OAI211_X1 g305(.A(new_n497), .B(new_n499), .C1(new_n506), .C2(G43gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(KEYINPUT94), .B2(new_n502), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n502), .A2(KEYINPUT94), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n503), .B(KEYINPUT95), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(new_n500), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n505), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT17), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(G1gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(G1gat), .B2(new_n515), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G8gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n513), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT18), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT96), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n519), .B(new_n513), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n522), .B(KEYINPUT13), .Z(new_n528));
  AOI22_X1  g327(.A1(new_n524), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(KEYINPUT96), .A3(new_n525), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G197gat), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT11), .B(G169gat), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT12), .Z(new_n537));
  OAI21_X1  g336(.A(new_n496), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n529), .A2(KEYINPUT97), .A3(new_n539), .A4(new_n531), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n538), .A2(new_n540), .B1(new_n537), .B2(new_n532), .ZN(new_n541));
  XNOR2_X1  g340(.A(G57gat), .B(G64gat), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT98), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G71gat), .B(G78gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G85gat), .A2(G92gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT101), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT101), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n548), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G99gat), .B(G106gat), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT102), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(G85gat), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT8), .A2(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n550), .A2(new_n554), .A3(new_n556), .A4(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n555), .A2(KEYINPUT102), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n561), .A2(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n547), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n562), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n546), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT103), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT105), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n567), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT103), .A3(new_n547), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n574), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT104), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n565), .A2(new_n577), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT10), .B1(new_n570), .B2(new_n574), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT104), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n572), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT106), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI211_X1 g385(.A(KEYINPUT106), .B(new_n572), .C1(new_n579), .C2(new_n583), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n575), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(G176gat), .B(G204gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n579), .A2(new_n583), .ZN(new_n594));
  INV_X1    g393(.A(new_n572), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n575), .A3(new_n591), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n546), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G127gat), .ZN(new_n604));
  XOR2_X1   g403(.A(G183gat), .B(G211gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n520), .B1(new_n600), .B2(new_n546), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT99), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n273), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n606), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n514), .A2(new_n567), .A3(new_n566), .ZN(new_n616));
  AND2_X1   g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n573), .A2(new_n513), .B1(KEYINPUT41), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n622));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n621), .B(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n599), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n495), .A2(new_n541), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n470), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  INV_X1    g429(.A(new_n628), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n463), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT16), .B(G8gat), .Z(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G8gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT42), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n633), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(G1325gat));
  AND2_X1   g440(.A1(new_n485), .A2(new_n483), .ZN(new_n642));
  OAI21_X1  g441(.A(G15gat), .B1(new_n631), .B2(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n447), .A2(G15gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n631), .B2(new_n644), .ZN(G1326gat));
  INV_X1    g444(.A(new_n393), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT43), .B(G22gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  AND3_X1   g448(.A1(new_n493), .A2(KEYINPUT92), .A3(new_n487), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT92), .B1(new_n493), .B2(new_n487), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n541), .ZN(new_n653));
  INV_X1    g452(.A(new_n625), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n598), .A2(new_n614), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n470), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n656), .A2(G29gat), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT45), .Z(new_n659));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n487), .A2(KEYINPUT108), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n642), .A2(new_n663), .A3(new_n486), .A4(new_n482), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n493), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n625), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n652), .A2(new_n661), .B1(new_n660), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n598), .B(KEYINPUT107), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n669), .A2(new_n541), .A3(new_n614), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G29gat), .B1(new_n671), .B2(new_n657), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n659), .A2(new_n672), .ZN(G1328gat));
  NOR3_X1   g472(.A1(new_n656), .A2(G36gat), .A3(new_n463), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT46), .ZN(new_n675));
  OAI21_X1  g474(.A(G36gat), .B1(new_n671), .B2(new_n463), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1329gat));
  NOR2_X1   g476(.A1(new_n495), .A2(new_n541), .ZN(new_n678));
  INV_X1    g477(.A(G43gat), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n678), .A2(new_n679), .A3(new_n448), .A4(new_n655), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n671), .A2(new_n642), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(KEYINPUT47), .B(new_n680), .C1(new_n681), .C2(new_n679), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1330gat));
  INV_X1    g485(.A(new_n506), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n660), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n489), .A2(new_n494), .A3(new_n661), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n688), .A2(new_n646), .A3(new_n689), .A4(new_n670), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n667), .A2(KEYINPUT110), .A3(new_n646), .A4(new_n670), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n646), .A2(new_n687), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT109), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT48), .B1(new_n656), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n690), .A2(new_n506), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n678), .A2(new_n655), .A3(new_n696), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT48), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(KEYINPUT111), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n698), .B1(new_n692), .B2(new_n693), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n703), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(G1331gat));
  NOR4_X1   g508(.A1(new_n668), .A2(new_n653), .A3(new_n615), .A4(new_n625), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n665), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n657), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT112), .B(G57gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1332gat));
  NOR2_X1   g513(.A1(new_n711), .A2(new_n463), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  AND2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n715), .B2(new_n716), .ZN(G1333gat));
  OAI21_X1  g518(.A(G71gat), .B1(new_n711), .B2(new_n642), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n447), .A2(G71gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n711), .B2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g522(.A1(new_n711), .A2(new_n393), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g524(.A1(new_n653), .A2(new_n614), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(new_n598), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n667), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G85gat), .B1(new_n728), .B2(new_n657), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  INV_X1    g529(.A(new_n726), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n666), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n665), .A2(KEYINPUT51), .A3(new_n625), .A4(new_n726), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n599), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n558), .A3(new_n470), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n735), .ZN(G1336gat));
  OAI21_X1  g535(.A(G92gat), .B1(new_n728), .B2(new_n463), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n668), .B1(new_n732), .B2(new_n733), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n265), .A2(new_n559), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT52), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n737), .B(new_n743), .C1(new_n739), .C2(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n728), .B2(new_n642), .ZN(new_n746));
  INV_X1    g545(.A(G99gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n734), .A2(new_n747), .A3(new_n448), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1338gat));
  NAND4_X1  g548(.A1(new_n688), .A2(new_n646), .A3(new_n689), .A4(new_n727), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G106gat), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT53), .B1(new_n751), .B2(KEYINPUT113), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n393), .A2(G106gat), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n738), .A2(new_n753), .B1(new_n750), .B2(G106gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n752), .B(new_n754), .ZN(G1339gat));
  NAND2_X1  g554(.A1(new_n596), .A2(KEYINPUT106), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n584), .A2(new_n585), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n594), .B2(new_n595), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n579), .A2(new_n583), .A3(new_n572), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n591), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT55), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n765), .A2(new_n653), .A3(new_n597), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n538), .A2(new_n540), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n527), .A2(new_n528), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n536), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT115), .Z(new_n772));
  AND2_X1   g571(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n598), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n625), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n766), .A2(new_n597), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n768), .A2(new_n625), .A3(new_n772), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n765), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n615), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n627), .B2(new_n653), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n599), .A2(new_n626), .A3(KEYINPUT114), .A4(new_n541), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n657), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n431), .A2(new_n434), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n646), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(new_n463), .ZN(new_n789));
  AOI21_X1  g588(.A(G113gat), .B1(new_n789), .B2(new_n653), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n780), .A2(new_n784), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n393), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT116), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n794), .A3(new_n393), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n657), .A2(new_n265), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n448), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n541), .A2(new_n315), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n790), .B1(new_n799), .B2(new_n800), .ZN(G1340gat));
  AOI21_X1  g600(.A(G120gat), .B1(new_n789), .B2(new_n598), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n668), .A2(new_n316), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n799), .B2(new_n803), .ZN(G1341gat));
  INV_X1    g603(.A(G127gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n805), .A3(new_n614), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n796), .A2(new_n615), .A3(new_n798), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n805), .ZN(G1342gat));
  NAND2_X1  g607(.A1(new_n625), .A2(new_n463), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n809), .B(KEYINPUT117), .Z(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n788), .A2(new_n321), .A3(new_n811), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT56), .Z(new_n813));
  NOR3_X1   g612(.A1(new_n796), .A2(new_n654), .A3(new_n798), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n321), .B2(new_n814), .ZN(G1343gat));
  NAND2_X1  g614(.A1(new_n642), .A2(new_n797), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n393), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n767), .A2(new_n774), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n541), .B1(new_n763), .B2(new_n764), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n776), .A2(new_n822), .B1(new_n598), .B2(new_n773), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT118), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n824), .A3(new_n654), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n614), .B1(new_n825), .B2(new_n778), .ZN(new_n826));
  INV_X1    g625(.A(new_n784), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n818), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n791), .A2(new_n646), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n817), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n816), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n541), .A2(new_n268), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n642), .A2(new_n646), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT119), .Z(new_n834));
  NAND4_X1  g633(.A1(new_n785), .A2(new_n834), .A3(new_n463), .A4(new_n653), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n831), .A2(new_n832), .B1(new_n268), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT120), .B(KEYINPUT58), .C1(new_n836), .C2(KEYINPUT121), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838));
  INV_X1    g637(.A(new_n816), .ZN(new_n839));
  INV_X1    g638(.A(new_n818), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n654), .B1(new_n823), .B2(KEYINPUT118), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n819), .A2(new_n820), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n778), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n615), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n840), .B1(new_n844), .B2(new_n784), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT57), .B1(new_n791), .B2(new_n646), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n839), .B(new_n832), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n835), .A2(new_n268), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n838), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n849), .B2(new_n838), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n837), .B1(new_n851), .B2(new_n853), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n627), .A2(new_n653), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n817), .B(new_n646), .C1(new_n826), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n829), .A2(KEYINPUT57), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n598), .A3(new_n839), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n831), .A2(new_n861), .A3(new_n598), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n785), .A2(new_n834), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(new_n463), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n864), .B2(new_n598), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n860), .B(new_n862), .C1(new_n279), .C2(new_n865), .ZN(G1345gat));
  AND3_X1   g665(.A1(new_n863), .A2(new_n463), .A3(new_n614), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n615), .A2(new_n281), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n869), .A2(new_n281), .B1(new_n831), .B2(new_n870), .ZN(G1346gat));
  NAND3_X1  g670(.A1(new_n863), .A2(new_n274), .A3(new_n811), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n831), .A2(new_n625), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n274), .ZN(G1347gat));
  AOI21_X1  g673(.A(new_n470), .B1(new_n780), .B2(new_n784), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n265), .A3(new_n787), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n653), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n470), .A2(new_n463), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n448), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n793), .B2(new_n795), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n653), .A2(G169gat), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(G1348gat));
  INV_X1    g682(.A(G176gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n877), .A2(new_n884), .A3(new_n598), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n881), .A2(new_n669), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n884), .ZN(G1349gat));
  INV_X1    g686(.A(G183gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n881), .B2(new_n614), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n877), .A2(new_n219), .A3(new_n614), .ZN(new_n890));
  XNOR2_X1  g689(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n889), .B2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1350gat));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n220), .A3(new_n625), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n625), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(KEYINPUT61), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n220), .B1(new_n898), .B2(KEYINPUT61), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n897), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(G1351gat));
  AND2_X1   g702(.A1(new_n642), .A2(new_n879), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n858), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(G197gat), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(new_n541), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n875), .A2(new_n642), .A3(new_n265), .A4(new_n646), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT125), .Z(new_n909));
  AOI21_X1  g708(.A(G197gat), .B1(new_n909), .B2(new_n653), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n907), .A2(new_n910), .ZN(G1352gat));
  XNOR2_X1  g710(.A(KEYINPUT126), .B(G204gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n908), .A2(new_n599), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT62), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n856), .A2(new_n669), .A3(new_n857), .A4(new_n904), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n912), .B1(new_n915), .B2(KEYINPUT127), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1353gat));
  NAND3_X1  g717(.A1(new_n909), .A2(new_n207), .A3(new_n614), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n856), .A2(new_n614), .A3(new_n857), .A4(new_n904), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n920), .B2(G211gat), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n920), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(G1354gat));
  OAI21_X1  g722(.A(G218gat), .B1(new_n905), .B2(new_n654), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n208), .A3(new_n625), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1355gat));
endmodule


