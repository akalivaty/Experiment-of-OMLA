//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n438, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G96), .ZN(new_n438));
  INV_X1    g013(.A(new_n438), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G132), .A4(new_n438), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(new_n461));
  INV_X1    g036(.A(G2106), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(new_n455), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n466), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n475), .A2(G137), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(G101), .A3(G2104), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n473), .A2(new_n479), .A3(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n478), .A2(new_n474), .A3(G2105), .A4(new_n469), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT71), .ZN(new_n490));
  AND4_X1   g065(.A1(new_n476), .A2(new_n478), .A3(new_n474), .A4(new_n469), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(G136), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n478), .A2(new_n474), .A3(new_n496), .A4(new_n469), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n467), .A2(new_n469), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(G114), .B2(new_n476), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n482), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n500), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT72), .B1(new_n508), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(new_n518), .A3(new_n514), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n507), .A2(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n522), .B1(new_n528), .B2(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(new_n522), .A3(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n521), .B1(new_n530), .B2(new_n531), .ZN(G166));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n533), .B1(new_n524), .B2(new_n525), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n536), .B(new_n533), .C1(new_n524), .C2(new_n525), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n513), .A2(G51), .A3(G543), .A4(new_n514), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n538), .A2(KEYINPUT75), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT75), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n513), .A2(G89), .A3(new_n518), .A4(new_n514), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n543), .B1(new_n542), .B2(new_n545), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n540), .A2(new_n541), .B1(new_n546), .B2(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n516), .B2(new_n517), .ZN(new_n553));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT77), .B(new_n554), .C1(new_n526), .C2(new_n552), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n556), .A2(G651), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n513), .A2(G52), .A3(G543), .A4(new_n514), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n513), .A2(G90), .A3(new_n518), .A4(new_n514), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n550), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n556), .A2(G651), .A3(new_n557), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G171));
  NAND2_X1  g141(.A1(G68), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G56), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n526), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n509), .A2(new_n512), .B1(new_n508), .B2(G651), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(G81), .A3(new_n518), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(G43), .A3(G543), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  NAND4_X1  g151(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  NAND4_X1  g155(.A1(new_n513), .A2(G91), .A3(new_n518), .A4(new_n514), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT79), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n571), .A2(new_n583), .A3(G91), .A4(new_n518), .ZN(new_n584));
  NAND2_X1  g159(.A1(G78), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G65), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n526), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n582), .A2(new_n584), .B1(G651), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G53), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT9), .B1(new_n515), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT9), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n571), .A2(new_n591), .A3(G53), .A4(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n588), .A2(new_n593), .ZN(G299));
  INV_X1    g169(.A(G171), .ZN(G301));
  INV_X1    g170(.A(G166), .ZN(G303));
  NAND3_X1  g171(.A1(new_n571), .A2(G49), .A3(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n571), .A2(G87), .A3(new_n518), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G288));
  NAND4_X1  g175(.A1(new_n513), .A2(G48), .A3(G543), .A4(new_n514), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n571), .A2(new_n603), .A3(G48), .A4(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT80), .B1(new_n526), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n518), .A2(new_n608), .A3(G61), .ZN(new_n609));
  NAND2_X1  g184(.A1(G73), .A2(G543), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G651), .ZN(new_n612));
  AND3_X1   g187(.A1(new_n513), .A2(new_n518), .A3(new_n514), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G86), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n605), .A2(new_n612), .A3(new_n614), .ZN(G305));
  INV_X1    g190(.A(new_n515), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G47), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT82), .B(G85), .Z(new_n619));
  OAI221_X1 g194(.A(new_n617), .B1(new_n511), .B2(new_n618), .C1(new_n519), .C2(new_n619), .ZN(G290));
  XNOR2_X1  g195(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n613), .A2(G92), .A3(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n621), .B1(new_n519), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G66), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(new_n516), .B2(new_n517), .ZN(new_n627));
  AND2_X1   g202(.A1(G79), .A2(G543), .ZN(new_n628));
  OAI21_X1  g203(.A(G651), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n571), .A2(G54), .A3(G543), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n623), .A2(new_n625), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(G171), .B2(G868), .ZN(G284));
  XOR2_X1   g208(.A(G284), .B(KEYINPUT84), .Z(G321));
  MUX2_X1   g209(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g210(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g211(.A(new_n631), .ZN(new_n637));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G860), .ZN(G148));
  OAI21_X1  g214(.A(KEYINPUT85), .B1(new_n575), .B2(G868), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G868), .ZN(new_n642));
  MUX2_X1   g217(.A(KEYINPUT85), .B(new_n640), .S(new_n642), .Z(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g219(.A(G123), .ZN(new_n645));
  OR3_X1    g220(.A1(new_n485), .A2(KEYINPUT87), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(KEYINPUT87), .B1(new_n485), .B2(new_n645), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  INV_X1    g223(.A(G111), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(G2105), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n491), .B2(G135), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(G2096), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(G2096), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  NAND2_X1  g232(.A1(KEYINPUT86), .A2(G2100), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(KEYINPUT86), .B2(G2100), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n659), .B1(new_n661), .B2(new_n658), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n653), .A2(new_n654), .A3(new_n662), .ZN(G156));
  XOR2_X1   g238(.A(KEYINPUT15), .B(G2435), .Z(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT89), .B(G2438), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2427), .B(G2430), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n669), .A3(new_n667), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(KEYINPUT14), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT90), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1341), .B(G1348), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2443), .B(G2446), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n676), .B(new_n679), .Z(new_n680));
  XNOR2_X1  g255(.A(G2451), .B(G2454), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT91), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G14), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n676), .B(new_n679), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n682), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(G401));
  XNOR2_X1  g263(.A(G2084), .B(G2090), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT92), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2067), .B(G2678), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(KEYINPUT17), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  AOI21_X1  g270(.A(KEYINPUT18), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2100), .ZN(new_n697));
  NOR2_X1   g272(.A1(G2072), .A2(G2078), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n444), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n693), .B2(KEYINPUT18), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(G2096), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n697), .B(new_n701), .ZN(G227));
  XNOR2_X1  g277(.A(G1971), .B(G1976), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT19), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G1956), .B(G2474), .Z(new_n706));
  XOR2_X1   g281(.A(G1961), .B(G1966), .Z(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT20), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n707), .ZN(new_n711));
  NOR3_X1   g286(.A1(new_n705), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n705), .B2(new_n711), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(G1991), .B(G1996), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n715), .ZN(new_n719));
  INV_X1    g294(.A(new_n717), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n714), .A2(new_n715), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(G1981), .B(G1986), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n718), .B2(new_n722), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(G229));
  NAND3_X1  g301(.A1(new_n483), .A2(G119), .A3(new_n484), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G107), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n491), .B2(G131), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n727), .A2(KEYINPUT93), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G25), .B(new_n736), .S(G29), .Z(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT97), .ZN(new_n742));
  OR2_X1    g317(.A1(G16), .A2(G24), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(G290), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G1986), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n746), .B2(new_n745), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n739), .B1(new_n738), .B2(new_n740), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(G6), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G305), .B2(new_n744), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT32), .B(G1981), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT95), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n744), .A2(G22), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G166), .B2(new_n744), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1971), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n744), .A2(G23), .ZN(new_n761));
  INV_X1    g336(.A(G288), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n744), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT33), .B(G1976), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT96), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n763), .B(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n756), .A2(new_n757), .A3(new_n760), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(KEYINPUT34), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(KEYINPUT34), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n751), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n486), .A2(G129), .ZN(new_n773));
  INV_X1    g348(.A(G105), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n774), .A2(new_n468), .A3(G2105), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT26), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n775), .B(new_n777), .C1(new_n491), .C2(G141), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT100), .ZN(new_n780));
  INV_X1    g355(.A(G29), .ZN(new_n781));
  OR3_X1    g356(.A1(new_n780), .A2(KEYINPUT101), .A3(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(G29), .A2(G32), .ZN(new_n783));
  OAI211_X1 g358(.A(KEYINPUT101), .B(new_n783), .C1(new_n780), .C2(new_n781), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT102), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n785), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n781), .A2(G35), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n781), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT29), .B(G2090), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n744), .A2(G5), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G171), .B2(new_n744), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(G1961), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G34), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT24), .ZN(new_n798));
  AOI21_X1  g373(.A(G29), .B1(new_n797), .B2(KEYINPUT24), .ZN(new_n799));
  AOI22_X1  g374(.A1(G160), .A2(G29), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G2084), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G19), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n575), .B2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n801), .B1(G1341), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G27), .A2(G29), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G164), .B2(G29), .ZN(new_n806));
  INV_X1    g381(.A(G2078), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n803), .A2(G1341), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G2067), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n781), .A2(G26), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT28), .Z(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(G116), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G2105), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n491), .B2(G140), .ZN(new_n817));
  INV_X1    g392(.A(G128), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n485), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(G29), .ZN(new_n820));
  AOI211_X1 g395(.A(new_n804), .B(new_n810), .C1(new_n811), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n744), .A2(G20), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT23), .Z(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G299), .B2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1956), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n781), .A2(G33), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n491), .A2(G139), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT25), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n498), .A2(G127), .ZN(new_n831));
  INV_X1    g406(.A(G115), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n468), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n476), .B1(new_n833), .B2(KEYINPUT99), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n826), .B1(new_n836), .B2(new_n781), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G2072), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n800), .A2(G2084), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT105), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n820), .A2(new_n811), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n796), .A2(new_n821), .A3(new_n825), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n744), .A2(G4), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n637), .B2(new_n744), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1348), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n794), .B2(G1961), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT30), .B(G28), .ZN(new_n848));
  OR2_X1    g423(.A1(KEYINPUT31), .A2(G11), .ZN(new_n849));
  NAND2_X1  g424(.A1(KEYINPUT31), .A2(G11), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n848), .A2(new_n781), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n652), .B2(new_n781), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT104), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n744), .A2(G21), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(G168), .B2(new_n744), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT103), .B(G1966), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n847), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n788), .A2(new_n843), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n771), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n751), .A2(new_n769), .A3(new_n860), .A4(new_n768), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n772), .A2(new_n859), .A3(new_n861), .ZN(G150));
  INV_X1    g437(.A(G150), .ZN(G311));
  XNOR2_X1  g438(.A(KEYINPUT106), .B(G55), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n616), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n511), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n613), .A2(G93), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n574), .A2(KEYINPUT107), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n570), .A2(new_n572), .A3(new_n573), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n637), .A2(G559), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n881));
  AOI21_X1  g456(.A(G860), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n869), .A2(G860), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT37), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G145));
  XNOR2_X1  g461(.A(new_n652), .B(new_n493), .ZN(new_n887));
  XNOR2_X1  g462(.A(G160), .B(KEYINPUT108), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n887), .B(new_n888), .Z(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n819), .B(G164), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n736), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n734), .A2(KEYINPUT109), .A3(new_n735), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n491), .A2(G142), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n476), .A2(G118), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  INV_X1    g474(.A(G130), .ZN(new_n900));
  OAI221_X1 g475(.A(new_n897), .B1(new_n898), .B2(new_n899), .C1(new_n485), .C2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n656), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n891), .A3(new_n894), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n896), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n902), .ZN(new_n905));
  INV_X1    g480(.A(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n895), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n779), .A2(new_n836), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n780), .B2(new_n836), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n904), .B2(new_n907), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n890), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n904), .A2(new_n907), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n909), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n889), .A3(new_n911), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g495(.A1(new_n874), .A2(new_n876), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(new_n641), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  NOR2_X1   g498(.A1(G299), .A2(new_n631), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n622), .B1(new_n613), .B2(G92), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n630), .A2(new_n629), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n927), .A2(new_n623), .B1(new_n588), .B2(new_n593), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n923), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G299), .A2(new_n631), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n927), .A2(new_n593), .A3(new_n588), .A4(new_n623), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n922), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n924), .B2(new_n928), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n935), .B1(new_n922), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  XNOR2_X1  g517(.A(G290), .B(G288), .ZN(new_n943));
  XNOR2_X1  g518(.A(G166), .B(G305), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n935), .B(new_n947), .C1(new_n922), .C2(new_n940), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n942), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n942), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G868), .B2(new_n870), .ZN(G295));
  OAI21_X1  g527(.A(new_n951), .B1(G868), .B2(new_n870), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  INV_X1    g529(.A(new_n547), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n538), .A2(new_n539), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT75), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n538), .A2(KEYINPUT75), .A3(new_n539), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n564), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT78), .B1(new_n563), .B2(new_n564), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n957), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(G286), .A2(new_n565), .A3(new_n562), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n877), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n874), .A4(new_n876), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n933), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(KEYINPUT112), .A3(new_n969), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n921), .A2(new_n972), .A3(new_n965), .A4(new_n966), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n924), .A2(new_n928), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n976), .B2(new_n946), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n971), .A2(new_n934), .A3(new_n973), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n939), .A2(new_n968), .A3(new_n969), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n939), .A2(new_n968), .A3(KEYINPUT113), .A4(new_n969), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n945), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n977), .A2(new_n978), .A3(new_n985), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n928), .B(new_n924), .C1(new_n971), .C2(new_n973), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n945), .B1(new_n987), .B2(new_n970), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n978), .B1(new_n977), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n954), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n977), .A2(new_n988), .A3(new_n978), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n977), .B2(new_n985), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT44), .B(new_n991), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  AOI211_X1 g570(.A(KEYINPUT114), .B(new_n992), .C1(new_n977), .C2(new_n985), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n990), .B1(new_n995), .B2(new_n996), .ZN(G397));
  INV_X1    g572(.A(G1956), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n500), .B2(new_n505), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AND4_X1   g577(.A1(G40), .A2(new_n473), .A3(new_n479), .A4(new_n480), .ZN(new_n1003));
  NOR2_X1   g578(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(G164), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n998), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n588), .A2(new_n1009), .A3(new_n593), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n473), .A2(new_n479), .A3(G40), .A4(new_n480), .ZN(new_n1011));
  INV_X1    g586(.A(new_n505), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n498), .A2(new_n499), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G1384), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1011), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1000), .A2(new_n1017), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT56), .B(G2072), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1022), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1011), .B1(new_n1016), .B2(new_n1004), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1956), .B1(new_n1026), .B2(new_n1001), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1024), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT122), .B1(new_n1000), .B2(new_n1011), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1000), .A2(new_n1011), .A3(KEYINPUT122), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n811), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1348), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n631), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1023), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1003), .A2(new_n1016), .A3(new_n1038), .A4(new_n999), .ZN(new_n1039));
  AOI21_X1  g614(.A(G2067), .B1(new_n1039), .B2(new_n1030), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1348), .B1(new_n1026), .B2(new_n1001), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n637), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT60), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  OR4_X1    g618(.A1(KEYINPUT60), .A2(new_n1040), .A3(new_n1041), .A4(new_n631), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT61), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1028), .A2(new_n1023), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1028), .B2(new_n1023), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1043), .B(new_n1044), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT58), .B(G1341), .Z(new_n1049));
  NAND3_X1  g624(.A1(new_n1039), .A2(new_n1030), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1996), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1019), .A2(new_n1051), .A3(new_n1020), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n574), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT123), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1053), .A2(KEYINPUT123), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT59), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1059), .B2(new_n1055), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1037), .B1(new_n1048), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(G166), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n531), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n529), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT55), .B(G8), .C1(new_n1066), .C2(new_n521), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G2090), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1026), .A2(new_n1069), .A3(new_n1001), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1018), .B1(new_n500), .B2(new_n505), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1020), .A2(new_n1003), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1072), .B2(G1971), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1068), .B1(new_n1073), .B2(G8), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1073), .A2(G8), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1064), .A2(new_n1076), .A3(new_n1067), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1074), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1961), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1020), .A2(new_n807), .A3(new_n1003), .A4(new_n1071), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1019), .A2(KEYINPUT53), .A3(new_n807), .A4(new_n1020), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(KEYINPUT127), .A3(G171), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G171), .A2(KEYINPUT127), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1082), .A2(new_n1085), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(KEYINPUT54), .A3(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n597), .A2(new_n598), .A3(G1976), .A4(new_n599), .ZN(new_n1092));
  OAI211_X1 g667(.A(G8), .B(new_n1092), .C1(new_n1000), .C2(new_n1011), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1093), .A2(KEYINPUT118), .A3(KEYINPUT52), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT118), .B1(new_n1093), .B2(KEYINPUT52), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n762), .B2(G1976), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1094), .A2(new_n1095), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n611), .A2(G651), .B1(new_n613), .B2(G86), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n605), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1100), .B2(new_n605), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1000), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1063), .B1(new_n1105), .B2(new_n1003), .ZN(new_n1106));
  NAND2_X1  g681(.A1(G305), .A2(G1981), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(new_n1101), .A3(new_n605), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(KEYINPUT49), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1104), .A2(new_n1109), .A3(KEYINPUT119), .A4(new_n1106), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1098), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1080), .A2(new_n1091), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT126), .B(KEYINPUT54), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1087), .A2(G171), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1087), .A2(G171), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G2084), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1026), .A2(new_n1121), .A3(new_n1001), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n856), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT125), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n1122), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1129), .A3(G168), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n1063), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(G8), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(G286), .A2(G8), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1061), .A2(new_n1120), .A3(new_n1141), .ZN(new_n1142));
  AND4_X1   g717(.A1(G171), .A2(new_n1080), .A3(new_n1114), .A4(new_n1087), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1137), .A2(new_n1144), .A3(new_n1140), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1130), .A2(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT62), .B1(new_n1146), .B2(new_n1139), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1134), .A2(G286), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1080), .A2(new_n1114), .A3(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT121), .B(KEYINPUT63), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1080), .A2(new_n1114), .A3(new_n1153), .A4(new_n1149), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1114), .A2(new_n1075), .A3(new_n1079), .ZN(new_n1155));
  NOR2_X1   g730(.A1(G288), .A2(G1976), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT120), .Z(new_n1157));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1106), .B1(new_n1158), .B2(new_n1102), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1154), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1142), .A2(new_n1148), .A3(new_n1152), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1020), .A2(new_n1011), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1051), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT115), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n780), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1162), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n819), .B(new_n811), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n779), .A2(G1996), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n736), .B(new_n739), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT116), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1166), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1172), .B2(new_n1171), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(G290), .B(G1986), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1162), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1161), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n739), .ZN(new_n1179));
  NOR4_X1   g754(.A1(new_n1165), .A2(new_n1169), .A3(new_n1179), .A4(new_n736), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n819), .A2(G2067), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1162), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1166), .A2(G1986), .A3(G290), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1164), .A2(KEYINPUT46), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT115), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1163), .B(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT46), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n779), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1167), .A2(new_n1190), .ZN(new_n1191));
  OAI22_X1  g766(.A1(new_n1185), .A2(new_n1189), .B1(new_n1166), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1192), .A2(KEYINPUT47), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1192), .A2(KEYINPUT47), .ZN(new_n1194));
  OAI221_X1 g769(.A(new_n1182), .B1(new_n1175), .B2(new_n1184), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1178), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g772(.A1(G227), .A2(new_n464), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n1199), .B1(new_n724), .B2(new_n725), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1200), .B1(new_n684), .B2(new_n687), .ZN(new_n1201));
  OAI211_X1 g775(.A(new_n1201), .B(new_n919), .C1(new_n986), .C2(new_n989), .ZN(G225));
  INV_X1    g776(.A(G225), .ZN(G308));
endmodule


