

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U324 ( .A(n361), .B(n360), .Z(n292) );
  XOR2_X1 U325 ( .A(n384), .B(n393), .Z(n293) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n426) );
  XNOR2_X1 U327 ( .A(n427), .B(n426), .ZN(n448) );
  XNOR2_X1 U328 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n411) );
  XNOR2_X1 U329 ( .A(n362), .B(n292), .ZN(n363) );
  XNOR2_X1 U330 ( .A(n412), .B(n411), .ZN(n528) );
  XNOR2_X1 U331 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n295) );
  XNOR2_X1 U335 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U337 ( .A(G169GAT), .B(n296), .Z(n416) );
  XOR2_X1 U338 ( .A(G134GAT), .B(G99GAT), .Z(n298) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U341 ( .A(G183GAT), .B(G71GAT), .Z(n300) );
  XNOR2_X1 U342 ( .A(G176GAT), .B(KEYINPUT88), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U344 ( .A(n302), .B(n301), .Z(n312) );
  XOR2_X1 U345 ( .A(KEYINPUT87), .B(KEYINPUT84), .Z(n304) );
  XNOR2_X1 U346 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n310) );
  XOR2_X1 U348 ( .A(G15GAT), .B(G127GAT), .Z(n372) );
  XOR2_X1 U349 ( .A(G120GAT), .B(KEYINPUT0), .Z(n306) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n433) );
  XOR2_X1 U352 ( .A(n372), .B(n433), .Z(n308) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U357 ( .A(n416), .B(n313), .ZN(n476) );
  XNOR2_X1 U358 ( .A(G106GAT), .B(G78GAT), .ZN(n314) );
  XNOR2_X1 U359 ( .A(n314), .B(G148GAT), .ZN(n359) );
  XOR2_X1 U360 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n316) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n428) );
  XNOR2_X1 U363 ( .A(n359), .B(n428), .ZN(n329) );
  XOR2_X1 U364 ( .A(G22GAT), .B(G155GAT), .Z(n371) );
  XOR2_X1 U365 ( .A(G197GAT), .B(KEYINPUT21), .Z(n422) );
  XOR2_X1 U366 ( .A(n371), .B(n422), .Z(n318) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U369 ( .A(G50GAT), .B(G162GAT), .Z(n398) );
  XOR2_X1 U370 ( .A(n319), .B(n398), .Z(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT23), .B(G204GAT), .Z(n321) );
  XNOR2_X1 U372 ( .A(G218GAT), .B(G211GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U374 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n323) );
  XNOR2_X1 U375 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n472) );
  XOR2_X1 U380 ( .A(KEYINPUT70), .B(G8GAT), .Z(n331) );
  XNOR2_X1 U381 ( .A(G22GAT), .B(G197GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n347) );
  XOR2_X1 U383 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n333) );
  XNOR2_X1 U384 ( .A(G43GAT), .B(G29GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U386 ( .A(KEYINPUT8), .B(n334), .Z(n399) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XOR2_X1 U388 ( .A(G141GAT), .B(G15GAT), .Z(n336) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(G113GAT), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U391 ( .A(G36GAT), .B(G50GAT), .Z(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n399), .B(n341), .ZN(n345) );
  XOR2_X1 U395 ( .A(G1GAT), .B(KEYINPUT29), .Z(n343) );
  XNOR2_X1 U396 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n546) );
  XOR2_X1 U400 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n349) );
  XNOR2_X1 U401 ( .A(G120GAT), .B(KEYINPUT76), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n366) );
  INV_X1 U403 ( .A(KEYINPUT72), .ZN(n350) );
  NAND2_X1 U404 ( .A1(n350), .A2(G57GAT), .ZN(n353) );
  INV_X1 U405 ( .A(G57GAT), .ZN(n351) );
  NAND2_X1 U406 ( .A1(n351), .A2(KEYINPUT72), .ZN(n352) );
  NAND2_X1 U407 ( .A1(n353), .A2(n352), .ZN(n355) );
  XNOR2_X1 U408 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n384) );
  XOR2_X1 U410 ( .A(G99GAT), .B(G85GAT), .Z(n393) );
  NAND2_X1 U411 ( .A1(G230GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n293), .B(n356), .ZN(n364) );
  XOR2_X1 U413 ( .A(G64GAT), .B(G92GAT), .Z(n358) );
  XNOR2_X1 U414 ( .A(G176GAT), .B(G204GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n414) );
  XNOR2_X1 U416 ( .A(n359), .B(n414), .ZN(n362) );
  XOR2_X1 U417 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n361) );
  XNOR2_X1 U418 ( .A(KEYINPUT31), .B(KEYINPUT75), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n366), .B(n365), .ZN(n574) );
  XOR2_X1 U420 ( .A(KEYINPUT65), .B(KEYINPUT41), .Z(n367) );
  XOR2_X1 U421 ( .A(n574), .B(n367), .Z(n548) );
  OR2_X1 U422 ( .A1(n546), .A2(n548), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n368), .B(KEYINPUT46), .ZN(n403) );
  XOR2_X1 U424 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n370) );
  XNOR2_X1 U425 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n376) );
  XOR2_X1 U427 ( .A(n371), .B(G78GAT), .Z(n374) );
  XNOR2_X1 U428 ( .A(G1GAT), .B(n372), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U430 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U431 ( .A1(G231GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U433 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n380) );
  XNOR2_X1 U434 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U436 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U437 ( .A(G8GAT), .B(G183GAT), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n383), .B(G211GAT), .ZN(n413) );
  XNOR2_X1 U439 ( .A(n384), .B(n413), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n553) );
  XOR2_X1 U441 ( .A(n553), .B(KEYINPUT114), .Z(n561) );
  XOR2_X1 U442 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n392) );
  XOR2_X1 U443 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n388) );
  XNOR2_X1 U444 ( .A(G106GAT), .B(G92GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n390) );
  XNOR2_X1 U446 ( .A(G36GAT), .B(G190GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n389), .B(G218GAT), .ZN(n415) );
  XNOR2_X1 U448 ( .A(n390), .B(n415), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n397) );
  XOR2_X1 U450 ( .A(G134GAT), .B(KEYINPUT78), .Z(n429) );
  XOR2_X1 U451 ( .A(n393), .B(n429), .Z(n395) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U454 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n557) );
  INV_X1 U457 ( .A(n557), .ZN(n563) );
  NOR2_X1 U458 ( .A1(n561), .A2(n563), .ZN(n402) );
  NAND2_X1 U459 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n404), .B(KEYINPUT47), .ZN(n410) );
  XNOR2_X1 U461 ( .A(KEYINPUT36), .B(n557), .ZN(n583) );
  NOR2_X1 U462 ( .A1(n553), .A2(n583), .ZN(n406) );
  XNOR2_X1 U463 ( .A(KEYINPUT67), .B(KEYINPUT45), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n408) );
  NAND2_X1 U465 ( .A1(n546), .A2(n574), .ZN(n407) );
  NOR2_X1 U466 ( .A1(n408), .A2(n407), .ZN(n409) );
  NOR2_X1 U467 ( .A1(n410), .A2(n409), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n420) );
  XOR2_X1 U469 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n418) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U473 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n423) );
  XOR2_X1 U475 ( .A(n424), .B(n423), .Z(n466) );
  BUF_X1 U476 ( .A(n466), .Z(n520) );
  XOR2_X1 U477 ( .A(n520), .B(KEYINPUT120), .Z(n425) );
  NOR2_X1 U478 ( .A1(n528), .A2(n425), .ZN(n427) );
  XOR2_X1 U479 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U481 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U482 ( .A(n432), .B(KEYINPUT93), .Z(n435) );
  XNOR2_X1 U483 ( .A(n433), .B(KEYINPUT92), .ZN(n434) );
  XNOR2_X1 U484 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U485 ( .A(G85GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(G127GAT), .ZN(n436) );
  XNOR2_X1 U487 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U488 ( .A(n439), .B(n438), .Z(n447) );
  XOR2_X1 U489 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n441) );
  XNOR2_X1 U490 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U492 ( .A(G57GAT), .B(G155GAT), .Z(n443) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(G148GAT), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n447), .B(n446), .ZN(n517) );
  NOR2_X1 U497 ( .A1(n448), .A2(n517), .ZN(n449) );
  XOR2_X1 U498 ( .A(KEYINPUT66), .B(n449), .Z(n570) );
  NOR2_X1 U499 ( .A1(n472), .A2(n570), .ZN(n450) );
  XNOR2_X1 U500 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NOR2_X1 U501 ( .A1(n476), .A2(n451), .ZN(n564) );
  XNOR2_X1 U502 ( .A(KEYINPUT109), .B(n548), .ZN(n533) );
  NAND2_X1 U503 ( .A1(n564), .A2(n533), .ZN(n457) );
  XOR2_X1 U504 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n453) );
  XNOR2_X1 U505 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n455) );
  XOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT122), .Z(n454) );
  XOR2_X1 U508 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n459) );
  XNOR2_X1 U509 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U511 ( .A(KEYINPUT101), .B(n460), .Z(n482) );
  NOR2_X1 U512 ( .A1(n553), .A2(n563), .ZN(n461) );
  XNOR2_X1 U513 ( .A(KEYINPUT16), .B(n461), .ZN(n479) );
  INV_X1 U514 ( .A(n476), .ZN(n530) );
  AND2_X1 U515 ( .A1(n520), .A2(n530), .ZN(n462) );
  NOR2_X1 U516 ( .A1(n472), .A2(n462), .ZN(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(n463), .Z(n469) );
  XOR2_X1 U518 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n465) );
  NAND2_X1 U519 ( .A1(n472), .A2(n476), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n465), .B(n464), .ZN(n569) );
  XOR2_X1 U521 ( .A(n466), .B(KEYINPUT27), .Z(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT96), .ZN(n474) );
  NOR2_X1 U523 ( .A1(n569), .A2(n474), .ZN(n545) );
  XNOR2_X1 U524 ( .A(n545), .B(KEYINPUT98), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n517), .A2(n470), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n471), .B(KEYINPUT99), .ZN(n478) );
  INV_X1 U528 ( .A(n517), .ZN(n543) );
  XOR2_X1 U529 ( .A(n472), .B(KEYINPUT28), .Z(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT68), .B(n473), .Z(n524) );
  OR2_X1 U531 ( .A1(n474), .A2(n524), .ZN(n475) );
  NOR2_X1 U532 ( .A1(n543), .A2(n475), .ZN(n529) );
  NAND2_X1 U533 ( .A1(n529), .A2(n476), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n490) );
  NAND2_X1 U535 ( .A1(n479), .A2(n490), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n480), .B(KEYINPUT100), .ZN(n505) );
  INV_X1 U537 ( .A(n546), .ZN(n571) );
  NAND2_X1 U538 ( .A1(n571), .A2(n574), .ZN(n492) );
  NOR2_X1 U539 ( .A1(n505), .A2(n492), .ZN(n486) );
  NAND2_X1 U540 ( .A1(n486), .A2(n517), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(G1324GAT) );
  NAND2_X1 U542 ( .A1(n520), .A2(n486), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U545 ( .A1(n486), .A2(n530), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n486), .A2(n524), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT104), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(n488), .ZN(G1327GAT) );
  INV_X1 U550 ( .A(n553), .ZN(n577) );
  NOR2_X1 U551 ( .A1(n583), .A2(n577), .ZN(n489) );
  NAND2_X1 U552 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n491), .Z(n515) );
  NOR2_X1 U554 ( .A1(n492), .A2(n515), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n503), .A2(n517), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT105), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n498) );
  NAND2_X1 U561 ( .A1(n503), .A2(n520), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n501) );
  NAND2_X1 U565 ( .A1(n530), .A2(n503), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U567 ( .A(G43GAT), .B(n502), .Z(G1330GAT) );
  NAND2_X1 U568 ( .A1(n503), .A2(n524), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  NAND2_X1 U571 ( .A1(n546), .A2(n533), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n505), .A2(n514), .ZN(n511) );
  NAND2_X1 U573 ( .A1(n517), .A2(n511), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n520), .A2(n511), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n511), .A2(n530), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n509), .B(KEYINPUT110), .ZN(n510) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U581 ( .A1(n511), .A2(n524), .ZN(n512) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n519) );
  NOR2_X1 U584 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U585 ( .A(KEYINPUT111), .B(n516), .Z(n525) );
  NAND2_X1 U586 ( .A1(n517), .A2(n525), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n520), .A2(n525), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT113), .Z(n523) );
  NAND2_X1 U591 ( .A1(n525), .A2(n530), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U597 ( .A1(n528), .A2(n531), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n571), .A2(n540), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n535) );
  NAND2_X1 U601 ( .A1(n540), .A2(n533), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n538) );
  NAND2_X1 U605 ( .A1(n540), .A2(n561), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U609 ( .A1(n540), .A2(n563), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n528), .A2(n543), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n556) );
  NOR2_X1 U613 ( .A1(n546), .A2(n556), .ZN(n547) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  NOR2_X1 U615 ( .A1(n556), .A2(n548), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n550) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n556), .ZN(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT118), .B(n554), .Z(n555) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n571), .A2(n564), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n571), .A2(n578), .ZN(n572) );
  XOR2_X1 U638 ( .A(n573), .B(n572), .Z(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U640 ( .A(n578), .ZN(n582) );
  OR2_X1 U641 ( .A1(n582), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n581) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n585) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(n585), .B(n584), .Z(G1355GAT) );
endmodule

