//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n190), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(KEYINPUT75), .ZN(new_n194));
  NOR2_X1   g008(.A1(G119), .A2(G128), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G119), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G128), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT65), .A2(G119), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT65), .A2(G119), .ZN(new_n201));
  OAI21_X1  g015(.A(G128), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n195), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n198), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(KEYINPUT75), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(KEYINPUT23), .A3(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n200), .B2(new_n201), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n199), .A2(new_n206), .B1(new_n212), .B2(G110), .ZN(new_n213));
  INV_X1    g027(.A(G125), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G140), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G140), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT76), .B1(new_n219), .B2(G125), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(new_n214), .A3(G140), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n215), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n218), .B1(new_n223), .B2(new_n217), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G146), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n226), .B(new_n218), .C1(new_n223), .C2(new_n217), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n212), .A2(G110), .B1(new_n204), .B2(new_n205), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n214), .A2(G140), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n216), .A2(new_n230), .A3(new_n226), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n224), .B2(G146), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n213), .A2(new_n228), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n193), .B1(new_n233), .B2(KEYINPUT77), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n199), .A2(new_n206), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n212), .A2(G110), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n221), .B1(new_n214), .B2(G140), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n219), .A2(KEYINPUT76), .A3(G125), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n216), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT16), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n226), .B1(new_n240), .B2(new_n218), .ZN(new_n241));
  INV_X1    g055(.A(new_n227), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n235), .B(new_n236), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n229), .A2(new_n232), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n233), .A2(KEYINPUT77), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n234), .B1(new_n249), .B2(new_n193), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT25), .B1(new_n250), .B2(new_n188), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT77), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT77), .B1(new_n243), .B2(new_n244), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n193), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n234), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n189), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n189), .A2(G902), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G101), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT26), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G101), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT69), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT69), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g083(.A1(G237), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n266), .A2(G101), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n264), .A2(KEYINPUT26), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT69), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n271), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n263), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n272), .B1(new_n268), .B2(new_n269), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n271), .A3(new_n278), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n262), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G143), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT1), .B1(new_n285), .B2(G146), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(G146), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n226), .A2(G143), .ZN(new_n288));
  OAI211_X1 g102(.A(G128), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT11), .ZN(new_n290));
  INV_X1    g104(.A(G134), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(G137), .ZN(new_n292));
  INV_X1    g106(.A(G137), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT11), .A3(G134), .ZN(new_n294));
  INV_X1    g108(.A(G131), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(G137), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n292), .A2(new_n294), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n291), .A2(G137), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n293), .A2(G134), .ZN(new_n299));
  OAI21_X1  g113(.A(G131), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n226), .A2(G143), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n285), .A2(G146), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n301), .B(new_n302), .C1(KEYINPUT1), .C2(new_n208), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n289), .A2(new_n297), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n292), .A2(new_n294), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n299), .A2(G131), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n292), .A2(new_n294), .A3(new_n296), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n305), .A2(new_n306), .B1(new_n307), .B2(G131), .ZN(new_n308));
  AND2_X1   g122(.A1(KEYINPUT0), .A2(G128), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n301), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G143), .B(G146), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT0), .B(G128), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n304), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT65), .A2(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(G116), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n318), .A2(G116), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G113), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G113), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n321), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n321), .B2(new_n323), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n316), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n328), .ZN(new_n332));
  INV_X1    g146(.A(G116), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n200), .A2(new_n201), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n334), .B2(new_n322), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n321), .A2(new_n323), .A3(new_n328), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(KEYINPUT66), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n284), .B1(new_n315), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n304), .A2(KEYINPUT30), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n307), .A2(G131), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n313), .B1(new_n297), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT67), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n297), .ZN(new_n344));
  INV_X1    g158(.A(new_n313), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT30), .A4(new_n304), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n338), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n314), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n339), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n343), .A2(new_n348), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n350), .A3(new_n352), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT70), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n339), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n359), .A3(KEYINPUT31), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT31), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n339), .B(new_n361), .C1(new_n349), .C2(new_n353), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n357), .A2(KEYINPUT71), .A3(new_n361), .A4(new_n339), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n329), .A2(new_n330), .A3(new_n316), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT66), .B1(new_n335), .B2(new_n336), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n304), .B(new_n346), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n314), .A2(new_n337), .A3(new_n331), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT28), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT72), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n314), .B1(new_n337), .B2(new_n331), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(KEYINPUT28), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n369), .A2(KEYINPUT72), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n284), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n360), .A2(new_n366), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(G472), .A2(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT32), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n377), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT72), .B1(new_n369), .B2(new_n376), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT74), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n284), .B1(new_n371), .B2(KEYINPUT28), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT74), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n375), .A2(new_n389), .A3(new_n377), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n387), .A2(KEYINPUT29), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n369), .B1(new_n349), .B2(new_n353), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT29), .B1(new_n392), .B2(new_n284), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(KEYINPUT73), .A3(new_n375), .A4(new_n377), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n385), .A2(new_n386), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT73), .B1(new_n396), .B2(new_n388), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n188), .B(new_n391), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n381), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n383), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n398), .A2(G472), .B1(new_n380), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n261), .B1(new_n384), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G214), .B1(G237), .B2(G902), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT80), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(G234), .A2(G237), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(G952), .A3(new_n191), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT21), .B(G898), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(G902), .A3(G953), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G104), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT3), .B1(new_n413), .B2(G107), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n415));
  INV_X1    g229(.A(G107), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(G104), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(G107), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n420), .A3(G101), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(G101), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT78), .B(G101), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n423), .A2(new_n414), .A3(new_n417), .A4(new_n418), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(KEYINPUT4), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n331), .A2(new_n337), .A3(new_n421), .A4(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n334), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT81), .B1(new_n321), .B2(KEYINPUT5), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n321), .A2(KEYINPUT5), .A3(new_n323), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n430), .A2(new_n431), .A3(G113), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n413), .A2(G107), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n416), .A2(G104), .ZN(new_n435));
  OAI21_X1  g249(.A(G101), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n424), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n433), .A2(new_n336), .A3(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n426), .A2(new_n427), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n427), .B1(new_n426), .B2(new_n439), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G122), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT83), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n426), .A2(new_n439), .A3(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT6), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT84), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n289), .A2(new_n303), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n313), .A2(G125), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G224), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n453), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n449), .B2(new_n450), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n444), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n426), .A2(new_n439), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT82), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n426), .A2(new_n427), .A3(new_n439), .ZN(new_n462));
  INV_X1    g276(.A(new_n443), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n465));
  INV_X1    g279(.A(new_n446), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n447), .A2(new_n457), .A3(new_n459), .A4(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n442), .B(KEYINPUT8), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n430), .A2(new_n431), .A3(G113), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n432), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(new_n470), .B2(new_n471), .ZN(new_n474));
  AOI211_X1 g288(.A(new_n329), .B(new_n437), .C1(new_n472), .C2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n438), .B1(new_n433), .B2(new_n336), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI22_X1  g291(.A1(new_n454), .A2(new_n456), .B1(KEYINPUT7), .B2(new_n453), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n451), .A2(new_n479), .A3(new_n455), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n478), .A2(new_n445), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n468), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G210), .B1(G237), .B2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n468), .A2(new_n482), .A3(new_n484), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n412), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n425), .A2(new_n345), .A3(new_n421), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n424), .A2(new_n289), .A3(new_n303), .A4(new_n436), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(KEYINPUT10), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(KEYINPUT10), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n308), .B(new_n490), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT79), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G140), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n191), .A2(G227), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n495), .B1(new_n494), .B2(new_n498), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n437), .A2(new_n448), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n491), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT12), .B1(new_n502), .B2(new_n344), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n504), .B(new_n308), .C1(new_n501), .C2(new_n491), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n499), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n344), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n498), .B1(new_n509), .B2(new_n494), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n489), .B(new_n188), .C1(new_n507), .C2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n494), .A2(new_n498), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n494), .B1(new_n503), .B2(new_n505), .ZN(new_n513));
  INV_X1    g327(.A(new_n498), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n509), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G469), .B1(new_n515), .B2(G902), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G221), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT9), .B(G234), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n520), .B2(new_n188), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT87), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n223), .A2(new_n226), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n525), .A2(new_n231), .ZN(new_n526));
  INV_X1    g340(.A(G237), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n191), .A3(G214), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n285), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n270), .A2(G143), .A3(G214), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(KEYINPUT18), .A2(G131), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n528), .A2(new_n285), .ZN(new_n535));
  AOI21_X1  g349(.A(G143), .B1(new_n270), .B2(G214), .ZN(new_n536));
  OAI21_X1  g350(.A(G131), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n529), .A2(new_n295), .A3(new_n530), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n531), .A2(KEYINPUT17), .A3(G131), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n225), .A2(new_n540), .A3(new_n541), .A4(new_n227), .ZN(new_n542));
  XNOR2_X1  g356(.A(G113), .B(G122), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(new_n413), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n534), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT86), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n239), .A2(new_n546), .A3(KEYINPUT19), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT86), .B1(new_n223), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n216), .A2(new_n230), .A3(new_n548), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n547), .A2(new_n549), .A3(new_n226), .A4(new_n550), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n224), .A2(G146), .B1(new_n537), .B2(new_n539), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n544), .B1(new_n553), .B2(new_n534), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n524), .B1(new_n545), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(G475), .A2(G902), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n534), .A2(new_n542), .A3(new_n544), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n551), .A2(new_n552), .B1(new_n526), .B2(new_n533), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n557), .B(KEYINPUT87), .C1(new_n558), .C2(new_n544), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT20), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n557), .B1(new_n558), .B2(new_n544), .ZN(new_n562));
  NOR3_X1   g376(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G475), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n544), .B1(new_n534), .B2(new_n542), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n545), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n568), .B2(new_n188), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n208), .A2(G143), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT88), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n208), .A3(G143), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT88), .B1(new_n285), .B2(G128), .ZN(new_n576));
  AOI211_X1 g390(.A(G134), .B(new_n573), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n575), .ZN(new_n578));
  INV_X1    g392(.A(new_n573), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n291), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n572), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n574), .B1(new_n208), .B2(G143), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n285), .A2(KEYINPUT88), .A3(G128), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G134), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n578), .A2(new_n291), .A3(new_n579), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(KEYINPUT89), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G122), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G116), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n333), .A2(G122), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(G107), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT14), .B1(new_n588), .B2(G116), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT90), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT90), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n590), .A2(new_n595), .A3(KEYINPUT14), .ZN(new_n596));
  OR3_X1    g410(.A1(new_n588), .A2(KEYINPUT14), .A3(G116), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n594), .A2(new_n596), .A3(new_n597), .A4(new_n589), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n592), .B1(new_n598), .B2(G107), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n581), .A2(new_n587), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n573), .B(KEYINPUT13), .ZN(new_n601));
  INV_X1    g415(.A(new_n578), .ZN(new_n602));
  OAI21_X1  g416(.A(G134), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n591), .B(G107), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n586), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n519), .A2(new_n187), .A3(G953), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT91), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n600), .A2(new_n605), .A3(new_n607), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n606), .A2(KEYINPUT91), .A3(new_n608), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n188), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G478), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(KEYINPUT15), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(KEYINPUT15), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n620), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n612), .A2(new_n188), .A3(new_n613), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n523), .A2(new_n571), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n402), .A2(new_n488), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(new_n423), .Z(G3));
  INV_X1    g441(.A(new_n403), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n486), .B2(new_n487), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n615), .A2(G902), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n611), .A2(new_n610), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n607), .B1(new_n600), .B2(new_n605), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n613), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT93), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n606), .A2(new_n638), .A3(new_n608), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n611), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n634), .A2(new_n638), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT33), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n631), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n614), .A2(new_n615), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n560), .A2(KEYINPUT20), .B1(new_n562), .B2(new_n563), .ZN(new_n646));
  OAI22_X1  g460(.A1(new_n643), .A2(new_n645), .B1(new_n646), .B2(new_n569), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n629), .A2(new_n411), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n261), .A2(new_n523), .ZN(new_n650));
  INV_X1    g464(.A(G472), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n380), .B2(new_n188), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n381), .B2(new_n380), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  NAND2_X1  g471(.A1(new_n624), .A2(new_n570), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n555), .A2(new_n559), .A3(new_n563), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT94), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT94), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n555), .A2(new_n661), .A3(new_n559), .A4(new_n563), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n660), .A2(new_n662), .B1(KEYINPUT20), .B2(new_n560), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n629), .A2(new_n411), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n654), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n416), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(new_n193), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n245), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n259), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n258), .A2(KEYINPUT96), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT96), .ZN(new_n675));
  INV_X1    g489(.A(new_n189), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n254), .A2(new_n188), .A3(new_n255), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT25), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n676), .B1(new_n679), .B2(new_n256), .ZN(new_n680));
  INV_X1    g494(.A(new_n673), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n653), .A3(new_n625), .A4(new_n488), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  OR2_X1    g500(.A1(new_n410), .A2(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n407), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT97), .B1(new_n664), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT97), .ZN(new_n690));
  INV_X1    g504(.A(new_n688), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n658), .A2(new_n663), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n523), .B1(new_n401), .B2(new_n384), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n693), .A2(new_n629), .A3(new_n683), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NAND3_X1  g510(.A1(new_n571), .A2(new_n403), .A3(new_n624), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n683), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT98), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n521), .B1(new_n511), .B2(new_n516), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n688), .B(KEYINPUT39), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT40), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n380), .A2(new_n400), .ZN(new_n704));
  INV_X1    g518(.A(new_n359), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n358), .B1(new_n357), .B2(new_n339), .ZN(new_n706));
  INV_X1    g520(.A(new_n284), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n369), .B2(new_n370), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(G472), .B1(new_n709), .B2(G902), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT32), .B1(new_n380), .B2(new_n381), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n486), .A2(new_n487), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n714), .B(KEYINPUT38), .Z(new_n715));
  OR4_X1    g529(.A1(new_n699), .A2(new_n703), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(KEYINPUT99), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n647), .B2(new_n691), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n600), .A2(new_n605), .A3(new_n607), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n638), .B2(new_n634), .ZN(new_n721));
  INV_X1    g535(.A(new_n641), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n632), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT33), .B1(new_n612), .B2(new_n613), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n630), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n644), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n571), .A2(new_n726), .A3(KEYINPUT99), .A4(new_n688), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n719), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n629), .A3(new_n683), .A4(new_n694), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  NOR2_X1   g544(.A1(new_n500), .A2(new_n506), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n512), .A2(new_n495), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n510), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(G469), .B1(new_n733), .B2(G902), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n522), .A3(new_n511), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT100), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n734), .A2(KEYINPUT100), .A3(new_n522), .A4(new_n511), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n402), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n649), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT41), .B(G113), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  INV_X1    g557(.A(new_n665), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT101), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n745), .A3(new_n739), .A4(new_n402), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT101), .B1(new_n740), .B2(new_n665), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT102), .B(G116), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G18));
  NAND2_X1  g564(.A1(new_n401), .A2(new_n384), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n571), .A2(new_n624), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n683), .A2(new_n751), .A3(new_n411), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n754));
  INV_X1    g568(.A(new_n735), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n629), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n484), .B1(new_n468), .B2(new_n482), .ZN(new_n757));
  INV_X1    g571(.A(new_n487), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n755), .B(new_n403), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT103), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n753), .B1(new_n756), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n318), .ZN(G21));
  NAND3_X1  g576(.A1(new_n387), .A2(new_n372), .A3(new_n390), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT104), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT104), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n387), .A2(new_n765), .A3(new_n372), .A4(new_n390), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n284), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n360), .A2(new_n366), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n399), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n769), .A2(new_n261), .A3(new_n652), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n737), .A2(new_n411), .A3(new_n738), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n624), .A2(new_n403), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n569), .B1(new_n561), .B2(new_n564), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n758), .B2(new_n757), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n770), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G122), .ZN(G24));
  NOR2_X1   g592(.A1(new_n769), .A2(new_n652), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n683), .A3(new_n719), .A4(new_n727), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n760), .A2(new_n756), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G125), .ZN(G27));
  AND4_X1   g598(.A1(new_n486), .A2(new_n487), .A3(new_n403), .A4(new_n700), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT105), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(KEYINPUT42), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n728), .A2(new_n402), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n261), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n751), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n719), .A2(new_n727), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n486), .A2(new_n487), .A3(new_n403), .A4(new_n700), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G131), .ZN(G33));
  INV_X1    g611(.A(new_n663), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n569), .B1(new_n621), .B2(new_n623), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n688), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n690), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n664), .A2(KEYINPUT97), .A3(new_n688), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n402), .A2(new_n785), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT106), .B(G134), .Z(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G36));
  NAND2_X1  g619(.A1(new_n637), .A2(new_n642), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n806), .A2(new_n630), .B1(new_n615), .B2(new_n614), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n571), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(KEYINPUT43), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT107), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(KEYINPUT43), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT108), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n653), .B1(new_n682), .B2(new_n674), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT109), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n758), .A2(new_n757), .A3(new_n628), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n515), .A2(KEYINPUT45), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n515), .A2(KEYINPUT45), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(G469), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(G469), .A2(G902), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT46), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n511), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(KEYINPUT46), .A3(new_n824), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n521), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n701), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n820), .B(new_n830), .C1(new_n815), .C2(new_n816), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n818), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G137), .ZN(G39));
  XNOR2_X1  g647(.A(new_n829), .B(KEYINPUT47), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n820), .A2(new_n792), .A3(new_n751), .A4(new_n790), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  NOR3_X1   g651(.A1(new_n261), .A2(new_n711), .A3(new_n712), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n571), .A2(new_n807), .A3(new_n404), .A4(new_n521), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n734), .A2(new_n511), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT49), .Z(new_n841));
  NAND4_X1  g655(.A1(new_n715), .A2(new_n838), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n769), .A2(new_n261), .A3(new_n407), .A4(new_n652), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n813), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n715), .A2(new_n628), .A3(new_n755), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT50), .ZN(new_n847));
  INV_X1    g661(.A(new_n813), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n779), .A2(new_n683), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n819), .A2(new_n755), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT118), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n407), .B1(new_n850), .B2(KEYINPUT118), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n848), .A2(new_n849), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n851), .A2(new_n852), .A3(new_n838), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n571), .A2(new_n726), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n844), .A2(new_n820), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n521), .B1(new_n840), .B2(KEYINPUT116), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(KEYINPUT116), .B2(new_n840), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n834), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n847), .A2(KEYINPUT51), .A3(new_n857), .A4(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n848), .A2(new_n791), .A3(new_n853), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT48), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n813), .A2(new_n782), .A3(new_n843), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT119), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n855), .A2(new_n648), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(G952), .A3(new_n191), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n857), .A2(new_n870), .A3(new_n847), .A4(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n862), .B(new_n869), .C1(new_n872), .C2(KEYINPUT51), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n258), .A2(new_n700), .A3(new_n673), .A4(new_n688), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT113), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n680), .A2(new_n681), .A3(new_n691), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n700), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n713), .A2(new_n775), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n695), .A2(new_n729), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n780), .B1(new_n756), .B2(new_n760), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n875), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n694), .A2(new_n629), .A3(new_n683), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n693), .B2(new_n728), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n783), .A3(KEYINPUT114), .A4(new_n883), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT110), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n807), .B2(new_n773), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n571), .A2(new_n726), .A3(KEYINPUT110), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n773), .A2(KEYINPUT111), .A3(new_n624), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT111), .B1(new_n773), .B2(new_n624), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n894), .B(new_n895), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(new_n488), .A3(new_n653), .A4(new_n650), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n777), .A2(new_n899), .A3(new_n626), .A4(new_n684), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n741), .ZN(new_n901));
  INV_X1    g715(.A(new_n761), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n748), .A3(new_n902), .ZN(new_n903));
  NOR4_X1   g717(.A1(new_n663), .A2(new_n569), .A3(new_n624), .A4(new_n691), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n694), .A2(new_n819), .A3(new_n683), .A4(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT112), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(KEYINPUT112), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n803), .B1(new_n780), .B2(new_n793), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n796), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT52), .B1(new_n884), .B2(new_n885), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n892), .A2(new_n912), .A3(KEYINPUT53), .A4(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n886), .A2(KEYINPUT52), .A3(new_n889), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT52), .B1(new_n886), .B2(new_n889), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n900), .A2(new_n761), .A3(new_n741), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n909), .B1(new_n906), .B2(new_n907), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n918), .A3(new_n748), .A4(new_n796), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n915), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n874), .B(new_n914), .C1(new_n920), .C2(KEYINPUT53), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT115), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n892), .A2(new_n912), .A3(new_n913), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n916), .A2(new_n919), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n886), .A2(KEYINPUT52), .A3(new_n889), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(KEYINPUT53), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n874), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n892), .A2(new_n912), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n924), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT115), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n932), .A2(new_n933), .A3(new_n874), .A4(new_n914), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n873), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(G952), .A2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n842), .B1(new_n935), .B2(new_n936), .ZN(G75));
  NOR2_X1   g751(.A1(new_n191), .A2(G952), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT120), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n188), .B1(new_n932), .B2(new_n914), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT56), .B1(new_n941), .B2(G210), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n447), .A2(new_n459), .A3(new_n467), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n457), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT55), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n942), .A2(new_n945), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(G51));
  NAND2_X1  g762(.A1(new_n921), .A2(KEYINPUT121), .ZN(new_n949));
  INV_X1    g763(.A(new_n914), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT53), .B1(new_n926), .B2(new_n927), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT54), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n932), .A2(new_n953), .A3(new_n874), .A4(new_n914), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n824), .B(KEYINPUT57), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n510), .B2(new_n507), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n941), .A2(G469), .A3(new_n822), .A4(new_n821), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n938), .B1(new_n958), .B2(new_n959), .ZN(G54));
  NAND2_X1  g774(.A1(KEYINPUT58), .A2(G475), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT122), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n941), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n555), .A2(new_n559), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n965), .A2(new_n966), .A3(new_n938), .ZN(G60));
  XNOR2_X1  g781(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n615), .A2(new_n188), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n968), .B(new_n969), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n934), .B(new_n971), .C1(new_n922), .C2(new_n929), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n973));
  INV_X1    g787(.A(new_n806), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n974), .A2(new_n970), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n955), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n939), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(G63));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT60), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n932), .B2(new_n914), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n940), .B1(new_n984), .B2(new_n672), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n984), .A2(new_n250), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n985), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n987), .A2(new_n989), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(G66));
  NAND2_X1  g806(.A1(new_n903), .A2(new_n191), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT126), .Z(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n408), .B2(new_n452), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(G898), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n943), .B1(new_n997), .B2(G953), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n996), .B(new_n998), .Z(G69));
  NAND2_X1  g813(.A1(G900), .A2(G953), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n888), .A2(new_n783), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n829), .A2(new_n402), .A3(new_n701), .A4(new_n776), .ZN(new_n1002));
  AND4_X1   g816(.A1(new_n796), .A2(new_n836), .A3(new_n803), .A4(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n832), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1000), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n356), .A2(new_n352), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT127), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1006), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n716), .A2(new_n1001), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n791), .A2(new_n793), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n898), .A2(new_n701), .ZN(new_n1013));
  AOI22_X1  g827(.A1(new_n834), .A2(new_n835), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n832), .A2(new_n1011), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1009), .A2(G953), .ZN(new_n1017));
  AOI22_X1  g831(.A1(new_n1005), .A2(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  OAI21_X1  g836(.A(new_n1022), .B1(new_n1016), .B2(new_n903), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1023), .A2(new_n707), .A3(new_n392), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1022), .B1(new_n1004), .B2(new_n903), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n392), .A2(new_n707), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n938), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n925), .A2(new_n928), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1022), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n705), .A2(new_n706), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n392), .A2(new_n284), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1028), .B1(new_n1029), .B2(new_n1033), .ZN(G57));
endmodule


