

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770;

  INV_X1 U380 ( .A(n580), .ZN(n644) );
  NOR2_X2 U381 ( .A1(n765), .A2(n683), .ZN(n541) );
  XNOR2_X2 U382 ( .A(n525), .B(KEYINPUT35), .ZN(n765) );
  XNOR2_X2 U383 ( .A(n482), .B(n481), .ZN(n599) );
  XNOR2_X1 U384 ( .A(n418), .B(n417), .ZN(n580) );
  OR2_X1 U385 ( .A1(n730), .A2(G902), .ZN(n418) );
  NAND2_X2 U386 ( .A1(n644), .A2(n643), .ZN(n641) );
  AND2_X1 U387 ( .A1(n532), .A2(n531), .ZN(n683) );
  NAND2_X1 U388 ( .A1(n651), .A2(KEYINPUT31), .ZN(n420) );
  XNOR2_X1 U389 ( .A(n544), .B(KEYINPUT95), .ZN(n651) );
  NOR2_X1 U390 ( .A1(n543), .A2(n646), .ZN(n544) );
  AND2_X1 U391 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U392 ( .A(G146), .B(KEYINPUT68), .ZN(n414) );
  NAND2_X1 U393 ( .A1(n419), .A2(n421), .ZN(n554) );
  NOR2_X1 U394 ( .A1(n406), .A2(n405), .ZN(n419) );
  NAND2_X1 U395 ( .A1(n407), .A2(n425), .ZN(n406) );
  INV_X1 U396 ( .A(n750), .ZN(n434) );
  NAND2_X1 U397 ( .A1(n379), .A2(n567), .ZN(n378) );
  INV_X1 U398 ( .A(KEYINPUT33), .ZN(n467) );
  XNOR2_X1 U399 ( .A(n507), .B(G475), .ZN(n402) );
  OR2_X1 U400 ( .A1(n684), .A2(G902), .ZN(n403) );
  NAND2_X1 U401 ( .A1(n375), .A2(n611), .ZN(n374) );
  XNOR2_X1 U402 ( .A(n660), .B(n376), .ZN(n375) );
  INV_X1 U403 ( .A(KEYINPUT77), .ZN(n376) );
  AND2_X1 U404 ( .A1(n559), .A2(n681), .ZN(n560) );
  OR2_X1 U405 ( .A1(n719), .A2(n383), .ZN(n382) );
  NAND2_X1 U406 ( .A1(n436), .A2(n519), .ZN(n383) );
  XNOR2_X1 U407 ( .A(n463), .B(n462), .ZN(n470) );
  XNOR2_X1 U408 ( .A(n459), .B(n458), .ZN(n463) );
  XNOR2_X1 U409 ( .A(G122), .B(G107), .ZN(n509) );
  XNOR2_X1 U410 ( .A(n396), .B(KEYINPUT10), .ZN(n497) );
  XNOR2_X1 U411 ( .A(G125), .B(G140), .ZN(n396) );
  XNOR2_X1 U412 ( .A(n401), .B(n400), .ZN(n399) );
  XNOR2_X1 U413 ( .A(n496), .B(n495), .ZN(n400) );
  XNOR2_X1 U414 ( .A(n499), .B(n500), .ZN(n401) );
  XNOR2_X1 U415 ( .A(KEYINPUT12), .B(KEYINPUT98), .ZN(n495) );
  XNOR2_X1 U416 ( .A(G113), .B(G122), .ZN(n502) );
  XNOR2_X1 U417 ( .A(G146), .B(G143), .ZN(n501) );
  XNOR2_X1 U418 ( .A(G107), .B(G140), .ZN(n429) );
  XOR2_X1 U419 ( .A(G137), .B(KEYINPUT70), .Z(n438) );
  AND2_X1 U420 ( .A1(n409), .A2(n362), .ZN(n380) );
  INV_X1 U421 ( .A(KEYINPUT48), .ZN(n367) );
  AND2_X1 U422 ( .A1(n397), .A2(n373), .ZN(n372) );
  XNOR2_X1 U423 ( .A(G119), .B(G110), .ZN(n439) );
  XNOR2_X1 U424 ( .A(G146), .B(G128), .ZN(n442) );
  XNOR2_X1 U425 ( .A(n497), .B(n395), .ZN(n749) );
  INV_X1 U426 ( .A(n438), .ZN(n395) );
  XOR2_X1 U427 ( .A(KEYINPUT76), .B(KEYINPUT34), .Z(n493) );
  XNOR2_X1 U428 ( .A(n452), .B(KEYINPUT25), .ZN(n417) );
  XNOR2_X1 U429 ( .A(n528), .B(n527), .ZN(n533) );
  AND2_X1 U430 ( .A1(n627), .A2(n519), .ZN(n465) );
  XNOR2_X1 U431 ( .A(n521), .B(n520), .ZN(n551) );
  NOR2_X1 U432 ( .A1(n673), .A2(n672), .ZN(n677) );
  AND2_X1 U433 ( .A1(n640), .A2(n674), .ZN(n673) );
  AND2_X1 U434 ( .A1(n676), .A2(n364), .ZN(n387) );
  INV_X1 U435 ( .A(n420), .ZN(n405) );
  NAND2_X1 U436 ( .A1(n437), .A2(G902), .ZN(n385) );
  XOR2_X1 U437 ( .A(G119), .B(G113), .Z(n459) );
  XNOR2_X1 U438 ( .A(KEYINPUT88), .B(KEYINPUT72), .ZN(n458) );
  XNOR2_X1 U439 ( .A(G116), .B(KEYINPUT73), .ZN(n461) );
  XOR2_X1 U440 ( .A(KEYINPUT69), .B(G131), .Z(n500) );
  XOR2_X1 U441 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n496) );
  XOR2_X1 U442 ( .A(KEYINPUT102), .B(n553), .Z(n660) );
  INV_X1 U443 ( .A(KEYINPUT78), .ZN(n393) );
  XNOR2_X1 U444 ( .A(n371), .B(n370), .ZN(n369) );
  INV_X1 U445 ( .A(KEYINPUT46), .ZN(n370) );
  OR2_X1 U446 ( .A1(n763), .A2(n770), .ZN(n371) );
  XNOR2_X1 U447 ( .A(n414), .B(KEYINPUT4), .ZN(n433) );
  XNOR2_X1 U448 ( .A(KEYINPUT18), .B(G125), .ZN(n472) );
  XNOR2_X1 U449 ( .A(KEYINPUT89), .B(KEYINPUT17), .ZN(n473) );
  XNOR2_X1 U450 ( .A(n392), .B(n415), .ZN(n627) );
  XNOR2_X1 U451 ( .A(n509), .B(n377), .ZN(n510) );
  INV_X1 U452 ( .A(G116), .ZN(n377) );
  XNOR2_X1 U453 ( .A(n399), .B(n497), .ZN(n506) );
  XOR2_X1 U454 ( .A(KEYINPUT11), .B(G104), .Z(n503) );
  XNOR2_X1 U455 ( .A(n476), .B(n427), .ZN(n426) );
  XNOR2_X1 U456 ( .A(n428), .B(n438), .ZN(n427) );
  XNOR2_X1 U457 ( .A(n435), .B(n429), .ZN(n428) );
  AND2_X1 U458 ( .A1(n748), .A2(n363), .ZN(n388) );
  XNOR2_X1 U459 ( .A(KEYINPUT75), .B(KEYINPUT39), .ZN(n576) );
  NOR2_X1 U460 ( .A1(n597), .A2(n657), .ZN(n577) );
  NAND2_X1 U461 ( .A1(n545), .A2(KEYINPUT31), .ZN(n425) );
  NAND2_X1 U462 ( .A1(n423), .A2(n422), .ZN(n421) );
  NOR2_X1 U463 ( .A1(n545), .A2(KEYINPUT31), .ZN(n422) );
  NAND2_X1 U464 ( .A1(n381), .A2(n357), .ZN(n409) );
  NAND2_X1 U465 ( .A1(n413), .A2(n412), .ZN(n411) );
  OR2_X1 U466 ( .A1(n584), .A2(KEYINPUT19), .ZN(n412) );
  INV_X2 U467 ( .A(G953), .ZN(n755) );
  XNOR2_X1 U468 ( .A(n448), .B(n449), .ZN(n730) );
  XNOR2_X1 U469 ( .A(n540), .B(n539), .ZN(n766) );
  AND2_X1 U470 ( .A1(n551), .A2(n550), .ZN(n713) );
  AND2_X1 U471 ( .A1(n549), .A2(n548), .ZN(n698) );
  AND2_X1 U472 ( .A1(n677), .A2(n387), .ZN(n680) );
  XNOR2_X1 U473 ( .A(n708), .B(n416), .ZN(G48) );
  INV_X1 U474 ( .A(G146), .ZN(n416) );
  AND2_X1 U475 ( .A1(n584), .A2(KEYINPUT19), .ZN(n357) );
  XNOR2_X1 U476 ( .A(n403), .B(n402), .ZN(n552) );
  INV_X1 U477 ( .A(n552), .ZN(n550) );
  XOR2_X1 U478 ( .A(n457), .B(n456), .Z(n358) );
  XNOR2_X1 U479 ( .A(n368), .B(n367), .ZN(n748) );
  NOR2_X1 U480 ( .A1(n408), .A2(n411), .ZN(n359) );
  INV_X1 U481 ( .A(n436), .ZN(n437) );
  BUF_X1 U482 ( .A(n599), .Z(n391) );
  AND2_X1 U483 ( .A1(n498), .A2(G210), .ZN(n360) );
  NOR2_X1 U484 ( .A1(n611), .A2(n610), .ZN(n361) );
  AND2_X1 U485 ( .A1(n569), .A2(n490), .ZN(n362) );
  AND2_X1 U486 ( .A1(n717), .A2(n682), .ZN(n363) );
  AND2_X1 U487 ( .A1(n755), .A2(n638), .ZN(n364) );
  XOR2_X1 U488 ( .A(n634), .B(n633), .Z(n365) );
  NAND2_X2 U489 ( .A1(n384), .A2(n382), .ZN(n546) );
  NAND2_X1 U490 ( .A1(n389), .A2(n388), .ZN(n404) );
  XNOR2_X1 U491 ( .A(n366), .B(n571), .ZN(n572) );
  NAND2_X1 U492 ( .A1(n570), .A2(n584), .ZN(n366) );
  NAND2_X1 U493 ( .A1(n372), .A2(n369), .ZN(n368) );
  XNOR2_X1 U494 ( .A(n577), .B(n576), .ZN(n594) );
  XNOR2_X1 U495 ( .A(n562), .B(KEYINPUT85), .ZN(n379) );
  NOR2_X1 U496 ( .A1(n616), .A2(n361), .ZN(n373) );
  INV_X1 U497 ( .A(n660), .ZN(n613) );
  NAND2_X1 U498 ( .A1(n374), .A2(n614), .ZN(n398) );
  NOR2_X1 U499 ( .A1(n710), .A2(n713), .ZN(n553) );
  INV_X1 U500 ( .A(n389), .ZN(n739) );
  XNOR2_X2 U501 ( .A(n378), .B(KEYINPUT45), .ZN(n389) );
  NAND2_X1 U502 ( .A1(n390), .A2(n380), .ZN(n492) );
  INV_X1 U503 ( .A(n599), .ZN(n381) );
  NAND2_X1 U504 ( .A1(n719), .A2(n437), .ZN(n386) );
  XNOR2_X2 U505 ( .A(n392), .B(n426), .ZN(n719) );
  XNOR2_X2 U506 ( .A(n546), .B(KEYINPUT1), .ZN(n529) );
  XNOR2_X1 U507 ( .A(n464), .B(n358), .ZN(n415) );
  INV_X1 U508 ( .A(n411), .ZN(n390) );
  XNOR2_X2 U509 ( .A(n478), .B(n434), .ZN(n392) );
  XNOR2_X2 U510 ( .A(n394), .B(n393), .ZN(n543) );
  NOR2_X2 U511 ( .A1(n529), .A2(n641), .ZN(n394) );
  NAND2_X1 U512 ( .A1(n398), .A2(n615), .ZN(n397) );
  NAND2_X1 U513 ( .A1(n404), .A2(n617), .ZN(n619) );
  INV_X1 U514 ( .A(n404), .ZN(n624) );
  NAND2_X1 U515 ( .A1(n404), .A2(n675), .ZN(n676) );
  XNOR2_X1 U516 ( .A(n624), .B(KEYINPUT82), .ZN(n640) );
  INV_X1 U517 ( .A(n698), .ZN(n407) );
  INV_X1 U518 ( .A(n409), .ZN(n408) );
  NAND2_X1 U519 ( .A1(n410), .A2(n584), .ZN(n602) );
  INV_X1 U520 ( .A(n391), .ZN(n410) );
  NAND2_X1 U521 ( .A1(n599), .A2(n485), .ZN(n413) );
  NAND2_X1 U522 ( .A1(n533), .A2(n534), .ZN(n530) );
  AND2_X1 U523 ( .A1(n420), .A2(n425), .ZN(n424) );
  NAND2_X1 U524 ( .A1(n424), .A2(n421), .ZN(n709) );
  INV_X1 U525 ( .A(n651), .ZN(n423) );
  XNOR2_X2 U526 ( .A(n753), .B(G101), .ZN(n478) );
  XOR2_X1 U527 ( .A(n628), .B(KEYINPUT112), .Z(n430) );
  INV_X1 U528 ( .A(KEYINPUT3), .ZN(n460) );
  XNOR2_X1 U529 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U530 ( .A(n451), .B(KEYINPUT80), .ZN(n452) );
  INV_X1 U531 ( .A(n733), .ZN(n631) );
  INV_X1 U532 ( .A(KEYINPUT119), .ZN(n678) );
  AND2_X1 U533 ( .A1(n630), .A2(G953), .ZN(n733) );
  XNOR2_X2 U534 ( .A(G143), .B(KEYINPUT64), .ZN(n432) );
  INV_X1 U535 ( .A(G128), .ZN(n431) );
  XNOR2_X2 U536 ( .A(n432), .B(n431), .ZN(n508) );
  XNOR2_X2 U537 ( .A(n508), .B(n433), .ZN(n753) );
  XNOR2_X1 U538 ( .A(n500), .B(G134), .ZN(n750) );
  XNOR2_X1 U539 ( .A(G110), .B(G104), .ZN(n736) );
  XNOR2_X1 U540 ( .A(n736), .B(KEYINPUT74), .ZN(n476) );
  NAND2_X1 U541 ( .A1(G227), .A2(n755), .ZN(n435) );
  XOR2_X1 U542 ( .A(KEYINPUT71), .B(G469), .Z(n436) );
  XOR2_X1 U543 ( .A(KEYINPUT84), .B(KEYINPUT92), .Z(n440) );
  XNOR2_X1 U544 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U545 ( .A(n749), .B(n441), .ZN(n449) );
  XOR2_X1 U546 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n443) );
  XNOR2_X1 U547 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U548 ( .A(KEYINPUT23), .B(n444), .Z(n447) );
  NAND2_X1 U549 ( .A1(G234), .A2(n755), .ZN(n445) );
  XOR2_X1 U550 ( .A(KEYINPUT8), .B(n445), .Z(n515) );
  NAND2_X1 U551 ( .A1(G221), .A2(n515), .ZN(n446) );
  XNOR2_X1 U552 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U553 ( .A(KEYINPUT15), .B(G902), .ZN(n620) );
  NAND2_X1 U554 ( .A1(n620), .A2(G234), .ZN(n450) );
  XNOR2_X1 U555 ( .A(n450), .B(KEYINPUT20), .ZN(n453) );
  NAND2_X1 U556 ( .A1(G217), .A2(n453), .ZN(n451) );
  AND2_X1 U557 ( .A1(n453), .A2(G221), .ZN(n455) );
  XNOR2_X1 U558 ( .A(KEYINPUT93), .B(KEYINPUT21), .ZN(n454) );
  XNOR2_X1 U559 ( .A(n455), .B(n454), .ZN(n579) );
  INV_X1 U560 ( .A(n579), .ZN(n643) );
  XOR2_X1 U561 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n457) );
  XNOR2_X1 U562 ( .A(G137), .B(KEYINPUT79), .ZN(n456) );
  NOR2_X1 U563 ( .A1(G953), .A2(G237), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n470), .B(n360), .ZN(n464) );
  INV_X1 U565 ( .A(G902), .ZN(n519) );
  XNOR2_X2 U566 ( .A(n465), .B(G472), .ZN(n646) );
  INV_X1 U567 ( .A(KEYINPUT6), .ZN(n466) );
  XNOR2_X1 U568 ( .A(n646), .B(n466), .ZN(n582) );
  NOR2_X2 U569 ( .A1(n543), .A2(n582), .ZN(n468) );
  XNOR2_X1 U570 ( .A(n468), .B(n467), .ZN(n636) );
  XNOR2_X1 U571 ( .A(n509), .B(KEYINPUT16), .ZN(n469) );
  XNOR2_X1 U572 ( .A(n470), .B(n469), .ZN(n734) );
  NAND2_X1 U573 ( .A1(n755), .A2(G224), .ZN(n471) );
  XNOR2_X1 U574 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U575 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U576 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U578 ( .A(n479), .B(n734), .ZN(n691) );
  NAND2_X1 U579 ( .A1(n691), .A2(n620), .ZN(n482) );
  INV_X1 U580 ( .A(G237), .ZN(n480) );
  NAND2_X1 U581 ( .A1(n519), .A2(n480), .ZN(n483) );
  NAND2_X1 U582 ( .A1(n483), .A2(G210), .ZN(n481) );
  NAND2_X1 U583 ( .A1(n483), .A2(G214), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n484), .B(KEYINPUT90), .ZN(n584) );
  INV_X1 U585 ( .A(n584), .ZN(n656) );
  INV_X1 U586 ( .A(KEYINPUT19), .ZN(n485) );
  NAND2_X1 U587 ( .A1(G234), .A2(G237), .ZN(n486) );
  XNOR2_X1 U588 ( .A(n486), .B(KEYINPUT14), .ZN(n669) );
  INV_X1 U589 ( .A(G952), .ZN(n630) );
  NAND2_X1 U590 ( .A1(n755), .A2(n630), .ZN(n488) );
  NAND2_X1 U591 ( .A1(G953), .A2(n519), .ZN(n487) );
  AND2_X1 U592 ( .A1(n488), .A2(n487), .ZN(n489) );
  AND2_X1 U593 ( .A1(n669), .A2(n489), .ZN(n569) );
  NAND2_X1 U594 ( .A1(G953), .A2(G898), .ZN(n490) );
  INV_X1 U595 ( .A(KEYINPUT0), .ZN(n491) );
  XNOR2_X2 U596 ( .A(n492), .B(n491), .ZN(n549) );
  NAND2_X1 U597 ( .A1(n636), .A2(n549), .ZN(n494) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n524) );
  NAND2_X1 U599 ( .A1(G214), .A2(n498), .ZN(n499) );
  XNOR2_X1 U600 ( .A(n502), .B(n501), .ZN(n504) );
  XNOR2_X1 U601 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U602 ( .A(n506), .B(n505), .ZN(n684) );
  INV_X1 U603 ( .A(KEYINPUT13), .ZN(n507) );
  XNOR2_X1 U604 ( .A(n510), .B(KEYINPUT7), .ZN(n514) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n512) );
  XNOR2_X1 U606 ( .A(G134), .B(KEYINPUT99), .ZN(n511) );
  XNOR2_X1 U607 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U608 ( .A(n514), .B(n513), .Z(n517) );
  NAND2_X1 U609 ( .A1(G217), .A2(n515), .ZN(n516) );
  XNOR2_X1 U610 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U611 ( .A(n508), .B(n518), .ZN(n725) );
  NAND2_X1 U612 ( .A1(n725), .A2(n519), .ZN(n521) );
  XOR2_X1 U613 ( .A(KEYINPUT101), .B(G478), .Z(n520) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n522) );
  XNOR2_X1 U615 ( .A(KEYINPUT106), .B(n522), .ZN(n598) );
  XNOR2_X1 U616 ( .A(n598), .B(KEYINPUT81), .ZN(n523) );
  NAND2_X1 U617 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n658) );
  AND2_X1 U619 ( .A1(n658), .A2(n643), .ZN(n526) );
  NAND2_X1 U620 ( .A1(n549), .A2(n526), .ZN(n528) );
  INV_X1 U621 ( .A(KEYINPUT22), .ZN(n527) );
  BUF_X1 U622 ( .A(n529), .Z(n534) );
  XNOR2_X1 U623 ( .A(n530), .B(KEYINPUT105), .ZN(n532) );
  AND2_X1 U624 ( .A1(n646), .A2(n580), .ZN(n531) );
  AND2_X1 U625 ( .A1(n533), .A2(n582), .ZN(n558) );
  INV_X1 U626 ( .A(n534), .ZN(n535) );
  NOR2_X1 U627 ( .A1(n534), .A2(n644), .ZN(n536) );
  XNOR2_X1 U628 ( .A(KEYINPUT104), .B(n536), .ZN(n537) );
  NAND2_X1 U629 ( .A1(n558), .A2(n537), .ZN(n540) );
  INV_X1 U630 ( .A(KEYINPUT65), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n538), .B(KEYINPUT32), .ZN(n539) );
  NAND2_X1 U632 ( .A1(n541), .A2(n766), .ZN(n542) );
  NAND2_X1 U633 ( .A1(n542), .A2(KEYINPUT44), .ZN(n561) );
  INV_X1 U634 ( .A(n549), .ZN(n545) );
  BUF_X1 U635 ( .A(n546), .Z(n547) );
  NOR2_X1 U636 ( .A1(n547), .A2(n641), .ZN(n574) );
  AND2_X1 U637 ( .A1(n646), .A2(n574), .ZN(n548) );
  NOR2_X1 U638 ( .A1(n550), .A2(n551), .ZN(n710) );
  NAND2_X1 U639 ( .A1(n554), .A2(n660), .ZN(n556) );
  INV_X1 U640 ( .A(KEYINPUT103), .ZN(n555) );
  XNOR2_X1 U641 ( .A(n556), .B(n555), .ZN(n559) );
  AND2_X1 U642 ( .A1(n534), .A2(n644), .ZN(n557) );
  NAND2_X1 U643 ( .A1(n558), .A2(n557), .ZN(n681) );
  NAND2_X1 U644 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U645 ( .A1(n765), .A2(KEYINPUT44), .ZN(n563) );
  XNOR2_X1 U646 ( .A(n563), .B(KEYINPUT67), .ZN(n566) );
  INV_X1 U647 ( .A(n683), .ZN(n564) );
  AND2_X1 U648 ( .A1(n766), .A2(n564), .ZN(n565) );
  NAND2_X1 U649 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U650 ( .A1(G953), .A2(G900), .ZN(n568) );
  NAND2_X1 U651 ( .A1(n569), .A2(n568), .ZN(n578) );
  XOR2_X1 U652 ( .A(KEYINPUT30), .B(KEYINPUT107), .Z(n571) );
  INV_X1 U653 ( .A(n646), .ZN(n570) );
  NOR2_X1 U654 ( .A1(n578), .A2(n572), .ZN(n573) );
  NAND2_X1 U655 ( .A1(n574), .A2(n573), .ZN(n597) );
  INV_X1 U656 ( .A(KEYINPUT38), .ZN(n575) );
  XNOR2_X1 U657 ( .A(n391), .B(n575), .ZN(n657) );
  NAND2_X1 U658 ( .A1(n594), .A2(n713), .ZN(n717) );
  NOR2_X1 U659 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n581), .A2(n580), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n588), .A2(n582), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n710), .A2(n583), .ZN(n603) );
  NAND2_X1 U663 ( .A1(n584), .A2(n534), .ZN(n585) );
  NOR2_X1 U664 ( .A1(n603), .A2(n585), .ZN(n586) );
  XOR2_X1 U665 ( .A(n586), .B(KEYINPUT43), .Z(n587) );
  NAND2_X1 U666 ( .A1(n587), .A2(n391), .ZN(n682) );
  NOR2_X1 U667 ( .A1(n588), .A2(n646), .ZN(n589) );
  XOR2_X1 U668 ( .A(KEYINPUT28), .B(n589), .Z(n591) );
  XOR2_X1 U669 ( .A(n547), .B(KEYINPUT109), .Z(n590) );
  NOR2_X1 U670 ( .A1(n591), .A2(n590), .ZN(n607) );
  NOR2_X1 U671 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U672 ( .A1(n658), .A2(n661), .ZN(n592) );
  XNOR2_X1 U673 ( .A(KEYINPUT41), .B(n592), .ZN(n655) );
  AND2_X1 U674 ( .A1(n607), .A2(n655), .ZN(n593) );
  XNOR2_X1 U675 ( .A(n593), .B(KEYINPUT42), .ZN(n770) );
  AND2_X1 U676 ( .A1(n710), .A2(n594), .ZN(n596) );
  XNOR2_X1 U677 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n595) );
  XNOR2_X1 U678 ( .A(n596), .B(n595), .ZN(n763) );
  NOR2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n600), .A2(n410), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT108), .ZN(n768) );
  NOR2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT36), .B(n604), .Z(n605) );
  XNOR2_X1 U684 ( .A(n605), .B(KEYINPUT111), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n606), .A2(n535), .ZN(n716) );
  NAND2_X1 U686 ( .A1(n768), .A2(n716), .ZN(n616) );
  INV_X1 U687 ( .A(KEYINPUT47), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n607), .A2(n359), .ZN(n707) );
  NOR2_X1 U689 ( .A1(n707), .A2(KEYINPUT77), .ZN(n608) );
  NOR2_X1 U690 ( .A1(KEYINPUT83), .A2(n608), .ZN(n609) );
  NOR2_X1 U691 ( .A1(n613), .A2(n609), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(KEYINPUT83), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n707), .A2(n612), .ZN(n615) );
  INV_X1 U694 ( .A(KEYINPUT83), .ZN(n614) );
  NAND2_X1 U695 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n617) );
  INV_X1 U696 ( .A(n620), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n623) );
  INV_X1 U698 ( .A(KEYINPUT2), .ZN(n674) );
  NOR2_X1 U699 ( .A1(n620), .A2(n674), .ZN(n621) );
  OR2_X1 U700 ( .A1(n621), .A2(KEYINPUT66), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n624), .A2(KEYINPUT2), .ZN(n625) );
  AND2_X2 U703 ( .A1(n626), .A2(n625), .ZN(n718) );
  NAND2_X1 U704 ( .A1(n718), .A2(G472), .ZN(n629) );
  XOR2_X1 U705 ( .A(n627), .B(KEYINPUT62), .Z(n628) );
  XNOR2_X1 U706 ( .A(n629), .B(n430), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n635) );
  XOR2_X1 U708 ( .A(KEYINPUT87), .B(KEYINPUT113), .Z(n634) );
  XNOR2_X1 U709 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n635), .B(n365), .ZN(G57) );
  BUF_X1 U711 ( .A(n636), .Z(n637) );
  NAND2_X1 U712 ( .A1(n655), .A2(n637), .ZN(n638) );
  INV_X1 U713 ( .A(KEYINPUT82), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n534), .A2(n641), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n642), .B(KEYINPUT50), .ZN(n650) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(KEYINPUT49), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U719 ( .A(KEYINPUT117), .B(n648), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U722 ( .A(KEYINPUT51), .B(n653), .Z(n654) );
  NAND2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n666) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U726 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U728 ( .A1(n637), .A2(n664), .ZN(n665) );
  NAND2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n667) );
  XNOR2_X1 U731 ( .A(n668), .B(n667), .ZN(n671) );
  NAND2_X1 U732 ( .A1(n669), .A2(G952), .ZN(n670) );
  NOR2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U734 ( .A1(n674), .A2(n639), .ZN(n675) );
  XNOR2_X1 U735 ( .A(n678), .B(KEYINPUT53), .ZN(n679) );
  XNOR2_X1 U736 ( .A(n680), .B(n679), .ZN(G75) );
  XNOR2_X1 U737 ( .A(n681), .B(G101), .ZN(G3) );
  XNOR2_X1 U738 ( .A(n682), .B(G140), .ZN(G42) );
  XOR2_X1 U739 ( .A(n683), .B(G110), .Z(G12) );
  NAND2_X1 U740 ( .A1(n718), .A2(G475), .ZN(n686) );
  XNOR2_X1 U741 ( .A(n684), .B(KEYINPUT59), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U743 ( .A1(n687), .A2(n631), .ZN(n689) );
  INV_X1 U744 ( .A(KEYINPUT60), .ZN(n688) );
  XNOR2_X1 U745 ( .A(n689), .B(n688), .ZN(G60) );
  NAND2_X1 U746 ( .A1(n718), .A2(G210), .ZN(n693) );
  XOR2_X1 U747 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n690) );
  XNOR2_X1 U748 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U750 ( .A1(n694), .A2(n631), .ZN(n696) );
  INV_X1 U751 ( .A(KEYINPUT56), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n696), .B(n695), .ZN(G51) );
  NAND2_X1 U753 ( .A1(n698), .A2(n710), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n697), .B(G104), .ZN(G6) );
  XNOR2_X1 U755 ( .A(G107), .B(KEYINPUT26), .ZN(n702) );
  XOR2_X1 U756 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n700) );
  NAND2_X1 U757 ( .A1(n698), .A2(n713), .ZN(n699) );
  XNOR2_X1 U758 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U759 ( .A(n702), .B(n701), .ZN(G9) );
  INV_X1 U760 ( .A(n713), .ZN(n703) );
  NOR2_X1 U761 ( .A1(n707), .A2(n703), .ZN(n705) );
  XNOR2_X1 U762 ( .A(G128), .B(KEYINPUT29), .ZN(n704) );
  XNOR2_X1 U763 ( .A(n705), .B(n704), .ZN(G30) );
  INV_X1 U764 ( .A(n710), .ZN(n706) );
  NOR2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U766 ( .A1(n709), .A2(n710), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT116), .ZN(n712) );
  XNOR2_X1 U768 ( .A(G113), .B(n712), .ZN(G15) );
  NAND2_X1 U769 ( .A1(n709), .A2(n713), .ZN(n714) );
  XNOR2_X1 U770 ( .A(n714), .B(G116), .ZN(G18) );
  XOR2_X1 U771 ( .A(G125), .B(KEYINPUT37), .Z(n715) );
  XNOR2_X1 U772 ( .A(n716), .B(n715), .ZN(G27) );
  XNOR2_X1 U773 ( .A(G134), .B(n717), .ZN(G36) );
  BUF_X2 U774 ( .A(n718), .Z(n729) );
  NAND2_X1 U775 ( .A1(n729), .A2(G469), .ZN(n723) );
  XOR2_X1 U776 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n721) );
  XNOR2_X1 U777 ( .A(n719), .B(KEYINPUT120), .ZN(n720) );
  XNOR2_X1 U778 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U779 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n733), .A2(n724), .ZN(G54) );
  NAND2_X1 U781 ( .A1(n729), .A2(G478), .ZN(n727) );
  XNOR2_X1 U782 ( .A(n725), .B(KEYINPUT121), .ZN(n726) );
  XNOR2_X1 U783 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n733), .A2(n728), .ZN(G63) );
  NAND2_X1 U785 ( .A1(n729), .A2(G217), .ZN(n731) );
  XNOR2_X1 U786 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n733), .A2(n732), .ZN(G66) );
  NOR2_X1 U788 ( .A1(G898), .A2(n755), .ZN(n738) );
  XOR2_X1 U789 ( .A(G101), .B(n734), .Z(n735) );
  XNOR2_X1 U790 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U791 ( .A1(n738), .A2(n737), .ZN(n747) );
  NOR2_X1 U792 ( .A1(n739), .A2(G953), .ZN(n744) );
  NAND2_X1 U793 ( .A1(G953), .A2(G224), .ZN(n740) );
  XNOR2_X1 U794 ( .A(KEYINPUT61), .B(n740), .ZN(n741) );
  NAND2_X1 U795 ( .A1(n741), .A2(G898), .ZN(n742) );
  XOR2_X1 U796 ( .A(KEYINPUT122), .B(n742), .Z(n743) );
  NOR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U798 ( .A(KEYINPUT123), .B(n745), .ZN(n746) );
  XNOR2_X1 U799 ( .A(n747), .B(n746), .ZN(G69) );
  NAND2_X1 U800 ( .A1(n748), .A2(n363), .ZN(n754) );
  XNOR2_X1 U801 ( .A(n749), .B(KEYINPUT124), .ZN(n751) );
  XNOR2_X1 U802 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U803 ( .A(n753), .B(n752), .ZN(n757) );
  XNOR2_X1 U804 ( .A(n754), .B(n757), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n762) );
  XOR2_X1 U806 ( .A(G227), .B(n757), .Z(n758) );
  XNOR2_X1 U807 ( .A(n758), .B(KEYINPUT125), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(G900), .ZN(n760) );
  NAND2_X1 U809 ( .A1(G953), .A2(n760), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n762), .A2(n761), .ZN(G72) );
  XNOR2_X1 U811 ( .A(n763), .B(G131), .ZN(n764) );
  XNOR2_X1 U812 ( .A(n764), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U813 ( .A(n765), .B(G122), .Z(G24) );
  XNOR2_X1 U814 ( .A(n766), .B(G119), .ZN(n767) );
  XNOR2_X1 U815 ( .A(n767), .B(KEYINPUT126), .ZN(G21) );
  XOR2_X1 U816 ( .A(G143), .B(n768), .Z(n769) );
  XNOR2_X1 U817 ( .A(KEYINPUT115), .B(n769), .ZN(G45) );
  XOR2_X1 U818 ( .A(G137), .B(n770), .Z(G39) );
endmodule

