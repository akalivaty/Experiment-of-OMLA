

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  XNOR2_X1 U323 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n308) );
  XNOR2_X1 U324 ( .A(n325), .B(n308), .ZN(n310) );
  XNOR2_X1 U325 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n372) );
  XNOR2_X1 U326 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U327 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U328 ( .A(n320), .B(n319), .ZN(n321) );
  NOR2_X1 U329 ( .A1(n419), .A2(n525), .ZN(n458) );
  INV_X1 U330 ( .A(G218GAT), .ZN(n454) );
  XNOR2_X1 U331 ( .A(n451), .B(n450), .ZN(n541) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n457), .B(n456), .ZN(G1355GAT) );
  INV_X1 U334 ( .A(KEYINPUT54), .ZN(n396) );
  XOR2_X1 U335 ( .A(G43GAT), .B(G29GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(n293), .B(KEYINPUT67), .Z(n295) );
  XNOR2_X1 U339 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n359) );
  XOR2_X1 U341 ( .A(G113GAT), .B(G15GAT), .Z(n437) );
  XNOR2_X1 U342 ( .A(n359), .B(n437), .ZN(n299) );
  XOR2_X1 U343 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n297) );
  NAND2_X1 U344 ( .A1(G229GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n302) );
  XNOR2_X1 U347 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n300) );
  XOR2_X1 U348 ( .A(G1GAT), .B(KEYINPUT68), .Z(n338) );
  XNOR2_X1 U349 ( .A(n300), .B(n338), .ZN(n301) );
  XOR2_X1 U350 ( .A(n302), .B(n301), .Z(n304) );
  XOR2_X1 U351 ( .A(G141GAT), .B(G22GAT), .Z(n423) );
  XOR2_X1 U352 ( .A(G169GAT), .B(G8GAT), .Z(n378) );
  XNOR2_X1 U353 ( .A(n423), .B(n378), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n580) );
  XNOR2_X1 U355 ( .A(KEYINPUT69), .B(n580), .ZN(n542) );
  INV_X1 U356 ( .A(n542), .ZN(n470) );
  XOR2_X1 U357 ( .A(G78GAT), .B(G148GAT), .Z(n306) );
  XNOR2_X1 U358 ( .A(G106GAT), .B(G204GAT), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n426) );
  XNOR2_X1 U360 ( .A(G176GAT), .B(G92GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n307), .B(G64GAT), .ZN(n377) );
  XOR2_X1 U362 ( .A(n426), .B(n377), .Z(n322) );
  XOR2_X1 U363 ( .A(G57GAT), .B(KEYINPUT13), .Z(n325) );
  INV_X1 U364 ( .A(n310), .ZN(n309) );
  XOR2_X1 U365 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  NAND2_X1 U366 ( .A1(n309), .A2(n441), .ZN(n313) );
  INV_X1 U367 ( .A(n441), .ZN(n311) );
  NAND2_X1 U368 ( .A1(n311), .A2(n310), .ZN(n312) );
  NAND2_X1 U369 ( .A1(n313), .A2(n312), .ZN(n315) );
  NAND2_X1 U370 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n320) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n316), .B(KEYINPUT71), .ZN(n354) );
  XNOR2_X1 U374 ( .A(n354), .B(KEYINPUT70), .ZN(n318) );
  INV_X1 U375 ( .A(KEYINPUT32), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n469) );
  INV_X1 U377 ( .A(n469), .ZN(n367) );
  XOR2_X1 U378 ( .A(G127GAT), .B(G71GAT), .Z(n324) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(G183GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U381 ( .A(n326), .B(n325), .Z(n328) );
  XNOR2_X1 U382 ( .A(G22GAT), .B(G211GAT), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n342) );
  XOR2_X1 U384 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n330) );
  NAND2_X1 U385 ( .A1(G231GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U387 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n332) );
  XNOR2_X1 U388 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U390 ( .A(n334), .B(n333), .Z(n340) );
  XOR2_X1 U391 ( .A(G64GAT), .B(G78GAT), .Z(n336) );
  XNOR2_X1 U392 ( .A(G8GAT), .B(G155GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(n342), .B(n341), .Z(n577) );
  INV_X1 U397 ( .A(n577), .ZN(n587) );
  XOR2_X1 U398 ( .A(KEYINPUT72), .B(KEYINPUT74), .Z(n344) );
  XNOR2_X1 U399 ( .A(KEYINPUT73), .B(KEYINPUT75), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U401 ( .A(KEYINPUT11), .B(G162GAT), .Z(n346) );
  XNOR2_X1 U402 ( .A(G190GAT), .B(G134GAT), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(n348), .B(n347), .Z(n353) );
  XOR2_X1 U405 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n350) );
  NAND2_X1 U406 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(n351), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U410 ( .A(n354), .B(KEYINPUT65), .Z(n356) );
  XNOR2_X1 U411 ( .A(G218GAT), .B(G92GAT), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U413 ( .A(n358), .B(n357), .Z(n361) );
  XNOR2_X1 U414 ( .A(n359), .B(KEYINPUT9), .ZN(n360) );
  XOR2_X1 U415 ( .A(n361), .B(n360), .Z(n565) );
  XNOR2_X1 U416 ( .A(KEYINPUT36), .B(n565), .ZN(n498) );
  NAND2_X1 U417 ( .A1(n587), .A2(n498), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n362), .B(KEYINPUT111), .ZN(n363) );
  XOR2_X1 U419 ( .A(n363), .B(KEYINPUT45), .Z(n364) );
  NOR2_X1 U420 ( .A1(n367), .A2(n364), .ZN(n365) );
  XOR2_X1 U421 ( .A(KEYINPUT112), .B(n365), .Z(n366) );
  NOR2_X1 U422 ( .A1(n470), .A2(n366), .ZN(n375) );
  XOR2_X1 U423 ( .A(n367), .B(KEYINPUT41), .Z(n559) );
  NAND2_X1 U424 ( .A1(n559), .A2(n580), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n368), .B(KEYINPUT46), .ZN(n369) );
  NAND2_X1 U426 ( .A1(n369), .A2(n577), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n370), .B(KEYINPUT109), .ZN(n371) );
  INV_X1 U428 ( .A(n565), .ZN(n550) );
  NAND2_X1 U429 ( .A1(n371), .A2(n550), .ZN(n373) );
  NOR2_X1 U430 ( .A1(n375), .A2(n374), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n376), .B(KEYINPUT48), .ZN(n538) );
  XOR2_X1 U432 ( .A(n378), .B(n377), .Z(n380) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U435 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n382) );
  XNOR2_X1 U436 ( .A(G36GAT), .B(G204GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U438 ( .A(n384), .B(n383), .Z(n393) );
  XOR2_X1 U439 ( .A(KEYINPUT19), .B(G190GAT), .Z(n386) );
  XNOR2_X1 U440 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U442 ( .A(KEYINPUT17), .B(n387), .Z(n449) );
  XNOR2_X1 U443 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n388), .B(KEYINPUT21), .ZN(n389) );
  XOR2_X1 U445 ( .A(n389), .B(KEYINPUT88), .Z(n391) );
  XNOR2_X1 U446 ( .A(G197GAT), .B(G218GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n431) );
  XNOR2_X1 U448 ( .A(n449), .B(n431), .ZN(n392) );
  XOR2_X1 U449 ( .A(n393), .B(n392), .Z(n529) );
  INV_X1 U450 ( .A(n529), .ZN(n394) );
  NOR2_X1 U451 ( .A1(n538), .A2(n394), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n419) );
  XOR2_X1 U453 ( .A(G127GAT), .B(KEYINPUT0), .Z(n398) );
  XNOR2_X1 U454 ( .A(G134GAT), .B(KEYINPUT80), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n440) );
  XOR2_X1 U456 ( .A(G85GAT), .B(n440), .Z(n400) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(n401), .ZN(n418) );
  XOR2_X1 U460 ( .A(G148GAT), .B(G120GAT), .Z(n403) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(G113GAT), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n405) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U466 ( .A(n407), .B(n406), .Z(n416) );
  XOR2_X1 U467 ( .A(KEYINPUT2), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U468 ( .A(KEYINPUT89), .B(G155GAT), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U470 ( .A(KEYINPUT3), .B(n410), .Z(n432) );
  INV_X1 U471 ( .A(n432), .ZN(n414) );
  XOR2_X1 U472 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n412) );
  XNOR2_X1 U473 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U475 ( .A(n414), .B(n413), .Z(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U477 ( .A(n418), .B(n417), .Z(n482) );
  INV_X1 U478 ( .A(n482), .ZN(n525) );
  XOR2_X1 U479 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n421) );
  XNOR2_X1 U480 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U482 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U485 ( .A(n427), .B(n426), .Z(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT24), .B(KEYINPUT86), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n478) );
  XOR2_X1 U490 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n435) );
  XNOR2_X1 U491 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U493 ( .A(n436), .B(G99GAT), .Z(n439) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n445) );
  XOR2_X1 U496 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n451) );
  XOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT83), .Z(n447) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(KEYINPUT81), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  NOR2_X1 U504 ( .A1(n478), .A2(n541), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n452), .B(KEYINPUT26), .ZN(n554) );
  NAND2_X1 U506 ( .A1(n458), .A2(n554), .ZN(n453) );
  XNOR2_X1 U507 ( .A(KEYINPUT125), .B(n453), .ZN(n586) );
  NAND2_X1 U508 ( .A1(n586), .A2(n498), .ZN(n457) );
  XOR2_X1 U509 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n455) );
  INV_X1 U510 ( .A(G190GAT), .ZN(n465) );
  NAND2_X1 U511 ( .A1(n458), .A2(n478), .ZN(n460) );
  XOR2_X1 U512 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U514 ( .A1(n461), .A2(n541), .ZN(n576) );
  NOR2_X1 U515 ( .A1(n550), .A2(n576), .ZN(n463) );
  XNOR2_X1 U516 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  NOR2_X1 U519 ( .A1(n542), .A2(n576), .ZN(n466) );
  XNOR2_X1 U520 ( .A(n466), .B(KEYINPUT120), .ZN(n468) );
  INV_X1 U521 ( .A(G169GAT), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n468), .B(n467), .ZN(G1348GAT) );
  XOR2_X1 U523 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n489) );
  NAND2_X1 U524 ( .A1(n470), .A2(n469), .ZN(n501) );
  NAND2_X1 U525 ( .A1(n587), .A2(n550), .ZN(n471) );
  XNOR2_X1 U526 ( .A(n471), .B(KEYINPUT16), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT79), .ZN(n486) );
  XNOR2_X1 U528 ( .A(n529), .B(KEYINPUT27), .ZN(n476) );
  NAND2_X1 U529 ( .A1(n476), .A2(n525), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT95), .ZN(n555) );
  XOR2_X1 U531 ( .A(KEYINPUT28), .B(n478), .Z(n533) );
  INV_X1 U532 ( .A(n533), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n555), .A2(n474), .ZN(n539) );
  NOR2_X1 U534 ( .A1(n541), .A2(n539), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT96), .B(n475), .Z(n485) );
  NAND2_X1 U536 ( .A1(n554), .A2(n476), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n541), .A2(n529), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n478), .A2(n477), .ZN(n479) );
  XOR2_X1 U539 ( .A(KEYINPUT25), .B(n479), .Z(n480) );
  NAND2_X1 U540 ( .A1(n481), .A2(n480), .ZN(n483) );
  NAND2_X1 U541 ( .A1(n483), .A2(n482), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n485), .A2(n484), .ZN(n497) );
  NAND2_X1 U543 ( .A1(n486), .A2(n497), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT97), .B(n487), .Z(n512) );
  NOR2_X1 U545 ( .A1(n501), .A2(n512), .ZN(n495) );
  NAND2_X1 U546 ( .A1(n495), .A2(n525), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U548 ( .A(G1GAT), .B(n490), .Z(G1324GAT) );
  XOR2_X1 U549 ( .A(G8GAT), .B(KEYINPUT99), .Z(n492) );
  NAND2_X1 U550 ( .A1(n495), .A2(n529), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U553 ( .A1(n495), .A2(n541), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n533), .A2(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .Z(n504) );
  NAND2_X1 U558 ( .A1(n498), .A2(n497), .ZN(n499) );
  NOR2_X1 U559 ( .A1(n587), .A2(n499), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT37), .B(n500), .ZN(n524) );
  NOR2_X1 U561 ( .A1(n501), .A2(n524), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(KEYINPUT38), .ZN(n508) );
  NAND2_X1 U563 ( .A1(n525), .A2(n508), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NAND2_X1 U565 ( .A1(n508), .A2(n529), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n508), .A2(n541), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(KEYINPUT40), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n510) );
  NAND2_X1 U571 ( .A1(n508), .A2(n533), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  XNOR2_X1 U574 ( .A(KEYINPUT102), .B(KEYINPUT42), .ZN(n516) );
  XOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT103), .Z(n514) );
  INV_X1 U576 ( .A(n559), .ZN(n570) );
  OR2_X1 U577 ( .A1(n570), .A2(n580), .ZN(n523) );
  NOR2_X1 U578 ( .A1(n512), .A2(n523), .ZN(n519) );
  NAND2_X1 U579 ( .A1(n519), .A2(n525), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n529), .A2(n519), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n541), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n518), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U587 ( .A1(n519), .A2(n533), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(n522), .ZN(G1335GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n527) );
  NOR2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n534), .A2(n525), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  XOR2_X1 U595 ( .A(G92GAT), .B(KEYINPUT107), .Z(n531) );
  NAND2_X1 U596 ( .A1(n534), .A2(n529), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n541), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n536) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U603 ( .A(G106GAT), .B(n537), .Z(G1339GAT) );
  NOR2_X1 U604 ( .A1(n538), .A2(n539), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n542), .A2(n549), .ZN(n543) );
  XOR2_X1 U607 ( .A(G113GAT), .B(n543), .Z(G1340GAT) );
  NOR2_X1 U608 ( .A1(n570), .A2(n549), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U611 ( .A1(n577), .A2(n549), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT113), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  NOR2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U616 ( .A(KEYINPUT51), .B(KEYINPUT114), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  XOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT115), .Z(n558) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U621 ( .A1(n538), .A2(n556), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n566), .A2(n580), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n561) );
  NAND2_X1 U625 ( .A1(n566), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n587), .A2(n566), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT116), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n564), .ZN(G1346GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n568) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n576), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n572) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT121), .B(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1349GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U642 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1350GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  NAND2_X1 U645 ( .A1(n586), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n586), .A2(n367), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
endmodule

