//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1206, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  AND2_X1   g0008(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT66), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(new_n211), .A2(new_n212), .B1(G77), .B2(G244), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G50), .A2(G226), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G68), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n217), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(G58), .A2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n206), .B(new_n226), .C1(new_n229), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n246), .B(KEYINPUT68), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT69), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT70), .B(G107), .ZN(new_n249));
  INV_X1    g0049(.A(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n248), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G169), .ZN(new_n255));
  INV_X1    g0055(.A(new_n227), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G238), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT71), .B(G45), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n259), .B(G274), .C1(new_n263), .C2(G41), .ZN(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G232), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G226), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n268), .A2(new_n271), .B1(G33), .B2(G97), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n262), .B(new_n264), .C1(new_n272), .C2(new_n258), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT13), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n271), .B1(G232), .B2(new_n270), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G97), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(new_n262), .A4(new_n264), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n255), .B1(new_n274), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(KEYINPUT78), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n274), .A2(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G179), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n285), .A2(KEYINPUT77), .A3(KEYINPUT78), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT14), .B1(new_n285), .B2(KEYINPUT77), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n287), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n227), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n259), .B2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G68), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT12), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(G68), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n297), .A2(new_n300), .A3(G1), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n222), .A2(new_n301), .A3(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G20), .A2(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G50), .ZN(new_n305));
  INV_X1    g0105(.A(G77), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n228), .A2(G33), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT64), .B(G68), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n305), .B1(new_n306), .B2(new_n307), .C1(new_n308), .C2(new_n228), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n294), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n310), .A2(KEYINPUT76), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(KEYINPUT76), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT11), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT11), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n303), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n292), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n288), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n288), .A2(G190), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n231), .B2(G50), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  INV_X1    g0126(.A(new_n304), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n325), .B1(new_n326), .B2(new_n327), .C1(new_n307), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G50), .ZN(new_n330));
  INV_X1    g0130(.A(new_n298), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n329), .A2(new_n294), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n295), .A2(G50), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n265), .A2(new_n266), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n270), .A2(G222), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G223), .A2(G1698), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n281), .C1(G77), .C2(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n261), .A2(G226), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n264), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n255), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n334), .B(new_n342), .C1(G179), .C2(new_n341), .ZN(new_n343));
  XOR2_X1   g0143(.A(new_n343), .B(KEYINPUT72), .Z(new_n344));
  NAND2_X1  g0144(.A1(new_n331), .A2(new_n306), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n295), .A2(G77), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT8), .B(G58), .Z(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n304), .B1(G20), .B2(G77), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT15), .B(G87), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n307), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n350), .A2(KEYINPUT74), .A3(new_n294), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT74), .B1(new_n350), .B2(new_n294), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n345), .B(new_n346), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G238), .A2(G1698), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n335), .B(new_n354), .C1(new_n267), .C2(G1698), .ZN(new_n355));
  OR2_X1    g0155(.A1(KEYINPUT73), .A2(G107), .ZN(new_n356));
  NAND2_X1  g0156(.A1(KEYINPUT73), .A2(G107), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n355), .B(new_n281), .C1(new_n335), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n261), .A2(G244), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n264), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n353), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n344), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n341), .A2(G200), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT75), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n341), .A2(new_n364), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n334), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n370), .B(new_n373), .C1(new_n372), .C2(new_n334), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n368), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n362), .A2(G179), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n362), .A2(new_n255), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n353), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n328), .A2(new_n298), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n295), .B2(new_n328), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n265), .A2(new_n228), .A3(new_n266), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n275), .A2(new_n276), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n386), .B2(new_n228), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G58), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n231), .B1(new_n222), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(G20), .B1(G159), .B2(new_n304), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n294), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n308), .B1(new_n385), .B2(new_n387), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT16), .B1(new_n394), .B2(new_n391), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n382), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n269), .A2(G1698), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n397), .B1(G223), .B2(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n281), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n261), .A2(G232), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n264), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G169), .ZN(new_n404));
  INV_X1    g0204(.A(G179), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n396), .A2(KEYINPUT18), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n396), .A2(new_n406), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n396), .A2(KEYINPUT79), .A3(new_n406), .A4(KEYINPUT18), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n401), .A2(new_n364), .A3(new_n264), .A4(new_n402), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT80), .ZN(new_n417));
  INV_X1    g0217(.A(G274), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT71), .B(G45), .Z(new_n419));
  INV_X1    g0219(.A(G41), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n400), .A2(new_n281), .B1(new_n421), .B2(new_n259), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT80), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n364), .A4(new_n402), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n403), .A2(new_n320), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n417), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n415), .B1(new_n426), .B2(new_n396), .ZN(new_n427));
  INV_X1    g0227(.A(new_n382), .ZN(new_n428));
  INV_X1    g0228(.A(new_n294), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n230), .B1(new_n308), .B2(G58), .ZN(new_n430));
  INV_X1    g0230(.A(G159), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n430), .A2(new_n228), .B1(new_n431), .B2(new_n327), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n383), .A2(new_n384), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n386), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n218), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n429), .B1(new_n436), .B2(KEYINPUT16), .ZN(new_n437));
  INV_X1    g0237(.A(new_n395), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n428), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n417), .A2(new_n424), .A3(new_n425), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(KEYINPUT17), .A3(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n427), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n414), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n324), .A2(new_n377), .A3(new_n380), .A4(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n259), .A2(new_n250), .A3(G13), .A4(G20), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n259), .A2(G33), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n429), .A2(new_n298), .A3(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n293), .A2(new_n227), .B1(G20), .B2(new_n250), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(new_n228), .C1(G33), .C2(new_n279), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT20), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n446), .B1(new_n448), .B2(new_n250), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G303), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n265), .A2(new_n455), .A3(new_n266), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G264), .A2(G1698), .ZN(new_n457));
  INV_X1    g0257(.A(G257), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(G1698), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n456), .B(new_n281), .C1(new_n386), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n462), .B(G274), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n462), .B1(new_n464), .B2(new_n463), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G270), .A3(new_n258), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n460), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n460), .A2(new_n467), .A3(KEYINPUT84), .A4(new_n465), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n454), .A2(new_n470), .A3(G169), .A4(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT21), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n470), .A2(new_n471), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G200), .ZN(new_n475));
  INV_X1    g0275(.A(new_n454), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n476), .C1(new_n364), .C2(new_n474), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n468), .A2(new_n405), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n454), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n473), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1698), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(G244), .C1(new_n276), .C2(new_n275), .ZN(new_n483));
  INV_X1    g0283(.A(G244), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n265), .B2(new_n266), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(new_n450), .C1(new_n485), .C2(KEYINPUT4), .ZN(new_n486));
  OAI21_X1  g0286(.A(G250), .B1(new_n275), .B2(new_n276), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n270), .B1(new_n487), .B2(KEYINPUT4), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n281), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n466), .A2(G257), .A3(new_n258), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n465), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n493), .A3(new_n465), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G200), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n359), .B1(new_n385), .B2(new_n387), .ZN(new_n497));
  INV_X1    g0297(.A(G107), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT6), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(KEYINPUT81), .ZN(new_n502));
  OAI211_X1 g0302(.A(G97), .B(new_n498), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(KEYINPUT81), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n279), .A2(G107), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G20), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n327), .A2(new_n306), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n497), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n513), .A2(new_n294), .B1(new_n279), .B2(new_n331), .ZN(new_n514));
  INV_X1    g0314(.A(new_n448), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G97), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n489), .A2(new_n492), .A3(G190), .A4(new_n494), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n496), .A2(new_n514), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n331), .A2(new_n279), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n358), .B1(new_n433), .B2(new_n434), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n228), .B1(new_n503), .B2(new_n508), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n520), .A2(new_n521), .A3(new_n511), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n516), .B(new_n519), .C1(new_n522), .C2(new_n429), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n495), .A2(new_n255), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n489), .A2(new_n492), .A3(new_n405), .A4(new_n494), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n307), .B2(new_n279), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n228), .B(G68), .C1(new_n275), .C2(new_n276), .ZN(new_n530));
  INV_X1    g0330(.A(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n279), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n356), .B2(new_n357), .ZN(new_n533));
  NAND3_X1  g0333(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n534), .A2(new_n228), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n529), .B(new_n530), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n294), .ZN(new_n537));
  INV_X1    g0337(.A(new_n349), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n515), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n349), .A2(new_n331), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n223), .A2(new_n270), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n484), .A2(G1698), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n275), .C2(new_n276), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n258), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(G250), .B1(new_n461), .B2(G1), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n259), .A2(G45), .A3(G274), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n547), .A2(new_n548), .B1(new_n256), .B2(new_n257), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n405), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n255), .B1(new_n546), .B2(new_n549), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n541), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n536), .A2(new_n294), .B1(new_n331), .B2(new_n349), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n515), .A2(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n544), .A2(new_n545), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n281), .ZN(new_n557));
  INV_X1    g0357(.A(new_n549), .ZN(new_n558));
  AOI21_X1  g0358(.A(G200), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n546), .A2(G190), .A3(new_n549), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n554), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT83), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT83), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n553), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n527), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT23), .B1(new_n498), .B2(G20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n545), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n567), .B1(new_n358), .B2(KEYINPUT23), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(new_n228), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n228), .B(G87), .C1(new_n275), .C2(new_n276), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT22), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n335), .A2(KEYINPUT22), .A3(new_n228), .A4(G87), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n570), .A2(KEYINPUT24), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  AND2_X1   g0376(.A1(KEYINPUT73), .A2(G107), .ZN(new_n577));
  NOR2_X1   g0377(.A1(KEYINPUT73), .A2(G107), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT23), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n567), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(G20), .B1(new_n545), .B2(new_n567), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n573), .A2(new_n574), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n576), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(new_n584), .A3(new_n294), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n515), .A2(G107), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n298), .A2(G107), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT25), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  OR2_X1    g0389(.A1(G250), .A2(G1698), .ZN(new_n590));
  OAI221_X1 g0390(.A(new_n590), .B1(G257), .B2(new_n270), .C1(new_n275), .C2(new_n276), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n466), .A2(new_n258), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n281), .A2(new_n593), .B1(new_n594), .B2(G264), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT85), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n465), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n466), .A2(G264), .A3(new_n258), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n265), .A2(new_n266), .B1(new_n458), .B2(G1698), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n590), .B1(G33), .B2(G294), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n465), .B(new_n598), .C1(new_n600), .C2(new_n258), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT85), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n364), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n320), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n589), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(new_n595), .B2(new_n465), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n601), .A2(KEYINPUT85), .ZN(new_n607));
  OAI21_X1  g0407(.A(G169), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n601), .A2(new_n405), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(KEYINPUT86), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n255), .B1(new_n597), .B2(new_n602), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n609), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n605), .B1(new_n615), .B2(new_n589), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n445), .A2(new_n480), .A3(new_n566), .A4(new_n616), .ZN(G372));
  AND3_X1   g0417(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n564), .B1(new_n553), .B2(new_n561), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n553), .A2(new_n561), .A3(new_n564), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(KEYINPUT26), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT88), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n553), .A2(new_n561), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n563), .A2(new_n565), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT26), .A4(new_n618), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n622), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n553), .B(KEYINPUT87), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n518), .A2(new_n526), .A3(new_n623), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(new_n605), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n589), .B1(new_n613), .B2(new_n609), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n473), .A2(new_n634), .A3(new_n479), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n445), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n344), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n412), .A2(new_n407), .ZN(new_n640));
  INV_X1    g0440(.A(new_n380), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n292), .A2(new_n318), .B1(new_n323), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n442), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n376), .A2(new_n375), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n638), .A2(new_n646), .ZN(G369));
  NAND2_X1  g0447(.A1(new_n473), .A2(new_n479), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n259), .A2(new_n228), .A3(G13), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n476), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n648), .A2(KEYINPUT89), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n648), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n473), .A2(new_n477), .A3(new_n479), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT89), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n657), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n589), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n616), .B1(new_n663), .B2(new_n655), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n611), .B2(new_n614), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n654), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n662), .A2(G330), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n634), .A2(new_n654), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n654), .B1(new_n473), .B2(new_n479), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n616), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n204), .ZN(new_n673));
  OR3_X1    g0473(.A1(new_n673), .A2(KEYINPUT90), .A3(G41), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT90), .B1(new_n673), .B2(G41), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n533), .A2(new_n250), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n232), .B2(new_n676), .ZN(new_n680));
  XOR2_X1   g0480(.A(KEYINPUT91), .B(KEYINPUT92), .Z(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n680), .B(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n633), .B1(new_n665), .B2(new_n648), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n627), .A2(new_n625), .A3(new_n618), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n631), .B(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n684), .A2(new_n685), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n655), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n616), .A2(new_n566), .A3(new_n480), .A4(new_n655), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n478), .A2(new_n595), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n489), .A2(new_n492), .A3(new_n550), .A4(new_n494), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  OR3_X1    g0495(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n557), .A2(new_n558), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n595), .A2(new_n465), .B1(new_n697), .B2(KEYINPUT93), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT93), .ZN(new_n699));
  AOI21_X1  g0499(.A(G179), .B1(new_n550), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n474), .A2(new_n698), .A3(new_n495), .A4(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n695), .B1(new_n693), .B2(new_n694), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n654), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n692), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n654), .B1(new_n630), .B2(new_n636), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n691), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT95), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n713), .B(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n683), .B1(new_n715), .B2(G1), .ZN(G364));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n660), .A2(new_n658), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n717), .B(G330), .C1(new_n718), .C2(new_n657), .ZN(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT96), .B1(new_n661), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n676), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n300), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n259), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n722), .B(new_n728), .C1(G330), .C2(new_n662), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n728), .B1(new_n661), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n227), .B1(G20), .B2(new_n255), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n405), .A2(new_n320), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n228), .A2(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G317), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT33), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n739), .A2(KEYINPUT33), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G329), .ZN(new_n746));
  INV_X1    g0546(.A(G283), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n320), .A2(G179), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n736), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n742), .B(new_n746), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(G20), .A2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n735), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(G326), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n748), .A2(new_n752), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G303), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n405), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n752), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n335), .B1(new_n761), .B2(G322), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n228), .B1(new_n743), .B2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G294), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n755), .A2(new_n758), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n736), .A2(new_n759), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(G311), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n737), .A2(new_n218), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n763), .A2(new_n279), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n386), .B(new_n771), .C1(G77), .C2(new_n768), .ZN(new_n772));
  INV_X1    g0572(.A(new_n749), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G107), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n744), .A2(new_n431), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G50), .A2(new_n754), .B1(new_n757), .B2(G87), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n772), .A2(new_n774), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n770), .B(new_n778), .C1(G58), .C2(new_n761), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n734), .B1(new_n769), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n732), .A2(new_n734), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n673), .A2(new_n335), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n232), .B2(new_n263), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n248), .B2(G45), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n335), .A2(new_n204), .ZN(new_n786));
  INV_X1    g0586(.A(G355), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n786), .A2(new_n787), .B1(G116), .B2(new_n204), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n781), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n733), .A2(new_n780), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n729), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  INV_X1    g0593(.A(new_n734), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n768), .A2(G159), .B1(new_n761), .B2(G143), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n754), .A2(G137), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(new_n326), .C2(new_n737), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT34), .Z(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G50), .B2(new_n757), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n386), .B1(new_n745), .B2(G132), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n764), .A2(G58), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n773), .A2(G68), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n771), .B1(G311), .B2(new_n745), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n498), .B2(new_n756), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n386), .B1(new_n760), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n773), .A2(G87), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n250), .B2(new_n767), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n805), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n810), .B1(new_n747), .B2(new_n737), .C1(new_n455), .C2(new_n753), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n794), .B1(new_n803), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n734), .A2(new_n730), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n728), .B(new_n812), .C1(new_n306), .C2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT99), .Z(new_n815));
  NAND2_X1  g0615(.A1(new_n641), .A2(new_n655), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n353), .A2(new_n654), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n366), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n818), .B2(new_n641), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n815), .B1(new_n731), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n637), .A2(new_n655), .A3(new_n820), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n819), .B(KEYINPUT100), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n710), .ZN(new_n824));
  INV_X1    g0624(.A(new_n709), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n728), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n821), .A2(new_n827), .ZN(G384));
  NAND2_X1  g0628(.A1(new_n318), .A2(new_n654), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n319), .A2(new_n829), .A3(new_n323), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n292), .A2(new_n318), .A3(new_n654), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n819), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT106), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n704), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n703), .A2(KEYINPUT106), .A3(new_n654), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n705), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(new_n692), .A3(new_n707), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n652), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n436), .A2(KEYINPUT16), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n382), .B1(new_n840), .B2(new_n393), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n443), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n439), .A2(new_n440), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n396), .A2(new_n839), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n410), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n841), .B1(new_n406), .B2(new_n839), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n843), .A3(KEYINPUT37), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n851));
  INV_X1    g0651(.A(KEYINPUT104), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n846), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n845), .B(new_n853), .Z(new_n854));
  AOI21_X1  g0654(.A(new_n844), .B1(new_n442), .B2(new_n640), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n838), .A2(new_n857), .A3(KEYINPUT40), .ZN(new_n858));
  NOR2_X1   g0658(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n842), .A2(new_n847), .A3(new_n849), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n850), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n859), .B1(new_n863), .B2(new_n838), .ZN(new_n864));
  NAND2_X1  g0664(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n858), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT107), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n445), .A2(new_n837), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(G330), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n830), .A2(new_n831), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT102), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n654), .B(new_n819), .C1(new_n630), .C2(new_n636), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n816), .B(KEYINPUT101), .Z(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n822), .A2(KEYINPUT102), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n872), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n863), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n857), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n850), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n319), .A2(new_n654), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n412), .A2(new_n407), .A3(new_n652), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n691), .A2(new_n712), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n445), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n646), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n887), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n870), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n259), .B2(new_n724), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n250), .B1(new_n509), .B2(KEYINPUT35), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n894), .B(new_n229), .C1(KEYINPUT35), .C2(new_n509), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT36), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n233), .B1(new_n222), .B2(new_n389), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n897), .A2(new_n306), .B1(G50), .B2(new_n218), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(G1), .A3(new_n300), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n893), .A2(new_n896), .A3(new_n899), .ZN(G367));
  OAI21_X1  g0700(.A(new_n781), .B1(new_n204), .B2(new_n349), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n242), .B2(new_n782), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT114), .B(G137), .Z(new_n903));
  AOI22_X1  g0703(.A1(G150), .A2(new_n761), .B1(new_n745), .B2(new_n903), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n904), .B1(new_n218), .B2(new_n763), .C1(new_n431), .C2(new_n737), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n330), .A2(new_n767), .B1(new_n749), .B2(new_n306), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n905), .A2(new_n386), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(G143), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n907), .B1(new_n389), .B2(new_n756), .C1(new_n908), .C2(new_n753), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n757), .A2(KEYINPUT46), .A3(G116), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT113), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT46), .B1(new_n757), .B2(G116), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n359), .B2(new_n764), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n279), .A2(new_n749), .B1(new_n767), .B2(new_n747), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n737), .A2(new_n806), .B1(new_n760), .B2(new_n455), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n914), .A2(new_n915), .A3(new_n335), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n911), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(G311), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n917), .B1(new_n918), .B2(new_n753), .C1(new_n739), .C2(new_n744), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT47), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n902), .B1(new_n921), .B2(new_n734), .ZN(new_n922));
  INV_X1    g0722(.A(new_n732), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n554), .A2(new_n555), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n654), .ZN(new_n925));
  MUX2_X1   g0725(.A(new_n631), .B(new_n623), .S(new_n925), .Z(new_n926));
  OAI211_X1 g0726(.A(new_n922), .B(new_n727), .C1(new_n923), .C2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT115), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n618), .A2(new_n654), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n523), .A2(new_n654), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n518), .A2(new_n526), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n668), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT109), .B1(new_n671), .B2(new_n932), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT109), .ZN(new_n937));
  INV_X1    g0737(.A(new_n932), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n616), .A2(new_n937), .A3(new_n938), .A4(new_n670), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n665), .A2(new_n938), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n655), .B1(new_n943), .B2(new_n618), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n936), .A2(KEYINPUT42), .A3(new_n939), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT108), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n947), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n949), .A2(new_n950), .B1(KEYINPUT43), .B2(new_n926), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n946), .A2(new_n948), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT108), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n935), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n676), .B(KEYINPUT41), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n671), .B1(new_n667), .B2(new_n670), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n722), .A2(KEYINPUT112), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT112), .B1(new_n722), .B2(new_n960), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n960), .A2(new_n720), .A3(new_n661), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT111), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n671), .A2(new_n669), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n965), .B1(new_n966), .B2(new_n934), .ZN(new_n967));
  AOI211_X1 g0767(.A(KEYINPUT111), .B(new_n933), .C1(new_n671), .C2(new_n669), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT44), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n967), .B2(new_n968), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n671), .A2(new_n669), .A3(new_n933), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT45), .Z(new_n973));
  NAND3_X1  g0773(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n668), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n668), .A3(new_n973), .A4(new_n971), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n964), .A2(new_n976), .A3(new_n715), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n959), .B1(new_n978), .B2(new_n715), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n958), .B1(new_n979), .B2(new_n726), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n951), .A2(new_n956), .A3(new_n935), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT110), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n951), .A2(new_n956), .A3(KEYINPUT110), .A4(new_n935), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n929), .B1(new_n980), .B2(new_n985), .ZN(G387));
  OR3_X1    g0786(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n987));
  INV_X1    g0787(.A(new_n715), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n676), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n988), .B2(new_n987), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n664), .A2(new_n666), .A3(new_n732), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n678), .A2(new_n786), .B1(G107), .B2(new_n204), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT116), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n328), .A2(G50), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n461), .B1(new_n218), .B2(new_n306), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n996), .A2(new_n677), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n239), .B2(new_n263), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n993), .B1(new_n999), .B2(new_n782), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n781), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n727), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n349), .A2(new_n763), .B1(new_n760), .B2(new_n330), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n347), .B2(new_n738), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G159), .A2(new_n754), .B1(new_n757), .B2(G77), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G68), .A2(new_n768), .B1(new_n773), .B2(G97), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n386), .B1(new_n745), .B2(G150), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n738), .A2(G311), .B1(new_n754), .B2(G322), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n455), .B2(new_n767), .C1(new_n739), .C2(new_n760), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT48), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n747), .B2(new_n763), .C1(new_n806), .C2(new_n756), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT49), .Z(new_n1013));
  INV_X1    g0813(.A(G326), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n386), .B1(new_n744), .B2(new_n1014), .C1(new_n250), .C2(new_n749), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1008), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1002), .B1(new_n1016), .B2(new_n734), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n964), .A2(new_n726), .B1(new_n991), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n990), .A2(new_n1018), .ZN(G393));
  NAND3_X1  g0819(.A1(new_n976), .A2(KEYINPUT118), .A3(new_n977), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(KEYINPUT118), .B2(new_n976), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n987), .A2(new_n988), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n723), .B(new_n978), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n753), .A2(new_n326), .B1(new_n760), .B2(new_n431), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT51), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n808), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n386), .B(new_n1026), .C1(new_n308), .C2(new_n757), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n738), .A2(G50), .B1(new_n764), .B2(G77), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n328), .B2(new_n767), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT119), .Z(new_n1030));
  OAI211_X1 g0830(.A(new_n1027), .B(new_n1030), .C1(new_n908), .C2(new_n744), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n763), .A2(new_n250), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n335), .B1(new_n757), .B2(G283), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n774), .C1(new_n806), .C2(new_n767), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(G322), .C2(new_n745), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n455), .B2(new_n737), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n753), .A2(new_n739), .B1(new_n760), .B2(new_n918), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  OAI21_X1  g0838(.A(new_n1031), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n728), .B1(new_n1039), .B2(new_n734), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n933), .B2(new_n923), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n253), .A2(new_n782), .B1(G97), .B2(new_n673), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n781), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1021), .B2(new_n726), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1023), .A2(new_n1044), .ZN(G390));
  NAND3_X1  g0845(.A1(new_n445), .A2(G330), .A3(new_n837), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n889), .A2(new_n1046), .A3(new_n646), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n832), .A2(new_n837), .A3(G330), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(KEYINPUT120), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n872), .B1(new_n709), .B2(new_n819), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT120), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n832), .A2(new_n837), .A3(new_n1051), .A4(G330), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n876), .A2(new_n878), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n825), .A2(new_n820), .A3(new_n871), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n689), .A2(new_n655), .A3(new_n820), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n877), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n823), .A2(G330), .A3(new_n837), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1056), .B(new_n1059), .C1(new_n871), .C2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1047), .B1(new_n1055), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n882), .A2(new_n883), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n879), .B2(new_n884), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n884), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n857), .B(new_n1066), .C1(new_n1059), .C2(new_n872), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n1065), .A2(new_n1067), .A3(new_n1056), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1063), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1065), .A2(new_n1067), .A3(new_n1056), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n857), .A2(new_n1066), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n871), .B2(new_n1058), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n874), .A2(new_n873), .A3(new_n875), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT102), .B1(new_n822), .B2(new_n877), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n871), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1066), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1078), .B2(new_n1064), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1072), .B(new_n1062), .C1(new_n1079), .C2(new_n1069), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1071), .A2(new_n723), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT121), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1071), .A2(KEYINPUT121), .A3(new_n1080), .A4(new_n723), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1072), .B(new_n726), .C1(new_n1079), .C2(new_n1069), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1064), .A2(new_n730), .ZN(new_n1087));
  INV_X1    g0887(.A(G125), .ZN(new_n1088));
  INV_X1    g0888(.A(G132), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n335), .B1(new_n744), .B2(new_n1088), .C1(new_n1089), .C2(new_n760), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n757), .A2(G150), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT53), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(G159), .C2(new_n764), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n738), .A2(new_n903), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT54), .B(G143), .Z(new_n1095));
  NAND2_X1  g0895(.A1(new_n768), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n754), .A2(G128), .B1(new_n773), .B2(G50), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n802), .B1(new_n306), .B2(new_n763), .C1(new_n531), .C2(new_n756), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n386), .B1(new_n737), .B2(new_n358), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n767), .A2(new_n279), .B1(new_n744), .B2(new_n806), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n250), .B2(new_n760), .C1(new_n747), .C2(new_n753), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n794), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n728), .B(new_n1104), .C1(new_n328), .C2(new_n813), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1087), .A2(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1086), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1085), .A2(new_n1107), .ZN(G378));
  INV_X1    g0908(.A(KEYINPUT57), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1047), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1080), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n645), .A2(new_n343), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n334), .A2(new_n839), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1113), .B(new_n1116), .Z(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n866), .B2(G330), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n850), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n849), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n841), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n414), .B2(new_n442), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n1122), .B2(new_n839), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT38), .B1(new_n1123), .B2(new_n847), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n838), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n859), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n865), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n838), .A2(new_n857), .A3(KEYINPUT40), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1127), .A2(G330), .A3(new_n1128), .A4(new_n1117), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1112), .B1(new_n1118), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1127), .A2(G330), .A3(new_n1128), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1117), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n887), .A3(new_n1129), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1109), .B1(new_n1111), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1134), .A2(new_n887), .A3(new_n1129), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n887), .B1(new_n1134), .B2(new_n1129), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1080), .A2(new_n1110), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(KEYINPUT57), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1142), .A3(new_n723), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n728), .B1(new_n330), .B2(new_n813), .ZN(new_n1144));
  AOI21_X1  g0944(.A(G50), .B1(new_n266), .B2(new_n420), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n306), .A2(new_n756), .B1(new_n760), .B2(new_n498), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n1146), .C1(G68), .C2(new_n764), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n335), .B1(new_n773), .B2(G58), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n768), .A2(new_n538), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G97), .A2(new_n738), .B1(new_n745), .B2(G283), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G116), .B2(new_n754), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT58), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT122), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(G124), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(G124), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n745), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n768), .A2(G137), .B1(new_n761), .B2(G128), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n757), .A2(new_n1095), .B1(new_n764), .B2(G150), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n1088), .B2(new_n753), .C1(new_n1089), .C2(new_n737), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n420), .B(new_n1157), .C1(new_n1161), .C2(KEYINPUT59), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G33), .B(new_n1162), .C1(G159), .C2(new_n773), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(KEYINPUT59), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1145), .B(new_n1153), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1144), .B1(new_n794), .B2(new_n1165), .C1(new_n1133), .C2(new_n731), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1140), .B2(new_n726), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1143), .A2(new_n1168), .ZN(G375));
  INV_X1    g0969(.A(new_n959), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1055), .A2(new_n1047), .A3(new_n1061), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1063), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n725), .B1(new_n1055), .B2(new_n1061), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n872), .A2(new_n730), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n349), .A2(new_n763), .B1(new_n744), .B2(new_n455), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n749), .A2(new_n306), .B1(new_n756), .B2(new_n279), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n386), .B1(new_n767), .B2(new_n358), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n753), .A2(new_n806), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n250), .B2(new_n737), .C1(new_n747), .C2(new_n760), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n763), .A2(new_n330), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n753), .A2(new_n1089), .B1(new_n749), .B2(new_n389), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n761), .C2(new_n903), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n738), .A2(new_n1095), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n745), .A2(G128), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n335), .B1(new_n767), .B2(new_n326), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G159), .B2(new_n757), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n794), .B1(new_n1180), .B2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n728), .B(new_n1189), .C1(new_n218), .C2(new_n813), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1173), .B1(new_n1174), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1172), .A2(new_n1191), .ZN(G381));
  AND3_X1   g0992(.A1(new_n1081), .A2(new_n1107), .A3(KEYINPUT123), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT123), .B1(new_n1081), .B2(new_n1107), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1195), .A2(new_n1168), .A3(new_n1143), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n1191), .A3(new_n1172), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n990), .A2(new_n792), .A3(new_n1018), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(G387), .A2(G390), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1197), .A2(G384), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT124), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1203), .A2(new_n1204), .ZN(G407));
  NAND2_X1  g1005(.A1(new_n1196), .A2(new_n653), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G213), .B(new_n1206), .C1(new_n1203), .C2(new_n1204), .ZN(G409));
  INV_X1    g1007(.A(KEYINPUT127), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n976), .A2(new_n977), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n715), .B1(new_n1209), .B2(new_n987), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1170), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n957), .B1(new_n1211), .B2(new_n725), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n983), .A2(new_n984), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n928), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT126), .B1(new_n1214), .B2(G390), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1198), .ZN(new_n1217));
  INV_X1    g1017(.A(G390), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(G387), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G390), .B(new_n929), .C1(new_n980), .C2(new_n985), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1215), .A2(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .A4(new_n1217), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1140), .A2(new_n1170), .A3(new_n1141), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1168), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1107), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(G375), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G213), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(G343), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n676), .B1(new_n1171), .B2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1055), .A2(new_n1047), .A3(new_n1061), .A4(KEYINPUT60), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1063), .A3(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(G384), .A3(new_n1191), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G384), .B1(new_n1239), .B2(new_n1191), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1232), .A2(new_n1235), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT125), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1242), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1240), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1234), .A2(G2897), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1246), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1243), .A2(new_n1248), .A3(G2897), .A4(new_n1234), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1244), .A2(KEYINPUT62), .B1(new_n1245), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1243), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G378), .A2(new_n1168), .A3(new_n1143), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1234), .B(new_n1255), .C1(new_n1256), .C2(new_n1229), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT61), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1226), .B1(new_n1254), .B2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1232), .A2(KEYINPUT63), .A3(new_n1235), .A4(new_n1243), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1217), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1222), .B1(G387), .B2(new_n1218), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1265), .B2(new_n1223), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1234), .B1(new_n1256), .B2(new_n1229), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT63), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1267), .B1(new_n1244), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1208), .B1(new_n1260), .B2(new_n1271), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1257), .A2(new_n1258), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1244), .B2(KEYINPUT62), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1225), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1270), .A2(new_n1244), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1266), .A3(new_n1261), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1278), .A3(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1272), .A2(new_n1279), .ZN(G405));
  INV_X1    g1080(.A(new_n1256), .ZN(new_n1281));
  AND2_X1   g1081(.A1(G375), .A2(new_n1195), .ZN(new_n1282));
  OR3_X1    g1082(.A1(new_n1225), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1225), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1243), .ZN(G402));
endmodule


