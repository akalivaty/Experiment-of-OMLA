//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1239,
    new_n1240, new_n1241, new_n1242;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  OR3_X1    g0007(.A1(KEYINPUT65), .A2(G58), .A3(G68), .ZN(new_n208));
  OAI21_X1  g0008(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n208), .A2(G50), .A3(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n213), .ZN(new_n217));
  INV_X1    g0017(.A(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT64), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT0), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n215), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(new_n223), .B2(new_n222), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT1), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AND2_X1   g0028(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n227), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n233));
  INV_X1    g0033(.A(G58), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  INV_X1    g0035(.A(G257), .ZN(new_n236));
  OAI221_X1 g0036(.A(new_n233), .B1(new_n234), .B2(new_n235), .C1(new_n204), .C2(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(new_n231), .B2(KEYINPUT67), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n217), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g0039(.A(new_n225), .B1(new_n226), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g0040(.A(new_n240), .B1(new_n226), .B2(new_n239), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(KEYINPUT68), .Z(G361));
  XOR2_X1   g0042(.A(G226), .B(G232), .Z(new_n243));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G250), .B(G257), .Z(new_n248));
  XNOR2_X1  g0048(.A(G264), .B(G270), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G358));
  XOR2_X1   g0051(.A(G97), .B(G107), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G50), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G68), .ZN(new_n256));
  INV_X1    g0056(.A(G68), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G50), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(G58), .B(G77), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n254), .B(new_n261), .ZN(G351));
  NAND2_X1  g0062(.A1(new_n217), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n212), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n216), .B2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G77), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n216), .A2(G13), .A3(G20), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(G77), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT74), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n213), .A2(new_n271), .A3(KEYINPUT73), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT73), .B1(new_n213), .B2(new_n271), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n213), .A2(G33), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT15), .B(G87), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n276), .B1(new_n213), .B2(new_n202), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n268), .B1(new_n279), .B2(new_n264), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G107), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G238), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n286), .B1(new_n288), .B2(new_n289), .C1(new_n235), .C2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT70), .B1(G33), .B2(G41), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(new_n212), .ZN(new_n300));
  NAND3_X1  g0100(.A1(KEYINPUT70), .A2(G33), .A3(G41), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G244), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n294), .A2(new_n298), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n280), .B1(new_n281), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n294), .A2(new_n309), .A3(new_n298), .A4(new_n306), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT75), .B(G200), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n280), .B(new_n315), .C1(new_n316), .C2(new_n307), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT77), .ZN(new_n319));
  INV_X1    g0119(.A(new_n293), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n285), .A2(new_n290), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(G223), .B1(G77), .B2(new_n285), .ZN(new_n322));
  INV_X1    g0122(.A(G222), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n291), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n325), .B2(new_n324), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n297), .B1(new_n305), .B2(G226), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n314), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n265), .A2(G50), .ZN(new_n331));
  INV_X1    g0131(.A(G150), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n274), .A2(new_n332), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n269), .A2(new_n277), .B1(new_n213), .B2(new_n201), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n264), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n331), .B(new_n335), .C1(G50), .C2(new_n267), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT9), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n329), .A2(new_n316), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT10), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n339), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n330), .A4(new_n337), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n329), .A2(new_n281), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n336), .C1(G179), .C2(new_n329), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n274), .A2(new_n255), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n277), .A2(new_n202), .B1(new_n213), .B2(G68), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n264), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT78), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT78), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n264), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(KEYINPUT11), .A3(new_n353), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n267), .A2(G68), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT12), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n265), .B2(G68), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT79), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n356), .A2(KEYINPUT79), .A3(new_n357), .A4(new_n360), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G97), .ZN(new_n366));
  INV_X1    g0166(.A(G226), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n288), .B2(new_n235), .C1(new_n367), .C2(new_n291), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n293), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT13), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n297), .B1(new_n305), .B2(G238), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g0174(.A(G169), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT14), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n377), .B(G169), .C1(new_n373), .C2(new_n374), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n373), .A2(new_n374), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G179), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n365), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n363), .A2(new_n364), .ZN(new_n383));
  INV_X1    g0183(.A(G200), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n369), .A2(new_n371), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT13), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n384), .B1(new_n386), .B2(new_n372), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(G190), .B2(new_n379), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT80), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n383), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n383), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n382), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n285), .A2(G1698), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT82), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n321), .A2(new_n395), .A3(G226), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT82), .B1(new_n288), .B2(new_n367), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n293), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n297), .B1(new_n305), .B2(G232), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G169), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(G179), .A3(new_n400), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(G58), .B(G68), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n275), .A2(G159), .B1(G20), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n285), .A2(new_n213), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT7), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n406), .B1(new_n408), .B2(new_n257), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT16), .B(new_n406), .C1(new_n408), .C2(new_n257), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n264), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n269), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n267), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n265), .B2(new_n414), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(KEYINPUT81), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT81), .B1(new_n413), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n404), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n413), .A2(new_n416), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT81), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n417), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n404), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n401), .A2(G200), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n399), .A2(G190), .A3(new_n400), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n413), .A2(new_n428), .A3(new_n416), .A4(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n421), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  NOR4_X1   g0234(.A1(new_n319), .A2(new_n347), .A3(new_n392), .A4(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n282), .A2(new_n284), .A3(G250), .A4(new_n290), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n282), .A2(new_n284), .A3(G257), .A4(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G294), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n293), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n216), .A2(G45), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G41), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(KEYINPUT5), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n446), .A2(new_n296), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n302), .A2(new_n446), .A3(G264), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n440), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n384), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n440), .A2(new_n447), .A3(new_n316), .A4(new_n448), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G116), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G20), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT88), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n455), .A2(new_n456), .B1(new_n205), .B2(G20), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n455), .B2(new_n456), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n205), .A2(KEYINPUT88), .A3(KEYINPUT23), .A4(G20), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n282), .A2(new_n284), .A3(new_n213), .A4(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT22), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n287), .A2(new_n463), .A3(new_n213), .A4(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n460), .A2(new_n465), .A3(KEYINPUT24), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n264), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n267), .A2(G107), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT89), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT25), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(KEYINPUT25), .B2(new_n471), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(KEYINPUT25), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(KEYINPUT89), .B2(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n217), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n216), .A2(G33), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n477), .A2(new_n267), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n479), .A2(G107), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n452), .A2(new_n470), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n470), .A2(new_n481), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n449), .A2(G169), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT90), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT91), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n449), .B2(new_n309), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n302), .A2(new_n446), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n488), .A2(G264), .B1(new_n439), .B2(new_n293), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(KEYINPUT91), .A3(G179), .A4(new_n447), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT90), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n449), .A2(new_n491), .A3(G169), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n485), .A2(new_n487), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n482), .B1(new_n483), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n278), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n479), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n287), .A2(new_n213), .A3(G68), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n213), .B1(new_n366), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G87), .B2(new_n206), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n277), .B2(new_n204), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI22_X1  g0302(.A1(new_n502), .A2(new_n477), .B1(new_n267), .B2(new_n495), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n503), .A2(KEYINPUT86), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(KEYINPUT86), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n496), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G244), .ZN(new_n507));
  OAI221_X1 g0307(.A(new_n453), .B1(new_n288), .B2(new_n507), .C1(new_n289), .C2(new_n291), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n293), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n441), .A2(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n441), .A2(KEYINPUT85), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n510), .A2(G250), .A3(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(new_n302), .B1(G274), .B2(new_n442), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n309), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n281), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n506), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(G190), .A3(new_n513), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT87), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n503), .B(KEYINPUT86), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n514), .A2(new_n314), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n479), .A2(G87), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n518), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n408), .A2(new_n205), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n205), .A2(G97), .ZN(new_n529));
  XNOR2_X1  g0329(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n530));
  MUX2_X1   g0330(.A(new_n529), .B(new_n252), .S(new_n530), .Z(new_n531));
  OAI22_X1  g0331(.A1(new_n531), .A2(new_n213), .B1(new_n202), .B2(new_n274), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n264), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n267), .A2(G97), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n479), .B2(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n302), .A2(new_n446), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n447), .B1(new_n538), .B2(new_n236), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n393), .A2(KEYINPUT4), .A3(G244), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT4), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n291), .B2(new_n507), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n321), .A2(G250), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n540), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n539), .B1(new_n545), .B2(new_n293), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G190), .ZN(new_n547));
  INV_X1    g0347(.A(new_n546), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  OAI21_X1  g0350(.A(G200), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n537), .B(new_n547), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n281), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n546), .A2(new_n309), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n536), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n479), .A2(G116), .ZN(new_n557));
  INV_X1    g0357(.A(G116), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n263), .A2(new_n212), .B1(G20), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n543), .B(new_n213), .C1(G33), .C2(new_n204), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT20), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  OAI221_X1 g0362(.A(new_n557), .B1(G116), .B2(new_n267), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n488), .A2(G270), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n285), .A2(G303), .ZN(new_n565));
  INV_X1    g0365(.A(G264), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n288), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(G257), .B2(new_n393), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n447), .B(new_n564), .C1(new_n568), .C2(new_n320), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n563), .B1(new_n569), .B2(G200), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n316), .B2(new_n569), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n563), .A2(new_n569), .A3(G169), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n563), .A2(new_n569), .A3(KEYINPUT21), .A4(G169), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n569), .A2(new_n309), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n563), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n571), .A2(new_n574), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n556), .A2(new_n578), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n435), .A2(new_n494), .A3(new_n527), .A4(new_n579), .ZN(G372));
  INV_X1    g0380(.A(new_n433), .ZN(new_n581));
  INV_X1    g0381(.A(new_n313), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n390), .B2(new_n391), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n583), .B2(new_n382), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n413), .A2(new_n416), .B1(new_n402), .B2(new_n403), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n585), .B(new_n426), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n344), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(new_n346), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT26), .B1(new_n526), .B2(new_n555), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT92), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n517), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT92), .B1(new_n514), .B2(new_n281), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n516), .B(new_n506), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n555), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n522), .A2(new_n523), .A3(new_n524), .A4(new_n519), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n589), .B1(new_n596), .B2(KEYINPUT26), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n452), .A2(new_n470), .A3(new_n481), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n552), .A2(new_n598), .A3(new_n555), .A4(new_n595), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n574), .A2(new_n577), .A3(new_n575), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n493), .A2(new_n483), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n593), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n435), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n588), .A2(new_n606), .ZN(G369));
  NOR2_X1   g0407(.A1(new_n218), .A2(G20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n216), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n609), .A2(KEYINPUT27), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(KEYINPUT27), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(G213), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(G343), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n563), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n578), .B2(KEYINPUT93), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(KEYINPUT93), .B2(new_n578), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n600), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G330), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT95), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n483), .A2(new_n614), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n601), .A2(new_n598), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT94), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT94), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n601), .A2(new_n598), .A3(new_n625), .A4(new_n622), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n614), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n601), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n621), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  AOI211_X1 g0431(.A(KEYINPUT95), .B(new_n629), .C1(new_n624), .C2(new_n626), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n620), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n601), .A2(new_n614), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n627), .A2(new_n630), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT95), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n627), .A2(new_n621), .A3(new_n630), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n600), .A2(new_n628), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n636), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n635), .A2(new_n643), .ZN(G399));
  NAND3_X1  g0444(.A1(new_n220), .A2(KEYINPUT96), .A3(new_n443), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT96), .B1(new_n220), .B2(new_n443), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G1), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n210), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT28), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT29), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n599), .A2(new_n603), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n526), .A2(KEYINPUT26), .A3(new_n555), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n596), .A2(KEYINPUT26), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .A4(new_n593), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n654), .B1(new_n658), .B2(new_n628), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(KEYINPUT98), .A2(KEYINPUT30), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n515), .A2(new_n489), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT98), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT30), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n663), .A2(new_n546), .A3(new_n576), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n576), .A2(new_n546), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n515), .A2(new_n489), .A3(new_n662), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n668), .A2(new_n669), .B1(new_n664), .B2(new_n665), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n569), .A2(new_n514), .A3(new_n309), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(KEYINPUT97), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n449), .B(new_n548), .C1(new_n671), .C2(KEYINPUT97), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n667), .B(new_n670), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT31), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n674), .A2(new_n675), .A3(new_n614), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n579), .A2(new_n494), .A3(new_n527), .A4(new_n628), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n675), .B1(new_n674), .B2(new_n614), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n654), .B(new_n628), .C1(new_n597), .C2(new_n604), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n660), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n653), .B1(new_n683), .B2(G1), .ZN(G364));
  AOI21_X1  g0484(.A(new_n216), .B1(new_n608), .B2(G45), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n649), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n219), .A2(new_n285), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n687), .A2(G355), .B1(new_n558), .B2(new_n219), .ZN(new_n688));
  INV_X1    g0488(.A(G45), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n261), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n219), .A2(new_n287), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(G45), .B2(new_n210), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(G13), .A2(G33), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G20), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n212), .B1(G20), .B2(new_n281), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n686), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n697), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n213), .A2(G190), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n309), .A3(new_n384), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT99), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT99), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  XOR2_X1   g0506(.A(KEYINPUT100), .B(G159), .Z(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT32), .ZN(new_n709));
  INV_X1    g0509(.A(new_n314), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n213), .A2(new_n316), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n710), .A2(G179), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n713), .A2(G87), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n309), .A2(new_n384), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n309), .A2(G200), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n701), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n717), .A2(G50), .B1(new_n720), .B2(G77), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n711), .A2(new_n718), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n234), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n715), .A2(new_n701), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n316), .A2(G179), .A3(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n213), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n287), .B1(new_n724), .B2(new_n257), .C1(new_n726), .C2(new_n204), .ZN(new_n727));
  NOR4_X1   g0527(.A1(new_n709), .A2(new_n714), .A3(new_n723), .A4(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n701), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n710), .A2(G179), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT101), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G107), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n706), .A2(G329), .ZN(new_n734));
  INV_X1    g0534(.A(new_n726), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G294), .ZN(new_n736));
  INV_X1    g0536(.A(new_n724), .ZN(new_n737));
  XNOR2_X1  g0537(.A(KEYINPUT33), .B(G317), .ZN(new_n738));
  AOI22_X1  g0538(.A1(G326), .A2(new_n717), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n722), .ZN(new_n740));
  AOI22_X1  g0540(.A1(G322), .A2(new_n740), .B1(new_n720), .B2(G311), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n734), .A2(new_n736), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(G283), .B2(new_n732), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n287), .B1(new_n713), .B2(G303), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT102), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n728), .A2(new_n733), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n696), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n699), .B1(new_n700), .B2(new_n746), .C1(new_n619), .C2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n620), .ZN(new_n749));
  INV_X1    g0549(.A(new_n686), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n619), .A2(G330), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(G396));
  NAND2_X1  g0554(.A1(new_n605), .A2(new_n628), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n308), .A2(new_n312), .A3(new_n614), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT103), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n308), .A2(new_n312), .A3(KEYINPUT103), .A4(new_n614), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n313), .B(new_n317), .C1(new_n280), .C2(new_n628), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n755), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n762), .B(new_n628), .C1(new_n597), .C2(new_n604), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n680), .ZN(new_n767));
  INV_X1    g0567(.A(new_n680), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(new_n764), .A3(new_n765), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n750), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n763), .A2(new_n694), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n717), .A2(G137), .B1(new_n720), .B2(new_n707), .ZN(new_n772));
  INV_X1    g0572(.A(G143), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n772), .B1(new_n773), .B2(new_n722), .C1(new_n332), .C2(new_n724), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT34), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n732), .A2(G68), .ZN(new_n776));
  INV_X1    g0576(.A(G132), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n287), .B1(new_n234), .B2(new_n726), .C1(new_n705), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(G50), .B2(new_n713), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n732), .A2(G87), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n724), .A2(new_n782), .B1(new_n719), .B2(new_n558), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n285), .B1(new_n716), .B2(new_n784), .C1(new_n726), .C2(new_n204), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(G294), .C2(new_n740), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n706), .A2(G311), .B1(G107), .B2(new_n713), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n781), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n700), .B1(new_n780), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n697), .A2(new_n694), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n202), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n686), .B1(new_n771), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n770), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT104), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n770), .A2(KEYINPUT104), .A3(new_n792), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G384));
  INV_X1    g0598(.A(KEYINPUT35), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n531), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n531), .A2(new_n799), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n800), .A2(new_n801), .A3(G116), .A4(new_n214), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT36), .Z(new_n803));
  OAI211_X1 g0603(.A(new_n211), .B(G77), .C1(new_n234), .C2(new_n257), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n216), .B(G13), .C1(new_n804), .C2(new_n256), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT38), .ZN(new_n807));
  INV_X1    g0607(.A(new_n612), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n422), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n420), .A2(KEYINPUT18), .B1(new_n431), .B2(new_n432), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(new_n427), .ZN(new_n811));
  INV_X1    g0611(.A(new_n430), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT106), .B1(new_n812), .B2(new_n585), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n422), .A2(new_n404), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT106), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n815), .A3(new_n430), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n809), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT37), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n430), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n425), .B2(new_n404), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n425), .A2(new_n808), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n817), .A2(KEYINPUT37), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n807), .B1(new_n811), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n817), .A2(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n820), .A2(new_n821), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n809), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n434), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n826), .A2(new_n828), .A3(KEYINPUT38), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT107), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n375), .A2(KEYINPUT14), .B1(new_n379), .B2(G179), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n383), .B1(new_n832), .B2(new_n378), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT105), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT105), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n382), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n383), .A2(new_n628), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n383), .A2(new_n388), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT80), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n383), .A2(new_n388), .A3(new_n389), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n392), .A2(new_n838), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n845), .A2(new_n679), .A3(new_n762), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT107), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n823), .A2(new_n829), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n831), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT40), .ZN(new_n850));
  INV_X1    g0650(.A(new_n825), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n812), .A2(new_n585), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n818), .B1(new_n821), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n581), .A2(new_n586), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n851), .A2(new_n853), .B1(new_n854), .B2(new_n821), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n807), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n850), .B1(new_n856), .B2(new_n829), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n849), .A2(new_n850), .B1(new_n846), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n435), .A3(new_n679), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n846), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n823), .A2(new_n829), .A3(new_n847), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n847), .B1(new_n823), .B2(new_n829), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n845), .A2(new_n679), .A3(new_n762), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(G330), .B(new_n860), .C1(new_n864), .C2(KEYINPUT40), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n435), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n680), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n859), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n681), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n435), .B1(new_n659), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n588), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n869), .B(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n856), .A2(new_n874), .A3(new_n829), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n837), .A2(new_n614), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n586), .A2(new_n612), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n582), .A2(new_n628), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n765), .A2(new_n881), .B1(new_n843), .B2(new_n844), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n831), .A2(new_n882), .A3(new_n848), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n873), .A2(new_n884), .B1(new_n216), .B2(new_n608), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n873), .A2(new_n884), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n806), .B1(new_n885), .B2(new_n886), .ZN(G367));
  NAND2_X1  g0687(.A1(new_n522), .A2(new_n524), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n614), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n593), .A2(new_n595), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n593), .B2(new_n889), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n891), .A2(new_n747), .ZN(new_n892));
  INV_X1    g0692(.A(new_n691), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n698), .B1(new_n220), .B2(new_n278), .C1(new_n250), .C2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT112), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n686), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  INV_X1    g0697(.A(G311), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n716), .A2(new_n898), .B1(new_n722), .B2(new_n784), .ZN(new_n899));
  OAI221_X1 g0699(.A(new_n285), .B1(new_n719), .B2(new_n782), .C1(new_n726), .C2(new_n205), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n899), .B(new_n900), .C1(G294), .C2(new_n737), .ZN(new_n901));
  INV_X1    g0701(.A(new_n730), .ZN(new_n902));
  INV_X1    g0702(.A(G317), .ZN(new_n903));
  OAI221_X1 g0703(.A(new_n901), .B1(new_n204), .B2(new_n902), .C1(new_n903), .C2(new_n705), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n713), .A2(G116), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT46), .Z(new_n906));
  INV_X1    g0706(.A(new_n707), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n907), .A2(new_n724), .B1(new_n719), .B2(new_n255), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n706), .A2(G137), .B1(KEYINPUT113), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n713), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n909), .B1(new_n234), .B2(new_n910), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n287), .B1(new_n722), .B2(new_n332), .C1(new_n773), .C2(new_n716), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(G68), .B2(new_n735), .ZN(new_n913));
  OAI221_X1 g0713(.A(new_n913), .B1(KEYINPUT113), .B2(new_n908), .C1(new_n202), .C2(new_n902), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n904), .A2(new_n906), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT47), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n700), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n897), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n892), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT111), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n642), .B1(new_n631), .B2(new_n632), .ZN(new_n922));
  INV_X1    g0722(.A(new_n636), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n552), .B(new_n555), .C1(new_n537), .C2(new_n628), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n594), .A2(new_n614), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT45), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n922), .A2(new_n923), .ZN(new_n931));
  INV_X1    g0731(.A(new_n926), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT44), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT44), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n934), .B(new_n926), .C1(new_n922), .C2(new_n923), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n929), .A2(new_n930), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n634), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n643), .B2(new_n926), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(KEYINPUT44), .A3(new_n932), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n927), .B(new_n928), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n941), .A3(new_n635), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n633), .A2(new_n641), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n749), .A2(new_n922), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n749), .B1(new_n943), .B2(new_n922), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n682), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n937), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n947), .A2(new_n683), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n648), .B(KEYINPUT41), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT109), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n947), .B2(new_n683), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT109), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n685), .B(KEYINPUT110), .Z(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n891), .A2(KEYINPUT43), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n640), .A2(new_n642), .A3(new_n926), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT108), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT42), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n594), .B1(new_n552), .B2(new_n602), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n960), .A2(new_n961), .B1(new_n614), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n960), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n634), .A2(new_n926), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n891), .A2(KEYINPUT43), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n966), .B(new_n967), .Z(new_n968));
  XNOR2_X1  g0768(.A(new_n965), .B(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n921), .B1(new_n957), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n956), .B1(new_n952), .B2(new_n953), .ZN(new_n971));
  AOI211_X1 g0771(.A(KEYINPUT109), .B(new_n950), .C1(new_n947), .C2(new_n683), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n969), .B(new_n921), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n920), .B1(new_n970), .B2(new_n974), .ZN(G387));
  INV_X1    g0775(.A(KEYINPUT114), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n946), .B2(new_n649), .ZN(new_n977));
  INV_X1    g0777(.A(new_n946), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(KEYINPUT114), .A3(new_n648), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n944), .A2(new_n945), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n977), .B(new_n979), .C1(new_n683), .C2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n633), .A2(new_n696), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n287), .B1(new_n706), .B2(G326), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n558), .B2(new_n902), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n717), .A2(G322), .B1(new_n720), .B2(G303), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n898), .B2(new_n724), .C1(new_n903), .C2(new_n722), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT48), .Z(new_n987));
  INV_X1    g0787(.A(G294), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n910), .A2(new_n988), .B1(new_n726), .B2(new_n782), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT49), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n984), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n992), .B2(new_n991), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n722), .A2(new_n255), .B1(new_n719), .B2(new_n257), .ZN(new_n995));
  INV_X1    g0795(.A(G159), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n287), .B1(new_n716), .B2(new_n996), .C1(new_n726), .C2(new_n278), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n995), .B(new_n997), .C1(new_n414), .C2(new_n737), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n706), .A2(G150), .B1(G77), .B2(new_n713), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n204), .C2(new_n731), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n700), .B1(new_n994), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n247), .A2(new_n689), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n650), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1002), .A2(new_n691), .B1(new_n1003), .B2(new_n687), .ZN(new_n1004));
  AOI21_X1  g0804(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n270), .A2(new_n255), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n650), .B(new_n1005), .C1(new_n1006), .C2(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(KEYINPUT50), .B2(new_n1006), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1004), .A2(new_n1008), .B1(G107), .B2(new_n220), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n686), .B(new_n1001), .C1(new_n698), .C2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n980), .A2(new_n955), .B1(new_n982), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n981), .A2(new_n1011), .ZN(G393));
  INV_X1    g0812(.A(new_n937), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n942), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n978), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n648), .A3(new_n947), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n937), .A2(new_n942), .A3(new_n955), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n698), .B1(new_n204), .B2(new_n220), .C1(new_n254), .C2(new_n893), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n750), .A2(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n287), .B1(new_n724), .B2(new_n255), .C1(new_n726), .C2(new_n202), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n706), .B2(G143), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n716), .A2(new_n332), .B1(new_n722), .B2(new_n996), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT51), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n270), .A2(new_n720), .B1(new_n713), .B2(G68), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n781), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n287), .B1(new_n706), .B2(G322), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n733), .B(new_n1026), .C1(new_n782), .C2(new_n910), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT116), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n716), .A2(new_n903), .B1(new_n722), .B2(new_n898), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1029), .B(new_n1030), .Z(new_n1031));
  AOI22_X1  g0831(.A1(G303), .A2(new_n737), .B1(new_n720), .B2(G294), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n558), .C2(new_n726), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1025), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1019), .B1(new_n1034), .B2(new_n697), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n926), .B2(new_n747), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1016), .A2(new_n1017), .A3(new_n1036), .ZN(G390));
  INV_X1    g0837(.A(KEYINPUT119), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n677), .A2(new_n678), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n676), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1039), .A2(G330), .A3(new_n1040), .A4(new_n762), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n837), .A2(new_n842), .B1(new_n392), .B2(new_n838), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1038), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n658), .A2(new_n628), .A3(new_n762), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n881), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(KEYINPUT119), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n765), .A2(new_n881), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n588), .B(new_n871), .C1(new_n867), .C2(new_n680), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT118), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n882), .B2(new_n878), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1051), .A2(new_n845), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n878), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1059), .A2(KEYINPUT118), .A3(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1061), .A3(new_n876), .A4(new_n875), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1044), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1047), .A2(new_n845), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n878), .B(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n856), .A2(new_n829), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n1062), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1056), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n1044), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1054), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1062), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1070), .A2(new_n648), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n875), .A2(new_n876), .A3(new_n694), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G283), .A2(new_n717), .B1(new_n737), .B2(G107), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n558), .B2(new_n722), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n285), .B1(new_n719), .B2(new_n204), .C1(new_n726), .C2(new_n202), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n776), .B1(new_n988), .B2(new_n705), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n714), .B(new_n1082), .C1(new_n1083), .C2(KEYINPUT120), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(KEYINPUT120), .B2(new_n1083), .ZN(new_n1085));
  INV_X1    g0885(.A(G128), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n716), .A2(new_n1086), .B1(new_n722), .B2(new_n777), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n285), .B1(new_n737), .B2(G137), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n996), .B2(new_n726), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT54), .B(G143), .Z(new_n1090));
  AOI211_X1 g0890(.A(new_n1087), .B(new_n1089), .C1(new_n720), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n713), .A2(G150), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT53), .Z(new_n1093));
  AOI22_X1  g0893(.A1(new_n706), .A2(G125), .B1(G50), .B2(new_n730), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n700), .B1(new_n1085), .B2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n686), .B(new_n1096), .C1(new_n269), .C2(new_n790), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1077), .A2(new_n955), .B1(new_n1078), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1076), .A2(new_n1098), .ZN(G378));
  NAND2_X1  g0899(.A1(new_n336), .A2(new_n808), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n347), .B(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1101), .B(new_n1102), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n865), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1103), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n858), .A2(G330), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n884), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n955), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n686), .B1(new_n255), .B2(new_n790), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n271), .B(new_n443), .C1(new_n902), .C2(new_n907), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G124), .B2(new_n706), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n713), .A2(new_n1090), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G125), .A2(new_n717), .B1(new_n737), .B2(G132), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G128), .A2(new_n740), .B1(new_n720), .B2(G137), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n735), .A2(G150), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1119));
  OR2_X1    g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1113), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n730), .A2(G58), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n910), .B2(new_n202), .C1(new_n782), .C2(new_n705), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G97), .A2(new_n737), .B1(new_n740), .B2(G107), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n278), .B2(new_n719), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n287), .A2(G41), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n716), .B2(new_n558), .C1(new_n257), .C2(new_n726), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1129), .A2(KEYINPUT58), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(KEYINPUT58), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1127), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1132), .B(new_n255), .C1(G33), .C2(G41), .ZN(new_n1133));
  AND4_X1   g0933(.A1(new_n1122), .A2(new_n1130), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1111), .B1(new_n700), .B2(new_n1134), .C1(new_n1105), .C2(new_n695), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1110), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n865), .A2(new_n1103), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1105), .B1(new_n858), .B2(G330), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n884), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1140), .A2(new_n1141), .B1(new_n1055), .B2(new_n1075), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n648), .B1(new_n1142), .B2(KEYINPUT57), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1075), .A2(new_n1055), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1137), .B1(new_n1143), .B2(new_n1147), .ZN(G375));
  NAND3_X1  g0948(.A1(new_n1050), .A2(new_n1054), .A3(new_n1052), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1056), .A2(new_n949), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1042), .A2(KEYINPUT122), .A3(new_n694), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT122), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n845), .B2(new_n695), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n285), .B1(new_n722), .B2(new_n782), .C1(new_n726), .C2(new_n278), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n719), .A2(new_n205), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n716), .A2(new_n988), .B1(new_n724), .B2(new_n558), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n204), .B2(new_n910), .C1(new_n784), .C2(new_n705), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n731), .A2(new_n202), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G132), .A2(new_n717), .B1(new_n740), .B2(G137), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n720), .A2(G150), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n735), .A2(G50), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n285), .B1(new_n737), .B2(new_n1090), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1123), .B1(new_n910), .B2(new_n996), .C1(new_n1086), .C2(new_n705), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n1158), .A2(new_n1159), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n697), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n686), .B1(new_n257), .B2(new_n790), .ZN(new_n1168));
  AND4_X1   g0968(.A1(new_n1151), .A2(new_n1153), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1053), .B2(new_n955), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1150), .A2(new_n1170), .ZN(G381));
  OR2_X1    g0971(.A1(G393), .A2(G396), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(G384), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT123), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n920), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT111), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1177), .B2(new_n973), .ZN(new_n1178));
  INV_X1    g0978(.A(G390), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n649), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1142), .A2(KEYINPUT57), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1136), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(G378), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OR4_X1    g0985(.A1(G381), .A2(new_n1174), .A3(new_n1180), .A4(new_n1185), .ZN(G407));
  OAI211_X1 g0986(.A(G407), .B(G213), .C1(G343), .C2(new_n1185), .ZN(G409));
  NAND2_X1  g0987(.A1(G387), .A2(G390), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(G393), .B(G396), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1180), .A2(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT126), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1190), .B1(new_n1178), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1175), .B(G390), .C1(new_n1177), .C2(new_n973), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1177), .A2(new_n973), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1179), .B1(new_n1195), .B2(new_n920), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT127), .B1(new_n1191), .B2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1189), .A2(new_n1188), .A3(new_n1180), .A4(new_n1190), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1193), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT127), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(G375), .A2(G378), .ZN(new_n1203));
  INV_X1    g1003(.A(G213), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(G343), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1076), .A2(new_n1098), .A3(new_n1135), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n949), .B2(new_n1142), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT124), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1140), .A2(new_n1209), .A3(new_n1141), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n955), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1205), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1203), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1205), .A2(G2897), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT60), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1149), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1050), .A2(KEYINPUT60), .A3(new_n1054), .A4(new_n1052), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1216), .A2(new_n1056), .A3(new_n648), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1170), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(G384), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n797), .A2(new_n1218), .A3(new_n1170), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1214), .B1(new_n1222), .B2(KEYINPUT125), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT125), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1214), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1220), .A2(new_n1224), .A3(new_n1221), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1222), .A2(KEYINPUT125), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1223), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT61), .B1(new_n1213), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT62), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1203), .A2(new_n1212), .A3(new_n1230), .A4(new_n1222), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1203), .A2(new_n1212), .A3(new_n1222), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT62), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1229), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1198), .A2(new_n1202), .A3(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1232), .B(KEYINPUT63), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1236), .A2(new_n1200), .A3(new_n1199), .A4(new_n1229), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(G405));
  NAND2_X1  g1038(.A1(new_n1203), .A2(new_n1185), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1222), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1239), .B(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1241), .B(new_n1242), .ZN(G402));
endmodule


