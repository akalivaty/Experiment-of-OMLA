//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n188), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G116), .B(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  AOI21_X1  g020(.A(G101), .B1(new_n205), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n205), .A2(G107), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n204), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n205), .A2(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n209), .A2(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT75), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n201), .A2(KEYINPUT5), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n191), .A2(G119), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT5), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n196), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  AND4_X1   g040(.A1(new_n203), .A2(new_n216), .A3(new_n221), .A4(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G110), .B(G122), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT8), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n195), .A2(new_n202), .B1(new_n222), .B2(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n219), .A2(new_n220), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT80), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n203), .A2(new_n226), .ZN(new_n234));
  INV_X1    g048(.A(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n216), .A3(new_n221), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT80), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .A4(new_n229), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT1), .B1(new_n242), .B2(G146), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(G146), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G143), .ZN(new_n246));
  OAI211_X1 g060(.A(G128), .B(new_n243), .C1(new_n244), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(G146), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n248), .B(new_n249), .C1(KEYINPUT1), .C2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(G125), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT0), .A4(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n244), .A2(new_n246), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT0), .B(G128), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n252), .A2(new_n253), .B1(new_n257), .B2(G125), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n247), .A2(new_n251), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT79), .B1(new_n259), .B2(G125), .ZN(new_n260));
  INV_X1    g074(.A(G224), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT7), .B1(new_n261), .B2(G953), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n258), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n258), .B2(new_n260), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n240), .A2(new_n241), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n241), .B1(new_n240), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n206), .A2(new_n210), .A3(new_n214), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n206), .A2(new_n210), .A3(KEYINPUT74), .A4(new_n214), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n193), .A2(new_n194), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n203), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n212), .B1(new_n272), .B2(new_n273), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n220), .A2(KEYINPUT4), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT75), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT75), .B1(new_n219), .B2(new_n220), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n216), .A2(KEYINPUT76), .A3(new_n221), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n230), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT78), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n287), .A2(new_n288), .A3(new_n291), .A4(new_n230), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n283), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n228), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n269), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n292), .ZN(new_n296));
  INV_X1    g110(.A(new_n283), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n228), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT6), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n293), .B2(new_n228), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n301), .A3(new_n299), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n258), .A2(new_n260), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n261), .A2(G953), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n295), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n295), .B2(new_n308), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n187), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT82), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(KEYINPUT82), .B(new_n187), .C1(new_n310), .C2(new_n311), .ZN(new_n315));
  INV_X1    g129(.A(G469), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n247), .A2(new_n251), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT67), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n247), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n287), .A2(new_n321), .A3(new_n288), .A4(KEYINPUT10), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT11), .ZN(new_n323));
  INV_X1    g137(.A(G134), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(G137), .ZN(new_n325));
  INV_X1    g139(.A(G137), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT11), .A3(G134), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT64), .A3(G131), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT64), .A2(G131), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n327), .A3(new_n331), .A4(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n257), .B1(new_n274), .B2(new_n275), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n280), .B2(new_n281), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT10), .B1(new_n259), .B2(new_n235), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n322), .A2(new_n334), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n317), .A2(new_n231), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n285), .A2(new_n286), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n317), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT12), .B1(new_n342), .B2(new_n334), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT12), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n285), .A2(new_n259), .A3(new_n286), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n344), .B(new_n333), .C1(new_n345), .C2(new_n340), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n339), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G110), .B(G140), .ZN(new_n348));
  INV_X1    g162(.A(G953), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G227), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n348), .B(new_n350), .Z(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n322), .ZN(new_n353));
  INV_X1    g167(.A(new_n257), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n276), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n338), .B1(new_n355), .B2(new_n282), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n333), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n351), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n339), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G902), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n316), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n358), .B1(new_n357), .B2(new_n339), .ZN(new_n363));
  AND4_X1   g177(.A1(new_n339), .A2(new_n343), .A3(new_n346), .A4(new_n358), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n316), .B(new_n361), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT77), .ZN(new_n366));
  INV_X1    g180(.A(new_n339), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n274), .A2(G101), .ZN(new_n368));
  INV_X1    g182(.A(new_n281), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n337), .B1(new_n370), .B2(new_n335), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n334), .B1(new_n371), .B2(new_n322), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n351), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n339), .A2(new_n343), .A3(new_n346), .A4(new_n358), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n316), .A4(new_n361), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n362), .B1(new_n366), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G475), .ZN(new_n379));
  INV_X1    g193(.A(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G125), .ZN(new_n381));
  INV_X1    g195(.A(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G140), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT16), .ZN(new_n384));
  OR3_X1    g198(.A1(new_n382), .A2(KEYINPUT16), .A3(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n245), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(G146), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G131), .ZN(new_n391));
  INV_X1    g205(.A(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n349), .A3(G214), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n242), .ZN(new_n394));
  NOR2_X1   g208(.A1(G237), .A2(G953), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(G143), .A3(G214), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n391), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT17), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n391), .A3(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT85), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(new_n396), .ZN(new_n403));
  AND4_X1   g217(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT17), .A4(G131), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n397), .B2(KEYINPUT17), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n390), .B(new_n401), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT83), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n403), .B2(new_n407), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G125), .B(G140), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(new_n245), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n403), .A2(new_n407), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n406), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G113), .B(G122), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(new_n205), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n406), .A2(new_n418), .A3(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n379), .B1(new_n425), .B2(KEYINPUT86), .ZN(new_n426));
  INV_X1    g240(.A(new_n424), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n421), .B1(new_n406), .B2(new_n418), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n361), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(G475), .A2(G902), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n413), .B(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n433), .B1(new_n435), .B2(G146), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n413), .B(KEYINPUT19), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT84), .A3(new_n245), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n398), .A2(new_n400), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n388), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n421), .B1(new_n441), .B2(new_n418), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n432), .B1(new_n442), .B2(new_n427), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT20), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n388), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(new_n436), .B2(new_n438), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n416), .B1(new_n411), .B2(new_n409), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n422), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n424), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n432), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n426), .A2(new_n431), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n349), .A2(G952), .ZN(new_n453));
  NAND2_X1  g267(.A1(G234), .A2(G237), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT89), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(G902), .A3(G953), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(G898), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G122), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n463), .B2(G116), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(G116), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n191), .A3(G122), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n464), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  OAI21_X1  g284(.A(G107), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT88), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n473), .B(G107), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n191), .A2(G122), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n475), .A3(new_n209), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n242), .A2(G128), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n250), .A2(G143), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n477), .A2(new_n478), .A3(new_n324), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n324), .B1(new_n477), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n472), .A2(new_n474), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n478), .A3(new_n324), .ZN(new_n484));
  INV_X1    g298(.A(new_n476), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n209), .B1(new_n465), .B2(new_n475), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n242), .A2(G128), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT13), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n489), .B2(new_n477), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n242), .A2(KEYINPUT13), .A3(G128), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n324), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT9), .B(G234), .ZN(new_n495));
  INV_X1    g309(.A(G217), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n495), .A2(new_n496), .A3(G953), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n483), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n483), .B2(new_n494), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n361), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G478), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n501), .A2(KEYINPUT15), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n500), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n452), .A2(new_n462), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G221), .ZN(new_n505));
  INV_X1    g319(.A(new_n495), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(new_n361), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n378), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n314), .A2(new_n315), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT90), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n496), .B1(G234), .B2(new_n361), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n189), .A2(G128), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n250), .A2(KEYINPUT23), .A3(G119), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n189), .A2(G128), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(KEYINPUT23), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT72), .B(G110), .ZN(new_n516));
  XNOR2_X1  g330(.A(G119), .B(G128), .ZN(new_n517));
  INV_X1    g331(.A(G110), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT24), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G110), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI22_X1  g336(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n413), .A2(new_n245), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n388), .A3(new_n524), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n515), .A2(G110), .B1(new_n517), .B2(new_n522), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n527));
  AOI21_X1  g341(.A(G146), .B1(new_n384), .B2(new_n385), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n384), .A2(G146), .A3(new_n385), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n527), .B1(new_n389), .B2(new_n526), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n525), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n525), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n526), .B1(new_n529), .B2(new_n528), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT71), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n538), .B2(new_n530), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT22), .B(G137), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n349), .A2(G221), .A3(G234), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n539), .A2(KEYINPUT73), .A3(new_n544), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT25), .B1(new_n548), .B2(new_n361), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n550), .B(G902), .C1(new_n545), .C2(new_n547), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n511), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n511), .A2(G902), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(G472), .A2(G902), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n329), .A2(new_n391), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n391), .B1(G134), .B2(new_n326), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n328), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n247), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT67), .B1(new_n247), .B2(new_n251), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n333), .A2(new_n354), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT30), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n257), .B1(new_n330), .B2(new_n332), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT65), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n317), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n329), .A2(new_n391), .B1(new_n328), .B2(new_n558), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT65), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n565), .B(new_n278), .C1(new_n571), .C2(KEYINPUT30), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n395), .A2(G210), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT27), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT26), .B(G101), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n575), .B(new_n576), .Z(new_n577));
  AOI21_X1  g391(.A(new_n566), .B1(new_n321), .B2(new_n560), .ZN(new_n578));
  INV_X1    g392(.A(new_n278), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n572), .A2(new_n573), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT68), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n572), .A2(new_n580), .A3(KEYINPUT68), .A4(new_n573), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n572), .A2(new_n580), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT31), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT28), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n259), .B1(KEYINPUT65), .B2(new_n569), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n560), .A2(new_n567), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n564), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n278), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n563), .A2(new_n579), .A3(new_n564), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n588), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n577), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n587), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n556), .B1(new_n585), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT32), .ZN(new_n601));
  INV_X1    g415(.A(new_n556), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n593), .B1(new_n571), .B2(new_n579), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT28), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n595), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n605), .A2(new_n577), .B1(new_n586), .B2(KEYINPUT31), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n583), .A2(new_n584), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT32), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n565), .A2(new_n278), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n560), .A2(new_n567), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n570), .A3(new_n259), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT30), .B1(new_n614), .B2(new_n564), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n593), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT29), .B1(new_n616), .B2(new_n577), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT69), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n595), .A2(new_n598), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n594), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n577), .B1(new_n593), .B2(new_n588), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n604), .A2(KEYINPUT69), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n617), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT70), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT70), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n617), .A2(new_n620), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n621), .A2(KEYINPUT29), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n563), .A2(new_n579), .A3(new_n564), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n579), .B1(new_n563), .B2(new_n564), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT28), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n624), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n555), .B1(new_n611), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT90), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n314), .A2(new_n315), .A3(new_n635), .A4(new_n508), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n510), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  NOR2_X1   g452(.A1(new_n378), .A2(new_n507), .ZN(new_n639));
  INV_X1    g453(.A(new_n554), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n544), .B1(new_n533), .B2(new_n534), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n361), .B1(new_n643), .B2(new_n546), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n550), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n548), .A2(KEYINPUT25), .A3(new_n361), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n640), .B1(new_n647), .B2(new_n511), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n639), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(G472), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n361), .B1(new_n585), .B2(new_n599), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT91), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT92), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(new_n600), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n653), .B(KEYINPUT92), .C1(new_n652), .C2(new_n651), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n649), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT93), .Z(new_n659));
  AOI21_X1  g473(.A(KEYINPUT95), .B1(new_n500), .B2(new_n501), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n481), .B1(new_n471), .B2(KEYINPUT88), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n493), .B1(new_n661), .B2(new_n474), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT94), .B1(new_n662), .B2(new_n497), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n663), .B(KEYINPUT33), .C1(new_n498), .C2(new_n499), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n483), .A2(new_n494), .ZN(new_n665));
  INV_X1    g479(.A(new_n497), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n662), .A2(new_n497), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT33), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n667), .B(new_n668), .C1(KEYINPUT94), .C2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n501), .A2(G902), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n660), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n672), .ZN(new_n674));
  AOI211_X1 g488(.A(KEYINPUT95), .B(new_n674), .C1(new_n664), .C2(new_n670), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT96), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT95), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n671), .A2(new_n677), .A3(new_n672), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT96), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n674), .B1(new_n664), .B2(new_n670), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n660), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(G475), .B1(new_n429), .B2(new_n430), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n425), .A2(KEYINPUT86), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n450), .B1(new_n449), .B2(new_n432), .ZN(new_n685));
  INV_X1    g499(.A(new_n432), .ZN(new_n686));
  AOI211_X1 g500(.A(KEYINPUT20), .B(new_n686), .C1(new_n448), .C2(new_n424), .ZN(new_n687));
  OAI22_X1  g501(.A1(new_n683), .A2(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n682), .A2(new_n462), .A3(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n659), .A2(new_n312), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT97), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT34), .B(G104), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G6));
  INV_X1    g507(.A(new_n187), .ZN(new_n694));
  INV_X1    g508(.A(new_n309), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n696));
  INV_X1    g510(.A(new_n268), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n240), .A2(new_n266), .A3(new_n241), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n294), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n361), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n695), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n295), .A2(new_n308), .A3(new_n309), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n694), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT98), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n688), .A2(new_n461), .A3(new_n503), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n705), .B(new_n187), .C1(new_n310), .C2(new_n311), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT98), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n659), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT35), .B(G107), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G9));
  NOR2_X1   g525(.A1(new_n544), .A2(KEYINPUT36), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n533), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n553), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n647), .B2(new_n511), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n656), .B2(new_n657), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n510), .A2(new_n636), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT37), .B(G110), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G12));
  NOR3_X1   g534(.A1(new_n716), .A2(new_n378), .A3(new_n507), .ZN(new_n721));
  INV_X1    g535(.A(new_n610), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n608), .A2(new_n609), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n633), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n503), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n452), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n456), .B1(G900), .B2(new_n457), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT99), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n721), .A2(new_n724), .A3(new_n703), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT100), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n362), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n365), .A2(KEYINPUT77), .ZN(new_n734));
  AOI21_X1  g548(.A(G902), .B1(new_n373), .B2(new_n374), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n376), .B1(new_n735), .B2(new_n316), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n733), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n552), .A2(new_n714), .ZN(new_n738));
  INV_X1    g552(.A(new_n507), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n601), .A2(new_n610), .B1(new_n632), .B2(G472), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT100), .A3(new_n703), .A4(new_n729), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n732), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT101), .B(G128), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G30));
  XOR2_X1   g560(.A(new_n728), .B(KEYINPUT39), .Z(new_n747));
  NAND2_X1  g561(.A1(new_n639), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT40), .Z(new_n749));
  NOR2_X1   g563(.A1(new_n310), .A2(new_n311), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT38), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n628), .A2(new_n629), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n753), .A2(new_n577), .B1(new_n572), .B2(new_n580), .ZN(new_n754));
  OAI21_X1  g568(.A(G472), .B1(new_n754), .B2(G902), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n611), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n688), .A2(new_n725), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n738), .A2(new_n694), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n749), .A2(new_n752), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT102), .B(G143), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G45));
  AOI211_X1 g575(.A(new_n728), .B(new_n452), .C1(new_n676), .C2(new_n681), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n721), .A2(new_n724), .A3(new_n703), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G146), .ZN(G48));
  NOR2_X1   g578(.A1(new_n312), .A2(new_n689), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n366), .A2(new_n377), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT103), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n375), .A2(new_n361), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n507), .B1(new_n768), .B2(G469), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n765), .A2(new_n772), .A3(new_n634), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT41), .B(G113), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G15));
  NAND2_X1  g589(.A1(new_n708), .A2(new_n706), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n766), .A2(new_n769), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT103), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n724), .A2(new_n778), .A3(new_n648), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G116), .ZN(G18));
  NOR3_X1   g596(.A1(new_n688), .A2(new_n461), .A3(new_n725), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n738), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n777), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n724), .A3(new_n703), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G119), .ZN(G21));
  AOI211_X1 g602(.A(new_n694), .B(new_n757), .C1(new_n701), .C2(new_n702), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n598), .B1(new_n630), .B2(new_n595), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(KEYINPUT31), .B2(new_n586), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n607), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n556), .B(KEYINPUT104), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(G902), .B1(new_n606), .B2(new_n607), .ZN(new_n795));
  OAI22_X1  g609(.A1(new_n792), .A2(new_n794), .B1(new_n795), .B2(new_n650), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n555), .A3(new_n461), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n772), .A2(new_n789), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G122), .ZN(G24));
  NOR2_X1   g613(.A1(new_n796), .A2(new_n716), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n762), .A3(new_n703), .A4(new_n786), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G125), .ZN(G27));
  INV_X1    g616(.A(KEYINPUT42), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n310), .A2(new_n311), .A3(new_n694), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT105), .B1(new_n347), .B2(new_n351), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n360), .B2(KEYINPUT105), .ZN(new_n806));
  OAI21_X1  g620(.A(G469), .B1(new_n806), .B2(G902), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n507), .B1(new_n807), .B2(new_n766), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n724), .A2(new_n804), .A3(new_n648), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n762), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n804), .A2(new_n808), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT42), .A3(new_n634), .A4(new_n762), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G131), .ZN(G33));
  NAND4_X1  g629(.A1(new_n634), .A2(new_n729), .A3(new_n808), .A4(new_n804), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G134), .ZN(G36));
  AOI21_X1  g631(.A(KEYINPUT45), .B1(new_n352), .B2(new_n359), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n316), .B(new_n818), .C1(KEYINPUT45), .C2(new_n806), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n316), .A2(new_n361), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(KEYINPUT46), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n766), .B1(new_n821), .B2(KEYINPUT46), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n739), .A3(new_n747), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n682), .A2(new_n452), .ZN(new_n826));
  NAND2_X1  g640(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n656), .A3(new_n657), .A4(new_n738), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT44), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n804), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n825), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n832), .B2(new_n831), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G137), .ZN(G39));
  NAND3_X1  g651(.A1(new_n824), .A2(KEYINPUT47), .A3(new_n739), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n739), .B1(new_n822), .B2(new_n823), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT47), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n834), .A2(new_n810), .A3(new_n724), .A4(new_n648), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G140), .ZN(G42));
  INV_X1    g659(.A(KEYINPUT108), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n773), .A2(new_n798), .A3(new_n787), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n724), .A2(new_n778), .A3(new_n648), .A4(new_n779), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n706), .B2(new_n708), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n794), .B1(new_n791), .B2(new_n607), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n651), .B2(G472), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n648), .A3(new_n462), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n770), .A3(new_n771), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n312), .A2(new_n777), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n741), .A2(new_n784), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n854), .A2(new_n789), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n781), .A3(KEYINPUT108), .A4(new_n773), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n688), .A2(new_n725), .A3(new_n728), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n721), .A2(new_n724), .A3(new_n804), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n816), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n800), .A2(new_n762), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n804), .A2(new_n808), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT109), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT109), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n812), .A2(new_n865), .A3(new_n762), .A4(new_n800), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n861), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n850), .A2(new_n858), .A3(new_n867), .A4(new_n814), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n314), .A2(new_n315), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n682), .A2(new_n688), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n726), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n658), .A2(new_n869), .A3(new_n462), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n637), .A2(new_n718), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT110), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n850), .A2(new_n858), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT110), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n637), .A2(new_n718), .A3(new_n872), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n866), .A2(new_n864), .ZN(new_n878));
  INV_X1    g692(.A(new_n861), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n814), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n763), .A2(new_n801), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n732), .B2(new_n743), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n738), .A2(new_n728), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n789), .A2(new_n756), .A3(new_n808), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n884), .A2(KEYINPUT52), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n874), .A2(new_n882), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT111), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT53), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n892), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(new_n456), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n830), .A2(new_n648), .A3(new_n897), .A4(new_n852), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n834), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n766), .B1(new_n316), .B2(new_n735), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n739), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n842), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n751), .A2(new_n694), .A3(new_n786), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT115), .B1(new_n903), .B2(new_n898), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT50), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n830), .A2(new_n897), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n834), .A2(new_n777), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n800), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n756), .A2(new_n555), .A3(new_n456), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n910), .A2(new_n688), .A3(new_n682), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n902), .A2(new_n905), .A3(new_n908), .A4(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n855), .ZN(new_n915));
  OAI22_X1  g729(.A1(new_n898), .A2(new_n915), .B1(new_n910), .B2(new_n870), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n906), .A2(new_n634), .A3(new_n907), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT48), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(KEYINPUT48), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n912), .A2(KEYINPUT116), .A3(new_n913), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT116), .B1(new_n912), .B2(new_n913), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT53), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n773), .A2(new_n798), .A3(new_n787), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n814), .A2(new_n926), .A3(new_n781), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT113), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n814), .A2(new_n926), .A3(KEYINPUT113), .A4(new_n781), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(KEYINPUT53), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT52), .B1(new_n884), .B2(new_n886), .ZN(new_n932));
  INV_X1    g746(.A(new_n883), .ZN(new_n933));
  AND4_X1   g747(.A1(KEYINPUT52), .A2(new_n744), .A3(new_n933), .A4(new_n886), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n867), .A2(new_n637), .A3(new_n718), .A4(new_n872), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT112), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  AOI22_X1  g753(.A1(new_n892), .A2(new_n925), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n896), .A2(new_n924), .A3(KEYINPUT117), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(G953), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT117), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n896), .A2(new_n924), .A3(new_n945), .A4(new_n942), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n453), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n648), .A2(new_n187), .A3(new_n739), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT107), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n900), .B(KEYINPUT49), .Z(new_n950));
  NOR2_X1   g764(.A1(new_n756), .A2(new_n826), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n751), .A4(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n944), .A2(new_n947), .A3(new_n952), .ZN(G75));
  NOR2_X1   g767(.A1(new_n349), .A2(G952), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT118), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n940), .A2(new_n361), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT56), .B1(new_n957), .B2(G210), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n303), .A2(new_n304), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n307), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT55), .Z(new_n961));
  OR2_X1    g775(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n961), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n956), .B1(new_n962), .B2(new_n963), .ZN(G51));
  XNOR2_X1  g778(.A(new_n820), .B(KEYINPUT57), .ZN(new_n965));
  INV_X1    g779(.A(new_n941), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n850), .A2(new_n858), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n967), .A2(new_n873), .A3(new_n880), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n935), .B1(new_n968), .B2(new_n876), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT53), .B1(new_n969), .B2(new_n874), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n929), .A4(new_n930), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n937), .B(KEYINPUT112), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n966), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n892), .A2(new_n925), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n936), .A2(new_n939), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT119), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n941), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n940), .B2(new_n941), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n965), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n375), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n957), .A2(new_n819), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n954), .B1(new_n982), .B2(new_n983), .ZN(G54));
  AND2_X1   g798(.A1(KEYINPUT58), .A2(G475), .ZN(new_n985));
  OAI211_X1 g799(.A(G902), .B(new_n985), .C1(new_n970), .C2(new_n973), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n424), .A3(new_n448), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n957), .A2(new_n449), .A3(new_n985), .ZN(new_n988));
  INV_X1    g802(.A(new_n954), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT120), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT120), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n987), .A2(new_n988), .A3(new_n992), .A4(new_n989), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(G60));
  XOR2_X1   g808(.A(new_n671), .B(KEYINPUT121), .Z(new_n995));
  AOI22_X1  g809(.A1(new_n895), .A2(KEYINPUT54), .B1(new_n940), .B2(new_n941), .ZN(new_n996));
  NAND2_X1  g810(.A1(G478), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT59), .Z(new_n998));
  OAI21_X1  g812(.A(new_n995), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n995), .A2(new_n998), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n979), .B2(new_n980), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n999), .A2(new_n955), .A3(new_n1001), .ZN(G63));
  NAND2_X1  g816(.A1(G217), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT60), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n713), .B(new_n1005), .C1(new_n970), .C2(new_n973), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n940), .A2(new_n1004), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1006), .B(new_n955), .C1(new_n1007), .C2(new_n548), .ZN(new_n1008));
  XNOR2_X1  g822(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1008), .A2(KEYINPUT122), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1008), .B2(KEYINPUT122), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1010), .A2(new_n1011), .ZN(G66));
  NAND2_X1  g826(.A1(new_n875), .A2(new_n877), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n349), .ZN(new_n1014));
  OAI21_X1  g828(.A(G953), .B1(new_n459), .B2(new_n261), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n959), .B1(G898), .B2(new_n349), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT124), .Z(new_n1018));
  XNOR2_X1  g832(.A(new_n1016), .B(new_n1018), .ZN(G69));
  OAI21_X1  g833(.A(new_n565), .B1(new_n571), .B2(KEYINPUT30), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(new_n435), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G900), .A2(G953), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n836), .A2(new_n844), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n814), .A2(new_n816), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT126), .ZN(new_n1025));
  INV_X1    g839(.A(new_n825), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n634), .A3(new_n789), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1023), .A2(new_n884), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1021), .B(new_n1022), .C1(new_n1028), .C2(G953), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n759), .A2(new_n884), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1032));
  INV_X1    g846(.A(new_n634), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n871), .B(KEYINPUT125), .ZN(new_n1034));
  OR4_X1    g848(.A1(new_n1033), .A2(new_n1034), .A3(new_n748), .A4(new_n834), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1023), .A2(new_n1031), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  AND2_X1   g850(.A1(new_n1036), .A2(new_n349), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1029), .B1(new_n1037), .B2(new_n1021), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n349), .B1(G227), .B2(G900), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(G72));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT63), .Z(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n1036), .B2(new_n1013), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n616), .B(KEYINPUT127), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1043), .A2(new_n598), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1042), .B1(new_n1028), .B2(new_n1013), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1044), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1046), .A2(new_n577), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n616), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n586), .B1(new_n1049), .B2(new_n598), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n895), .A2(new_n1042), .A3(new_n1050), .ZN(new_n1051));
  AND4_X1   g865(.A1(new_n989), .A2(new_n1045), .A3(new_n1048), .A4(new_n1051), .ZN(G57));
endmodule


