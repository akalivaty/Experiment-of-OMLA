

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  INV_X1 U322 ( .A(G106GAT), .ZN(n362) );
  XNOR2_X1 U323 ( .A(n363), .B(n362), .ZN(n365) );
  XNOR2_X1 U324 ( .A(n365), .B(n364), .ZN(n409) );
  XNOR2_X1 U325 ( .A(n367), .B(n395), .ZN(n368) );
  NOR2_X1 U326 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U327 ( .A(n369), .B(n368), .ZN(n372) );
  NOR2_X1 U328 ( .A1(n512), .A2(n426), .ZN(n566) );
  XOR2_X1 U329 ( .A(n377), .B(n376), .Z(n572) );
  NOR2_X1 U330 ( .A1(n466), .A2(n446), .ZN(n558) );
  XOR2_X1 U331 ( .A(n463), .B(KEYINPUT28), .Z(n527) );
  XNOR2_X1 U332 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U333 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(G71GAT), .B(KEYINPUT83), .Z(n291) );
  XNOR2_X1 U335 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n291), .B(n290), .ZN(n309) );
  XOR2_X1 U337 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n293) );
  XNOR2_X1 U338 ( .A(G134GAT), .B(G190GAT), .ZN(n292) );
  XNOR2_X1 U339 ( .A(n293), .B(n292), .ZN(n295) );
  XOR2_X1 U340 ( .A(G43GAT), .B(G99GAT), .Z(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n305) );
  XOR2_X1 U342 ( .A(G183GAT), .B(KEYINPUT17), .Z(n297) );
  XNOR2_X1 U343 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n331) );
  XOR2_X1 U345 ( .A(G127GAT), .B(KEYINPUT0), .Z(n299) );
  XNOR2_X1 U346 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n311) );
  XNOR2_X1 U348 ( .A(n331), .B(n311), .ZN(n303) );
  XOR2_X1 U349 ( .A(G176GAT), .B(G120GAT), .Z(n301) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G113GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n307) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(n309), .B(n308), .Z(n466) );
  INV_X1 U357 ( .A(KEYINPUT55), .ZN(n445) );
  XNOR2_X1 U358 ( .A(G120GAT), .B(G148GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n310), .B(G57GAT), .ZN(n370) );
  XNOR2_X1 U360 ( .A(n311), .B(n370), .ZN(n330) );
  XOR2_X1 U361 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n313) );
  XNOR2_X1 U362 ( .A(KEYINPUT93), .B(KEYINPUT4), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U364 ( .A(KEYINPUT94), .B(KEYINPUT1), .Z(n315) );
  XNOR2_X1 U365 ( .A(KEYINPUT90), .B(KEYINPUT92), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U367 ( .A(n317), .B(n316), .Z(n328) );
  XOR2_X1 U368 ( .A(G155GAT), .B(KEYINPUT2), .Z(n319) );
  XNOR2_X1 U369 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n433) );
  XOR2_X1 U371 ( .A(n433), .B(KEYINPUT5), .Z(n321) );
  NAND2_X1 U372 ( .A1(G225GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U374 ( .A(G134GAT), .B(G162GAT), .Z(n410) );
  XOR2_X1 U375 ( .A(n410), .B(G85GAT), .Z(n324) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(G113GAT), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n322), .B(G1GAT), .ZN(n353) );
  XNOR2_X1 U378 ( .A(G29GAT), .B(n353), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n461) );
  XNOR2_X1 U383 ( .A(KEYINPUT95), .B(n461), .ZN(n512) );
  XOR2_X1 U384 ( .A(n331), .B(KEYINPUT96), .Z(n333) );
  NAND2_X1 U385 ( .A1(G226GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U387 ( .A(n334), .B(G92GAT), .Z(n336) );
  XOR2_X1 U388 ( .A(G169GAT), .B(G8GAT), .Z(n354) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(n354), .ZN(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U391 ( .A(G190GAT), .B(G218GAT), .Z(n402) );
  XOR2_X1 U392 ( .A(n337), .B(n402), .Z(n343) );
  XNOR2_X1 U393 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n338), .B(KEYINPUT86), .ZN(n339) );
  XOR2_X1 U395 ( .A(n339), .B(KEYINPUT87), .Z(n341) );
  XNOR2_X1 U396 ( .A(G197GAT), .B(G204GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n441) );
  XOR2_X1 U398 ( .A(G176GAT), .B(G64GAT), .Z(n366) );
  XNOR2_X1 U399 ( .A(n441), .B(n366), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n455) );
  XOR2_X1 U401 ( .A(G29GAT), .B(G36GAT), .Z(n345) );
  XNOR2_X1 U402 ( .A(G50GAT), .B(G43GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U404 ( .A(KEYINPUT7), .B(KEYINPUT68), .Z(n347) );
  XNOR2_X1 U405 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U407 ( .A(n349), .B(n348), .Z(n414) );
  XOR2_X1 U408 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n351) );
  XNOR2_X1 U409 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n414), .B(n352), .ZN(n361) );
  XOR2_X1 U412 ( .A(n354), .B(n353), .Z(n356) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U415 ( .A(G22GAT), .B(G15GAT), .Z(n383) );
  XOR2_X1 U416 ( .A(n357), .B(n383), .Z(n359) );
  XNOR2_X1 U417 ( .A(G197GAT), .B(KEYINPUT65), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U419 ( .A(n361), .B(n360), .Z(n567) );
  XNOR2_X1 U420 ( .A(G99GAT), .B(G85GAT), .ZN(n363) );
  XOR2_X1 U421 ( .A(KEYINPUT72), .B(G92GAT), .Z(n364) );
  XNOR2_X1 U422 ( .A(G204GAT), .B(n409), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n366), .B(KEYINPUT32), .ZN(n367) );
  XOR2_X1 U424 ( .A(G71GAT), .B(KEYINPUT13), .Z(n395) );
  XOR2_X1 U425 ( .A(KEYINPUT71), .B(G78GAT), .Z(n430) );
  XNOR2_X1 U426 ( .A(n430), .B(n370), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n377) );
  XOR2_X1 U428 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n374) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U431 ( .A(KEYINPUT73), .B(n375), .Z(n376) );
  XNOR2_X1 U432 ( .A(KEYINPUT41), .B(n572), .ZN(n544) );
  NOR2_X1 U433 ( .A1(n567), .A2(n544), .ZN(n379) );
  XOR2_X1 U434 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n400) );
  XOR2_X1 U436 ( .A(G57GAT), .B(G78GAT), .Z(n381) );
  XNOR2_X1 U437 ( .A(G127GAT), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U439 ( .A(n382), .B(G155GAT), .Z(n385) );
  XNOR2_X1 U440 ( .A(n383), .B(G183GAT), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n399) );
  XOR2_X1 U442 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n387) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U445 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n389) );
  XNOR2_X1 U446 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U448 ( .A(n391), .B(n390), .Z(n397) );
  XOR2_X1 U449 ( .A(KEYINPUT77), .B(G64GAT), .Z(n393) );
  XNOR2_X1 U450 ( .A(G8GAT), .B(G1GAT), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n576) );
  NAND2_X1 U455 ( .A1(n400), .A2(n576), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n401), .B(KEYINPUT115), .ZN(n415) );
  XOR2_X1 U457 ( .A(KEYINPUT64), .B(n402), .Z(n404) );
  NAND2_X1 U458 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U460 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n406) );
  XNOR2_X1 U461 ( .A(KEYINPUT74), .B(KEYINPUT10), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U463 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n414), .B(n413), .ZN(n550) );
  NAND2_X1 U467 ( .A1(n415), .A2(n550), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n416), .B(KEYINPUT47), .ZN(n423) );
  XOR2_X1 U469 ( .A(KEYINPUT45), .B(KEYINPUT116), .Z(n419) );
  INV_X1 U470 ( .A(n576), .ZN(n556) );
  XNOR2_X1 U471 ( .A(KEYINPUT36), .B(KEYINPUT105), .ZN(n417) );
  XOR2_X1 U472 ( .A(KEYINPUT75), .B(n550), .Z(n560) );
  XNOR2_X1 U473 ( .A(n417), .B(n560), .ZN(n579) );
  NAND2_X1 U474 ( .A1(n556), .A2(n579), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U476 ( .A(KEYINPUT70), .B(n567), .ZN(n521) );
  NAND2_X1 U477 ( .A1(n420), .A2(n521), .ZN(n421) );
  NOR2_X1 U478 ( .A1(n572), .A2(n421), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n424), .B(KEYINPUT48), .ZN(n523) );
  NOR2_X1 U480 ( .A1(n455), .A2(n523), .ZN(n425) );
  XOR2_X1 U481 ( .A(n425), .B(KEYINPUT54), .Z(n426) );
  XOR2_X1 U482 ( .A(G148GAT), .B(G162GAT), .Z(n428) );
  XNOR2_X1 U483 ( .A(G141GAT), .B(G106GAT), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U485 ( .A(n429), .B(G218GAT), .Z(n432) );
  XNOR2_X1 U486 ( .A(G50GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n437) );
  XOR2_X1 U488 ( .A(G22GAT), .B(n433), .Z(n435) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U491 ( .A(n437), .B(n436), .Z(n443) );
  XOR2_X1 U492 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n439) );
  XNOR2_X1 U493 ( .A(KEYINPUT89), .B(KEYINPUT22), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n463) );
  NAND2_X1 U497 ( .A1(n566), .A2(n463), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U499 ( .A(n544), .ZN(n529) );
  NAND2_X1 U500 ( .A1(n558), .A2(n529), .ZN(n450) );
  XOR2_X1 U501 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n448) );
  XNOR2_X1 U502 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n447) );
  XOR2_X1 U503 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n471) );
  OR2_X1 U504 ( .A1(n521), .A2(n572), .ZN(n485) );
  XOR2_X1 U505 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n452) );
  NAND2_X1 U506 ( .A1(n556), .A2(n560), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n469) );
  XNOR2_X1 U508 ( .A(n455), .B(KEYINPUT97), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n453), .B(KEYINPUT27), .ZN(n464) );
  INV_X1 U510 ( .A(n466), .ZN(n524) );
  NOR2_X1 U511 ( .A1(n524), .A2(n463), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT26), .ZN(n565) );
  NAND2_X1 U513 ( .A1(n464), .A2(n565), .ZN(n460) );
  INV_X1 U514 ( .A(n455), .ZN(n514) );
  NAND2_X1 U515 ( .A1(n524), .A2(n514), .ZN(n456) );
  NAND2_X1 U516 ( .A1(n456), .A2(n463), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n457), .B(KEYINPUT25), .ZN(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT98), .B(n458), .Z(n459) );
  NAND2_X1 U519 ( .A1(n460), .A2(n459), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n462), .A2(n461), .ZN(n468) );
  NAND2_X1 U521 ( .A1(n464), .A2(n512), .ZN(n522) );
  NOR2_X1 U522 ( .A1(n527), .A2(n522), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n482) );
  NAND2_X1 U525 ( .A1(n469), .A2(n482), .ZN(n497) );
  NOR2_X1 U526 ( .A1(n485), .A2(n497), .ZN(n480) );
  NAND2_X1 U527 ( .A1(n480), .A2(n512), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n472), .ZN(G1324GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n474) );
  NAND2_X1 U531 ( .A1(n480), .A2(n514), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(n475), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U535 ( .A1(n480), .A2(n524), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT102), .Z(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n480), .A2(n527), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U541 ( .A(G29GAT), .B(KEYINPUT39), .Z(n489) );
  XOR2_X1 U542 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n487) );
  NAND2_X1 U543 ( .A1(n579), .A2(n482), .ZN(n483) );
  NOR2_X1 U544 ( .A1(n556), .A2(n483), .ZN(n484) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n484), .ZN(n511) );
  OR2_X1 U546 ( .A1(n485), .A2(n511), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n495) );
  NAND2_X1 U548 ( .A1(n495), .A2(n512), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT104), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U551 ( .A1(n514), .A2(n495), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n493) );
  NAND2_X1 U554 ( .A1(n495), .A2(n524), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n495), .A2(n527), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n529), .A2(n567), .ZN(n510) );
  NOR2_X1 U561 ( .A1(n497), .A2(n510), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT108), .ZN(n506) );
  NAND2_X1 U563 ( .A1(n512), .A2(n506), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n502) );
  NAND2_X1 U566 ( .A1(n506), .A2(n514), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n503), .ZN(G1333GAT) );
  XOR2_X1 U569 ( .A(G71GAT), .B(KEYINPUT111), .Z(n505) );
  NAND2_X1 U570 ( .A1(n506), .A2(n524), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U573 ( .A1(n527), .A2(n506), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n517) );
  NAND2_X1 U577 ( .A1(n517), .A2(n512), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n517), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U581 ( .A1(n524), .A2(n517), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n527), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  INV_X1 U587 ( .A(n521), .ZN(n554) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n540) );
  NAND2_X1 U589 ( .A1(n540), .A2(n524), .ZN(n525) );
  XOR2_X1 U590 ( .A(KEYINPUT117), .B(n525), .Z(n526) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n554), .A2(n534), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U595 ( .A1(n534), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NAND2_X1 U597 ( .A1(n534), .A2(n556), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  INV_X1 U600 ( .A(n534), .ZN(n535) );
  NOR2_X1 U601 ( .A1(n535), .A2(n560), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n537) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT119), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n540), .A2(n565), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n567), .A2(n549), .ZN(n541) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n541), .Z(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n543) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n546) );
  NOR2_X1 U612 ( .A1(n544), .A2(n549), .ZN(n545) );
  XOR2_X1 U613 ( .A(n546), .B(n545), .Z(G1345GAT) );
  NOR2_X1 U614 ( .A1(n576), .A2(n549), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n558), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U625 ( .A(n558), .ZN(n559) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n564) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT125), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT126), .B(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n575) );
  NOR2_X1 U632 ( .A1(n575), .A2(n567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  INV_X1 U637 ( .A(n575), .ZN(n578) );
  AND2_X1 U638 ( .A1(n572), .A2(n578), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

