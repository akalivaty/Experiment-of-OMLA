//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT64), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G143), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT68), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n187), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n191), .A2(G128), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT69), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n205), .B1(new_n202), .B2(G143), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n193), .A2(new_n195), .A3(G128), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT69), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n204), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT71), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G137), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G134), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n216), .A2(G137), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(KEYINPUT11), .ZN(new_n224));
  OAI211_X1 g038(.A(KEYINPUT66), .B(new_n220), .C1(new_n216), .C2(G137), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n218), .A2(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n229), .B2(new_n223), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n208), .A2(new_n209), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n211), .A2(KEYINPUT69), .A3(new_n212), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n204), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n215), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n225), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT66), .B1(new_n219), .B2(new_n220), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(KEYINPUT67), .B(G131), .C1(new_n241), .C2(new_n221), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n226), .B1(new_n243), .B2(new_n227), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n203), .A2(new_n248), .B1(new_n211), .B2(new_n246), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n238), .A2(KEYINPUT30), .A3(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT2), .B(G113), .Z(new_n252));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n253));
  XNOR2_X1  g067(.A(G116), .B(G119), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G116), .ZN(new_n257));
  INV_X1    g071(.A(G116), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G119), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT2), .B(G113), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT70), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n249), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n188), .A2(new_n190), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n200), .B1(new_n268), .B2(new_n199), .ZN(new_n269));
  INV_X1    g083(.A(new_n248), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n191), .A2(new_n206), .A3(new_n246), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT65), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n245), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n233), .A2(new_n234), .B1(new_n198), .B2(new_n203), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(new_n231), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n265), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n251), .A2(new_n264), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n238), .A2(new_n263), .A3(new_n250), .ZN(new_n279));
  INV_X1    g093(.A(G237), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G210), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n282), .B(KEYINPUT27), .Z(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G101), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT31), .B1(new_n278), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n279), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n264), .B1(new_n274), .B2(new_n276), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n279), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n285), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n287), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n251), .A2(new_n264), .A3(new_n277), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n300));
  INV_X1    g114(.A(G472), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT72), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n300), .B1(new_n299), .B2(new_n304), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n297), .A2(new_n279), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n285), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(KEYINPUT74), .A3(new_n285), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n285), .B1(new_n279), .B2(new_n289), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT73), .B1(new_n315), .B2(new_n293), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n279), .A2(new_n292), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n314), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT75), .B1(new_n313), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT74), .B1(new_n308), .B2(new_n285), .ZN(new_n324));
  AOI211_X1 g138(.A(new_n310), .B(new_n286), .C1(new_n297), .C2(new_n279), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n314), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT29), .B1(new_n328), .B2(KEYINPUT73), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n326), .A2(new_n327), .A3(new_n321), .A4(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n315), .A2(new_n317), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n238), .A2(new_n263), .A3(new_n250), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n263), .B1(new_n238), .B2(new_n250), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT28), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G902), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n323), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n307), .B1(new_n336), .B2(G472), .ZN(new_n337));
  INV_X1    g151(.A(G128), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n339));
  OAI211_X1 g153(.A(G119), .B(new_n338), .C1(new_n339), .C2(KEYINPUT23), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n256), .B2(G128), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n256), .B2(G128), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G110), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT24), .B(G110), .Z(new_n348));
  XNOR2_X1  g162(.A(G119), .B(G128), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT76), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT16), .ZN(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G125), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n355), .A2(KEYINPUT16), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(G146), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(G146), .B1(new_n353), .B2(new_n356), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n347), .B(new_n351), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n353), .A2(KEYINPUT79), .A3(new_n356), .A4(G146), .ZN(new_n363));
  INV_X1    g177(.A(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n355), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n352), .A2(KEYINPUT80), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(new_n202), .ZN(new_n370));
  OAI22_X1  g184(.A1(new_n344), .A2(G110), .B1(new_n349), .B2(new_n348), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n362), .A2(new_n363), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n372), .A2(new_n373), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n360), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT22), .B(G137), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n360), .B(new_n379), .C1(new_n374), .C2(new_n375), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n302), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(KEYINPUT25), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n385), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(new_n382), .A3(new_n302), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(G234), .B2(new_n302), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n382), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n391), .A2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n392), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n337), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  INV_X1    g213(.A(G104), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G107), .ZN(new_n402));
  INV_X1    g216(.A(G107), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT83), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(G104), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(KEYINPUT83), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n401), .A2(G107), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n412));
  AOI21_X1  g226(.A(G101), .B1(new_n400), .B2(G107), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT85), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(G107), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n406), .B1(new_n416), .B2(G104), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G101), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n398), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n215), .A2(new_n237), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n245), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n416), .A2(new_n408), .B1(KEYINPUT3), .B2(new_n406), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n426), .B2(new_n413), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n400), .A2(G107), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n411), .A2(new_n412), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G101), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n425), .A3(G101), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT84), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n429), .A2(new_n435), .A3(new_n425), .A4(G101), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n249), .B(new_n431), .C1(new_n434), .C2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n211), .ZN(new_n439));
  OAI21_X1  g253(.A(G128), .B1(new_n200), .B2(new_n192), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n233), .A2(new_n234), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n418), .A2(new_n420), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n398), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n423), .A2(new_n424), .A3(new_n438), .A4(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G140), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n281), .A2(G227), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n445), .B(new_n446), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n415), .A2(new_n421), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT86), .B1(new_n450), .B2(new_n214), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n441), .A2(new_n442), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n275), .A2(new_n453), .A3(new_n415), .A4(new_n421), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n245), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n455), .A2(KEYINPUT87), .A3(new_n457), .A4(new_n245), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n449), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n423), .A2(new_n438), .A3(new_n443), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n245), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n444), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n447), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G469), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n302), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n460), .A2(new_n444), .A3(new_n461), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n447), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n444), .A2(new_n448), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n444), .A2(KEYINPUT88), .A3(new_n448), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n464), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(G469), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n468), .A2(new_n302), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n469), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G122), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI221_X4 g297(.A(new_n263), .B1(new_n427), .B2(new_n430), .C1(new_n433), .C2(new_n436), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n485), .A2(G113), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n254), .A2(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n260), .B2(new_n261), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n415), .B2(new_n421), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n483), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n264), .B(new_n431), .C1(new_n434), .C2(new_n437), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n486), .A2(new_n487), .B1(new_n254), .B2(new_n252), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n407), .A2(new_n414), .A3(KEYINPUT85), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n419), .B1(new_n418), .B2(new_n420), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n496), .A3(new_n482), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(KEYINPUT6), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n235), .A2(new_n364), .A3(new_n204), .ZN(new_n499));
  OAI21_X1  g313(.A(G125), .B1(new_n271), .B2(new_n272), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G224), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(G953), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n501), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT6), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n505), .B(new_n483), .C1(new_n484), .C2(new_n490), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n498), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n482), .B(KEYINPUT8), .Z(new_n508));
  NAND2_X1  g322(.A1(new_n489), .A2(new_n442), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n496), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n503), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n499), .A2(new_n500), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n499), .B2(new_n500), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n515), .B2(new_n497), .ZN(new_n516));
  OAI21_X1  g330(.A(G210), .B1(G237), .B2(G902), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n507), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n507), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n481), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT89), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n507), .A2(new_n516), .ZN(new_n522));
  INV_X1    g336(.A(new_n517), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n507), .A2(new_n516), .A3(new_n517), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT89), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n481), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT9), .B(G234), .ZN(new_n529));
  OAI21_X1  g343(.A(G221), .B1(new_n529), .B2(G902), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n480), .A2(new_n521), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n370), .B1(new_n187), .B2(new_n352), .ZN(new_n532));
  INV_X1    g346(.A(G214), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n533), .A2(G237), .A3(G953), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT91), .B1(new_n535), .B2(new_n199), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G143), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n280), .A2(new_n281), .A3(G214), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n537), .B1(KEYINPUT90), .B2(G143), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n227), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g358(.A1(KEYINPUT18), .A2(G131), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n539), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n532), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n368), .A2(new_n369), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n548), .B2(new_n352), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n268), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n539), .A2(new_n227), .A3(new_n542), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n362), .B(new_n363), .C1(new_n553), .C2(new_n543), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n547), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G113), .B(G122), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(new_n400), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n358), .A2(new_n359), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n539), .A2(new_n542), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G131), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n552), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT93), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n543), .A2(new_n565), .A3(KEYINPUT17), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(new_n543), .B2(KEYINPUT17), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n560), .B(new_n564), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n557), .B(KEYINPUT92), .Z(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n547), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(G475), .A2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n573), .A2(KEYINPUT94), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT20), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(KEYINPUT94), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT95), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n572), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT20), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT95), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n571), .A2(new_n583), .A3(new_n578), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G475), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n568), .A2(new_n547), .A3(new_n569), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n557), .B1(new_n568), .B2(new_n547), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n302), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n586), .B1(new_n589), .B2(KEYINPUT96), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n568), .A2(new_n547), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n558), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n592), .B2(new_n570), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(G128), .B(G143), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n216), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n258), .A2(KEYINPUT14), .A3(G122), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n258), .A2(G122), .ZN(new_n601));
  INV_X1    g415(.A(G122), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G116), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(G107), .B(new_n600), .C1(new_n604), .C2(KEYINPUT14), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n416), .A2(new_n601), .A3(new_n603), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n599), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n409), .A2(new_n410), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n601), .A2(new_n603), .B1(new_n409), .B2(new_n410), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n604), .A2(new_n609), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n606), .A2(new_n613), .A3(KEYINPUT97), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n598), .B2(new_n216), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n338), .A2(G143), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n199), .A2(G128), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n615), .A2(new_n617), .A3(new_n618), .A4(new_n216), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n612), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(KEYINPUT13), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n618), .ZN(new_n623));
  INV_X1    g437(.A(new_n618), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n623), .A2(KEYINPUT98), .B1(KEYINPUT13), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(new_n626), .A3(new_n618), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n216), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n607), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n529), .A2(new_n390), .A3(G953), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n607), .B(new_n630), .C1(new_n621), .C2(new_n628), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n302), .ZN(new_n635));
  INV_X1    g449(.A(G478), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(KEYINPUT15), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n634), .B2(new_n302), .ZN(new_n640));
  AOI211_X1 g454(.A(KEYINPUT100), .B(G902), .C1(new_n632), .C2(new_n633), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n638), .B1(new_n642), .B2(new_n637), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n281), .A2(G952), .ZN(new_n644));
  INV_X1    g458(.A(G234), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n280), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n302), .B(new_n281), .C1(G234), .C2(G237), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT21), .B(G898), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n531), .A2(new_n597), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n397), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G101), .ZN(G3));
  NAND2_X1  g469(.A1(new_n299), .A2(new_n302), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n656), .A2(G472), .B1(new_n304), .B2(new_n299), .ZN(new_n657));
  INV_X1    g471(.A(new_n396), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n530), .A4(new_n480), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT101), .ZN(new_n660));
  INV_X1    g474(.A(new_n520), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n651), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n634), .B(KEYINPUT33), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(G478), .A3(new_n302), .ZN(new_n664));
  INV_X1    g478(.A(new_n642), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n664), .B1(new_n665), .B2(G478), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n597), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT34), .B(G104), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  INV_X1    g485(.A(new_n643), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n575), .B1(new_n571), .B2(new_n572), .ZN(new_n673));
  AOI211_X1 g487(.A(KEYINPUT20), .B(new_n573), .C1(new_n559), .C2(new_n570), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n590), .A2(KEYINPUT102), .A3(new_n595), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT102), .B1(new_n590), .B2(new_n595), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n672), .B(new_n676), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n662), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n660), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT35), .B(G107), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  NOR2_X1   g498(.A1(new_n380), .A2(KEYINPUT36), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n376), .B(new_n685), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n389), .A2(new_n391), .B1(new_n394), .B2(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n597), .A3(new_n652), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n657), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n531), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT37), .B(G110), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  NOR2_X1   g506(.A1(new_n520), .A2(new_n687), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n694));
  OAI21_X1  g508(.A(G475), .B1(new_n593), .B2(new_n594), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n589), .A2(KEYINPUT96), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n675), .B(new_n643), .C1(new_n697), .C2(new_n677), .ZN(new_n698));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n647), .B1(new_n648), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n693), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n480), .A2(new_n530), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n335), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n329), .A2(new_n311), .A3(new_n312), .A4(new_n321), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n705), .B1(new_n706), .B2(KEYINPUT75), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n301), .B1(new_n707), .B2(new_n330), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n704), .B(KEYINPUT103), .C1(new_n307), .C2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n680), .A2(new_n700), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n530), .A3(new_n480), .A4(new_n693), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n710), .B1(new_n337), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G128), .ZN(G30));
  AND2_X1   g529(.A1(new_n480), .A2(new_n530), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n700), .B(KEYINPUT39), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT40), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n332), .A2(new_n333), .ZN(new_n721));
  AOI21_X1  g535(.A(G902), .B1(new_n721), .B2(new_n285), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n308), .A2(new_n286), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n301), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n306), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n518), .A2(new_n519), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT38), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n686), .A2(new_n394), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n392), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n597), .A2(new_n672), .A3(new_n481), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n720), .A2(new_n729), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  NAND2_X1  g551(.A1(new_n336), .A2(G472), .ZN(new_n738));
  INV_X1    g552(.A(new_n307), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n597), .A2(new_n666), .A3(new_n701), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n703), .A2(new_n520), .A3(new_n687), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G146), .ZN(G48));
  INV_X1    g558(.A(new_n530), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n467), .A2(new_n302), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G469), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  AOI21_X1  g562(.A(G902), .B1(new_n462), .B2(new_n466), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(new_n468), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n749), .A2(KEYINPUT105), .A3(new_n468), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n745), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n397), .A2(new_n668), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  NAND4_X1  g571(.A1(new_n740), .A2(new_n658), .A3(new_n681), .A4(new_n754), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G116), .ZN(G18));
  AOI211_X1 g573(.A(new_n745), .B(new_n520), .C1(new_n751), .C2(new_n753), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n740), .A2(new_n688), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G119), .ZN(G21));
  NAND2_X1  g576(.A1(new_n751), .A2(new_n753), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n585), .A2(new_n596), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n520), .A2(new_n764), .A3(new_n650), .A4(new_n643), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n530), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n286), .B1(new_n334), .B2(new_n290), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT106), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n235), .A2(new_n236), .A3(new_n204), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n236), .B1(new_n235), .B2(new_n204), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n770), .A2(new_n771), .A3(new_n231), .ZN(new_n772));
  INV_X1    g586(.A(new_n250), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n264), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n289), .B1(new_n774), .B2(new_n279), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n285), .B1(new_n775), .B2(new_n291), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT106), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n288), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n769), .A2(new_n778), .A3(new_n298), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n304), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n656), .A2(G472), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n658), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n766), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n602), .ZN(G24));
  INV_X1    g598(.A(new_n741), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n780), .A2(new_n785), .A3(new_n781), .A4(new_n733), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n760), .A2(new_n787), .A3(KEYINPUT107), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT107), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n749), .A2(new_n468), .ZN(new_n790));
  AOI211_X1 g604(.A(G469), .B(G902), .C1(new_n462), .C2(new_n466), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n791), .A3(new_n748), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n530), .B(new_n661), .C1(new_n792), .C2(new_n752), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n789), .B1(new_n793), .B2(new_n786), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G125), .ZN(G27));
  INV_X1    g610(.A(KEYINPUT42), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  INV_X1    g612(.A(new_n481), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n526), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT108), .B1(new_n730), .B2(new_n481), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n716), .A3(new_n785), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT109), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n797), .B(new_n804), .C1(new_n397), .C2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n658), .B1(new_n708), .B2(new_n307), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT109), .B(KEYINPUT42), .C1(new_n807), .C2(new_n803), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n227), .ZN(G33));
  OAI21_X1  g624(.A(new_n798), .B1(new_n526), .B2(new_n799), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n730), .A2(KEYINPUT108), .A3(new_n481), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n480), .A3(new_n812), .A4(new_n530), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n680), .A3(new_n700), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n397), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G134), .ZN(G36));
  NAND2_X1  g630(.A1(new_n764), .A2(new_n666), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT43), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n817), .B(KEYINPUT43), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT111), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n657), .A2(new_n687), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT44), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n802), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n828), .A2(new_n829), .B1(new_n826), .B2(new_n825), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n471), .A2(new_n476), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT45), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n471), .A2(KEYINPUT45), .A3(new_n476), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(G469), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n479), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT46), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n478), .B1(new_n837), .B2(new_n838), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n469), .B1(new_n843), .B2(KEYINPUT46), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n530), .B(new_n717), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n830), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G137), .ZN(G39));
  INV_X1    g662(.A(new_n802), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n740), .A2(new_n849), .A3(new_n658), .A4(new_n741), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n530), .B1(new_n842), .B2(new_n844), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT47), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(KEYINPUT47), .B(new_n530), .C1(new_n842), .C2(new_n844), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n850), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(KEYINPUT113), .B(G140), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(G42));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n734), .A2(new_n730), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n733), .A2(new_n700), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n530), .A4(new_n480), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n727), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n740), .B2(new_n742), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n714), .A2(new_n795), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT52), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n714), .A2(new_n795), .A3(new_n864), .A4(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n867), .B1(new_n866), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n733), .A2(new_n643), .A3(new_n701), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n813), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n397), .A2(new_n814), .B1(new_n875), .B2(new_n740), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n780), .A2(new_n781), .A3(new_n733), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT115), .B1(new_n803), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n813), .A2(new_n741), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n880));
  INV_X1    g694(.A(new_n877), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  AND4_X1   g697(.A1(new_n808), .A2(new_n806), .A3(new_n876), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n755), .A2(new_n758), .A3(new_n761), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n672), .A2(new_n585), .A3(new_n596), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n667), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n521), .A3(new_n528), .A4(new_n651), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n659), .A2(new_n888), .B1(new_n531), .B2(new_n689), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n783), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n654), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n884), .A2(KEYINPUT116), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n806), .A2(new_n876), .A3(new_n808), .A4(new_n883), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n397), .B(new_n754), .C1(new_n668), .C2(new_n681), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n654), .A3(new_n761), .A4(new_n890), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n859), .B1(new_n872), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n866), .A2(new_n869), .ZN(new_n901));
  AOI211_X1 g715(.A(KEYINPUT53), .B(new_n901), .C1(new_n893), .C2(new_n898), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n884), .A2(KEYINPUT53), .A3(new_n892), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n901), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n713), .A2(new_n709), .B1(new_n788), .B2(new_n794), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n868), .B1(new_n907), .B2(new_n864), .ZN(new_n908));
  INV_X1    g722(.A(new_n869), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT117), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT116), .B1(new_n884), .B2(new_n892), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n895), .A2(new_n897), .A3(new_n894), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  AOI211_X1 g728(.A(KEYINPUT54), .B(new_n906), .C1(new_n914), .C2(new_n859), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n904), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n851), .A2(new_n852), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n763), .B(KEYINPUT114), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n745), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n854), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT119), .B1(new_n822), .B2(new_n646), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n819), .A2(new_n922), .A3(new_n647), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n782), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n849), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n754), .A2(new_n799), .A3(new_n731), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT50), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n729), .A2(new_n396), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n754), .A2(new_n802), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n932), .A2(new_n647), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n597), .A2(new_n666), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n924), .A2(new_n933), .ZN(new_n936));
  AOI22_X1  g750(.A1(new_n934), .A2(new_n935), .B1(new_n936), .B2(new_n881), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n928), .A2(KEYINPUT51), .A3(new_n931), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n397), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT48), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n644), .B1(new_n926), .B2(new_n793), .ZN(new_n941));
  INV_X1    g755(.A(new_n667), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n934), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT120), .B1(new_n853), .B2(new_n855), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n917), .A2(new_n946), .A3(new_n854), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n947), .A3(new_n919), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n927), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n931), .A2(new_n937), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n944), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n916), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(G952), .B2(G953), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n918), .B(KEYINPUT49), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n817), .A2(new_n745), .A3(new_n799), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n956), .A2(new_n731), .A3(new_n932), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(G75));
  INV_X1    g773(.A(KEYINPUT56), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n906), .B1(new_n914), .B2(new_n859), .ZN(new_n961));
  NAND2_X1  g775(.A1(G210), .A2(G902), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n498), .A2(new_n506), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n504), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT55), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n960), .B(new_n968), .C1(new_n961), .C2(new_n962), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n281), .A2(G952), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT121), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n967), .A2(KEYINPUT121), .A3(new_n969), .A4(new_n971), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G51));
  NOR3_X1   g790(.A1(new_n961), .A2(new_n302), .A3(new_n839), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT122), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n478), .B(KEYINPUT57), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n914), .A2(new_n859), .ZN(new_n980));
  INV_X1    g794(.A(new_n906), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n903), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n979), .B1(new_n982), .B2(new_n915), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n467), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n970), .B1(new_n978), .B2(new_n984), .ZN(G54));
  NOR2_X1   g799(.A1(new_n961), .A2(new_n302), .ZN(new_n986));
  AND2_X1   g800(.A1(KEYINPUT58), .A2(G475), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n986), .A2(new_n571), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n571), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n988), .A2(new_n989), .A3(new_n970), .ZN(G60));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n663), .B(KEYINPUT123), .ZN(new_n992));
  NAND2_X1  g806(.A1(G478), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT59), .Z(new_n994));
  NOR2_X1   g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT53), .B1(new_n872), .B2(new_n899), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT54), .B1(new_n997), .B2(new_n906), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n980), .A2(new_n903), .A3(new_n981), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n991), .B1(new_n1000), .B2(new_n970), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n995), .B1(new_n982), .B2(new_n915), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1002), .A2(KEYINPUT124), .A3(new_n971), .ZN(new_n1003));
  INV_X1    g817(.A(new_n994), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n904), .B2(new_n915), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n992), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1001), .A2(new_n1003), .A3(new_n1006), .ZN(G63));
  NAND2_X1  g821(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G217), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT60), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n393), .B1(new_n961), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n970), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1010), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n686), .B(new_n1015), .C1(new_n997), .C2(new_n906), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1008), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  AND4_X1   g831(.A1(new_n1008), .A2(new_n1011), .A3(new_n1016), .A4(new_n1013), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(G66));
  OAI21_X1  g833(.A(G953), .B1(new_n649), .B2(new_n502), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(new_n892), .B2(G953), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n964), .B1(G898), .B2(new_n281), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1021), .B(new_n1022), .ZN(G69));
  AOI21_X1  g837(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n251), .A2(new_n277), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(new_n550), .ZN(new_n1026));
  NAND2_X1  g840(.A1(G900), .A2(G953), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n807), .A2(new_n730), .A3(new_n734), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n846), .B1(new_n830), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n907), .A2(new_n743), .ZN(new_n1030));
  AOI211_X1 g844(.A(new_n809), .B(new_n1030), .C1(new_n397), .C2(new_n814), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1029), .A2(new_n856), .A3(new_n1031), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1026), .B(new_n1027), .C1(new_n1032), .C2(G953), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1024), .B1(new_n1033), .B2(KEYINPUT126), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n736), .A2(new_n907), .A3(new_n743), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT62), .Z(new_n1036));
  INV_X1    g850(.A(new_n718), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n397), .A2(new_n1037), .A3(new_n802), .A4(new_n887), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n1036), .A2(new_n847), .A3(new_n856), .A4(new_n1038), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1039), .A2(new_n281), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1033), .B1(new_n1040), .B2(new_n1026), .ZN(new_n1041));
  AND2_X1   g855(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1042), .A2(new_n1043), .ZN(G72));
  NAND2_X1  g858(.A1(G472), .A2(G902), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1045), .B(KEYINPUT63), .Z(new_n1046));
  OAI21_X1  g860(.A(new_n1046), .B1(new_n1039), .B2(new_n897), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1047), .A2(new_n286), .A3(new_n308), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1046), .B1(new_n1032), .B2(new_n897), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n308), .A2(new_n286), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1050), .B(KEYINPUT127), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1048), .A2(new_n971), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n278), .A2(new_n287), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1046), .B1(new_n313), .B2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g869(.A1(new_n900), .A2(new_n902), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n1053), .A2(new_n1056), .ZN(G57));
endmodule


