//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n204), .A2(G1gat), .ZN(new_n208));
  OAI21_X1  g007(.A(G8gat), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n210), .C1(G1gat), .C2(new_n204), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT88), .B(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G43gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n214), .B(new_n215), .C1(new_n219), .C2(KEYINPUT89), .ZN(new_n220));
  NOR2_X1   g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT15), .ZN(new_n224));
  NAND2_X1  g023(.A1(G29gat), .A2(G36gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT90), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n220), .A2(new_n223), .A3(new_n224), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n225), .ZN(new_n229));
  INV_X1    g028(.A(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n212), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n232), .A2(new_n235), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n203), .B(new_n233), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT91), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n202), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n228), .A2(new_n231), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n233), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n203), .B(KEYINPUT13), .Z(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n239), .A2(new_n240), .A3(new_n202), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G197gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT11), .B(G169gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT12), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n250), .A2(new_n241), .A3(new_n248), .ZN(new_n259));
  INV_X1    g058(.A(new_n257), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT82), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT31), .B(G50gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n267), .B(KEYINPUT83), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G228gat), .ZN(new_n270));
  INV_X1    g069(.A(G233gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G197gat), .B(G204gat), .ZN(new_n277));
  INV_X1    g076(.A(G211gat), .ZN(new_n278));
  INV_X1    g077(.A(G218gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n277), .B1(KEYINPUT22), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n276), .B(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n273), .B1(new_n282), .B2(KEYINPUT29), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(G155gat), .B2(G162gat), .ZN(new_n286));
  AND2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n284), .A2(new_n286), .B1(KEYINPUT76), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G155gat), .B(G162gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI221_X1 g090(.A(new_n289), .B1(new_n287), .B2(KEYINPUT76), .C1(new_n284), .C2(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(KEYINPUT77), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT78), .ZN(new_n299));
  INV_X1    g098(.A(new_n293), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(KEYINPUT3), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(KEYINPUT78), .A3(new_n273), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT29), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n282), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n272), .B(new_n298), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G22gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n274), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT29), .B1(new_n281), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n307), .B2(new_n281), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n293), .B1(new_n309), .B2(new_n273), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n301), .A2(new_n302), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n313), .B2(new_n282), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n305), .B(new_n306), .C1(new_n314), .C2(new_n272), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n303), .A2(new_n304), .ZN(new_n317));
  OAI22_X1  g116(.A1(new_n317), .A2(new_n310), .B1(new_n270), .B2(new_n271), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n306), .B1(new_n318), .B2(new_n305), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n269), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT84), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n305), .B1(new_n314), .B2(new_n272), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G22gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n315), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT84), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n269), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n315), .A2(new_n267), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n319), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(KEYINPUT85), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n321), .A2(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT27), .B(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT28), .ZN(new_n335));
  NOR2_X1   g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n336), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(KEYINPUT26), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(G169gat), .B2(G176gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n339), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n344), .A2(KEYINPUT66), .A3(new_n346), .A4(new_n339), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT24), .B1(new_n351), .B2(new_n333), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT24), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(G183gat), .A3(G190gat), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT65), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n349), .B(new_n350), .C1(new_n355), .C2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n352), .B2(new_n354), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n361), .A2(new_n347), .A3(new_n359), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n343), .A2(new_n364), .A3(KEYINPUT73), .ZN(new_n365));
  INV_X1    g164(.A(G226gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(new_n271), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(KEYINPUT29), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n362), .B1(new_n358), .B2(new_n359), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(new_n342), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n365), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n370), .A2(KEYINPUT67), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT67), .ZN(new_n374));
  AOI211_X1 g173(.A(new_n374), .B(new_n362), .C1(new_n358), .C2(new_n359), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n367), .B(new_n343), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n304), .ZN(new_n378));
  INV_X1    g177(.A(new_n371), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n370), .A2(new_n342), .A3(new_n369), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n367), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n343), .B1(new_n373), .B2(new_n375), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n368), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n383), .A3(new_n282), .ZN(new_n384));
  XNOR2_X1  g183(.A(G8gat), .B(G36gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  NAND3_X1  g186(.A1(new_n378), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(new_n384), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT74), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT74), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n378), .A2(new_n384), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n387), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT30), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n378), .A2(new_n384), .A3(KEYINPUT30), .A4(new_n387), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT75), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT40), .ZN(new_n400));
  XNOR2_X1  g199(.A(G113gat), .B(G120gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(KEYINPUT1), .ZN(new_n402));
  XOR2_X1   g201(.A(G127gat), .B(G134gat), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n293), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(KEYINPUT4), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n404), .B1(new_n297), .B2(KEYINPUT3), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n311), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n410), .B2(new_n311), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT39), .ZN(new_n416));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G1gat), .B(G29gat), .Z(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n405), .ZN(new_n426));
  INV_X1    g225(.A(new_n404), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(new_n297), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n417), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT39), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n415), .B2(new_n418), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n400), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n409), .B(new_n433), .C1(new_n413), .C2(new_n414), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n406), .A2(KEYINPUT80), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n404), .A2(new_n293), .A3(KEYINPUT80), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n408), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n417), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n410), .A2(new_n311), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT79), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n441), .B2(new_n412), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT5), .B1(new_n428), .B2(new_n417), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n434), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n424), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n441), .A2(new_n412), .B1(new_n407), .B2(new_n408), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT39), .B(new_n429), .C1(new_n447), .C2(new_n417), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n448), .A2(KEYINPUT40), .A3(new_n419), .A4(new_n424), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n432), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n331), .B1(new_n399), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  INV_X1    g252(.A(new_n368), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n364), .A2(new_n374), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n370), .A2(KEYINPUT67), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n457), .B2(new_n343), .ZN(new_n458));
  INV_X1    g257(.A(new_n367), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n365), .B2(new_n371), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n304), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n461), .A2(KEYINPUT86), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n377), .A2(new_n304), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n461), .B2(KEYINPUT86), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n453), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n378), .A2(new_n384), .A3(new_n453), .ZN(new_n466));
  INV_X1    g265(.A(new_n387), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n452), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n452), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n378), .A2(new_n384), .A3(new_n391), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n391), .B1(new_n378), .B2(new_n384), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n434), .B(new_n424), .C1(new_n442), .C2(new_n443), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n446), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n445), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n481), .A3(new_n388), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n395), .A3(new_n398), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n451), .A2(new_n482), .B1(new_n483), .B2(new_n331), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G43gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT69), .ZN(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT64), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n404), .B1(new_n457), .B2(new_n343), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n382), .A2(new_n427), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT68), .ZN(new_n496));
  INV_X1    g295(.A(new_n490), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n457), .A2(new_n404), .A3(new_n343), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n382), .A2(new_n427), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT32), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n493), .A2(KEYINPUT68), .A3(KEYINPUT32), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n495), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n488), .A2(new_n494), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n493), .A2(KEYINPUT32), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n493), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n498), .A2(new_n499), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n489), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n516), .A2(KEYINPUT34), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n512), .A2(KEYINPUT34), .A3(new_n490), .ZN(new_n518));
  OAI22_X1  g317(.A1(new_n505), .A2(new_n511), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n518), .B1(new_n516), .B2(KEYINPUT34), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n521), .A2(new_n504), .A3(new_n509), .A4(new_n510), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n519), .B2(new_n522), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n484), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n319), .A2(new_n328), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n330), .A2(new_n527), .A3(new_n315), .A4(new_n267), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n325), .B1(new_n324), .B2(new_n269), .ZN(new_n529));
  AOI211_X1 g328(.A(KEYINPUT84), .B(new_n268), .C1(new_n323), .C2(new_n315), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n531), .A2(new_n519), .A3(new_n522), .ZN(new_n532));
  INV_X1    g331(.A(new_n483), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n519), .A3(new_n522), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT35), .B1(new_n536), .B2(new_n483), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n263), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n540));
  OR2_X1    g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT94), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544));
  AND2_X1   g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(KEYINPUT8), .ZN(new_n549));
  OR2_X1    g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G85gat), .A2(G92gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n548), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n549), .A2(new_n554), .A3(new_n550), .A4(new_n555), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(new_n547), .A3(new_n543), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n236), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n540), .B1(new_n561), .B2(new_n238), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n242), .A2(KEYINPUT17), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(KEYINPUT95), .A3(new_n236), .A4(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT41), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n242), .B2(new_n560), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n565), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n568), .A2(KEYINPUT41), .ZN(new_n574));
  XNOR2_X1  g373(.A(G134gat), .B(G162gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n567), .B1(new_n565), .B2(new_n571), .ZN(new_n578));
  OR3_X1    g377(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n573), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(G57gat), .A2(G64gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G57gat), .A2(G64gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G71gat), .B(G78gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(G71gat), .B2(G78gat), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n587), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n234), .B1(new_n594), .B2(new_n593), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT93), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n599), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n581), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n558), .B1(new_n547), .B2(new_n543), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n609));
  OAI22_X1  g408(.A1(new_n608), .A2(new_n609), .B1(new_n591), .B2(new_n592), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n548), .B(new_n558), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n557), .A2(KEYINPUT96), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n590), .ZN(new_n614));
  INV_X1    g413(.A(new_n588), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n560), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G120gat), .B(G148gat), .Z(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n560), .A2(new_n593), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n619), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(new_n628), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n622), .B(new_n627), .C1(new_n631), .C2(new_n621), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT99), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT10), .B1(new_n612), .B2(new_n619), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n620), .B1(new_n634), .B2(new_n629), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n635), .A2(new_n636), .A3(new_n622), .A4(new_n627), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n627), .B1(new_n635), .B2(new_n622), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT100), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642));
  AOI211_X1 g441(.A(new_n642), .B(new_n639), .C1(new_n633), .C2(new_n637), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n607), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n539), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n481), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g448(.A(new_n210), .B1(new_n647), .B2(new_n399), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT30), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n397), .B1(new_n652), .B2(new_n388), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT16), .B(G8gat), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n646), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(KEYINPUT42), .B2(new_n655), .ZN(G1325gat));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n523), .B2(new_n524), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n509), .A2(new_n510), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n521), .B1(new_n660), .B2(new_n504), .ZN(new_n661));
  INV_X1    g460(.A(new_n522), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT36), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(KEYINPUT101), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n646), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n661), .A2(new_n662), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(G15gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n667), .B1(new_n646), .B2(new_n670), .ZN(G1326gat));
  NOR2_X1   g470(.A1(new_n646), .A2(new_n531), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT43), .B(G22gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n581), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n526), .B2(new_n538), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n579), .A2(new_n580), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n483), .A2(new_n331), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n432), .A2(new_n449), .A3(new_n446), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n531), .B1(new_n653), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n478), .A2(new_n479), .A3(new_n388), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n469), .B2(new_n474), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n665), .B2(new_n659), .ZN(new_n686));
  INV_X1    g485(.A(new_n538), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n679), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n678), .B1(new_n688), .B2(new_n675), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n644), .B(KEYINPUT102), .Z(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(new_n263), .A3(new_n606), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT103), .B1(new_n692), .B2(new_n480), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n689), .A2(new_n694), .A3(new_n481), .A4(new_n691), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(G29gat), .A3(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n644), .A2(new_n606), .A3(new_n581), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n480), .A2(G29gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n539), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n696), .A2(new_n700), .ZN(G1328gat));
  OAI21_X1  g500(.A(G36gat), .B1(new_n692), .B2(new_n653), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n653), .A2(G36gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n539), .A2(new_n697), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT46), .Z(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(G1329gat));
  NOR2_X1   g505(.A1(new_n666), .A2(new_n213), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n689), .A2(new_n691), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n539), .A2(new_n668), .A3(new_n697), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n709), .A2(new_n213), .B1(KEYINPUT104), .B2(KEYINPUT47), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g510(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1330gat));
  NAND2_X1  g512(.A1(new_n331), .A2(G50gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n689), .A2(new_n691), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n539), .A2(new_n331), .A3(new_n697), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n717), .A2(new_n216), .B1(new_n718), .B2(KEYINPUT48), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n718), .A2(KEYINPUT48), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1331gat));
  NOR3_X1   g521(.A1(new_n523), .A2(new_n524), .A3(new_n658), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT101), .B1(new_n663), .B2(new_n664), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n484), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n538), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n607), .A2(new_n262), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n690), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT106), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n481), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g532(.A(new_n653), .B(new_n730), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n666), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n726), .A2(new_n729), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT107), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT108), .B1(new_n730), .B2(new_n669), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n729), .A3(new_n742), .A4(new_n668), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n737), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT50), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n740), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n331), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n526), .A2(new_n538), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n676), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n262), .A2(new_n606), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT109), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(new_n644), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n581), .B1(new_n725), .B2(new_n538), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n753), .B(new_n756), .C1(new_n757), .C2(KEYINPUT44), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n480), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n726), .A2(new_n679), .A3(new_n755), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n757), .A2(KEYINPUT51), .A3(new_n755), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n644), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n766), .A2(new_n480), .A3(G85gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n759), .B1(new_n765), .B2(new_n767), .ZN(G1336gat));
  OAI21_X1  g567(.A(KEYINPUT110), .B1(new_n758), .B2(new_n653), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n689), .A2(new_n770), .A3(new_n399), .A4(new_n756), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n771), .A3(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(new_n690), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n773), .A2(G92gat), .A3(new_n653), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n764), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G92gat), .B1(new_n758), .B2(new_n653), .ZN(new_n777));
  AND4_X1   g576(.A1(KEYINPUT51), .A2(new_n726), .A3(new_n679), .A4(new_n755), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n757), .B2(new_n755), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT52), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n776), .A2(new_n782), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n758), .B2(new_n666), .ZN(new_n784));
  OR3_X1    g583(.A1(new_n669), .A2(G99gat), .A3(new_n766), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n765), .B2(new_n785), .ZN(G1338gat));
  OAI21_X1  g585(.A(G106gat), .B1(new_n758), .B2(new_n531), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n773), .A2(G106gat), .A3(new_n531), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n778), .B2(new_n779), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n787), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n727), .B2(new_n766), .ZN(new_n797));
  NOR4_X1   g596(.A1(new_n607), .A2(new_n644), .A3(KEYINPUT112), .A4(new_n262), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n631), .A2(new_n621), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n800), .A2(KEYINPUT54), .A3(new_n635), .ZN(new_n801));
  INV_X1    g600(.A(new_n627), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n635), .B2(KEYINPUT54), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n804), .A2(KEYINPUT55), .B1(new_n633), .B2(new_n637), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n801), .B2(new_n803), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n262), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n256), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n237), .A2(new_n238), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n234), .A2(new_n242), .ZN(new_n811));
  OAI211_X1 g610(.A(G229gat), .B(G233gat), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n245), .A2(new_n247), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n809), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n259), .B2(new_n260), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n641), .B2(new_n643), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n808), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n581), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n679), .A2(new_n815), .A3(new_n807), .A4(new_n805), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n606), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n481), .B(new_n532), .C1(new_n799), .C2(new_n820), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n399), .B1(new_n821), .B2(KEYINPUT114), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n263), .A2(G113gat), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n824), .B(KEYINPUT115), .Z(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n821), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n653), .A3(new_n262), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT113), .B1(new_n828), .B2(G113gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(G1340gat));
  NOR2_X1   g630(.A1(new_n766), .A2(G120gat), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n822), .A2(new_n823), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n827), .A2(new_n653), .A3(new_n690), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n835), .A2(new_n836), .A3(G120gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n835), .B2(G120gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(G1341gat));
  INV_X1    g638(.A(new_n606), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(G127gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n822), .A2(new_n823), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(G127gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n821), .A2(new_n399), .A3(new_n840), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(G1342gat));
  NOR2_X1   g644(.A1(new_n581), .A2(G134gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n822), .A2(new_n823), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n827), .A2(new_n653), .A3(new_n679), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G134gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT118), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n848), .A2(new_n850), .A3(new_n851), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n399), .A2(new_n480), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n666), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n799), .ZN(new_n859));
  INV_X1    g658(.A(new_n820), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n531), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n262), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(G141gat), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  AND4_X1   g664(.A1(new_n679), .A2(new_n815), .A3(new_n807), .A4(new_n805), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n816), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n815), .B(KEYINPUT119), .C1(new_n641), .C2(new_n643), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n807), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT120), .B(new_n806), .C1(new_n801), .C2(new_n803), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n262), .A2(new_n805), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n866), .B1(new_n874), .B2(new_n581), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n875), .A2(KEYINPUT121), .A3(new_n606), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(new_n875), .B2(new_n606), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n859), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n865), .B1(new_n878), .B2(new_n331), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n865), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n858), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n263), .A2(new_n863), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n864), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT58), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  NOR4_X1   g686(.A1(new_n879), .A2(new_n881), .A3(new_n863), .A4(new_n263), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT122), .B(new_n887), .C1(new_n888), .C2(new_n864), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1344gat));
  AND2_X1   g689(.A1(new_n858), .A2(new_n861), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n644), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT57), .B(new_n331), .C1(new_n799), .C2(new_n820), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n727), .A2(new_n766), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n875), .B2(new_n606), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n897), .B2(new_n331), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n898), .B2(KEYINPUT124), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900));
  AOI211_X1 g699(.A(new_n900), .B(KEYINPUT57), .C1(new_n897), .C2(new_n331), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n858), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n903), .A2(KEYINPUT123), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n766), .B1(new_n903), .B2(KEYINPUT123), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n894), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  AOI211_X1 g706(.A(KEYINPUT59), .B(new_n892), .C1(new_n882), .C2(new_n644), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n893), .B1(new_n907), .B2(new_n908), .ZN(G1345gat));
  AOI21_X1  g708(.A(G155gat), .B1(new_n891), .B2(new_n606), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n606), .A2(G155gat), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT125), .Z(new_n912));
  AOI21_X1  g711(.A(new_n910), .B1(new_n882), .B2(new_n912), .ZN(G1346gat));
  INV_X1    g712(.A(G162gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n891), .A2(new_n914), .A3(new_n679), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n879), .A2(new_n881), .A3(new_n581), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n914), .ZN(G1347gat));
  AOI21_X1  g716(.A(new_n536), .B1(new_n859), .B2(new_n860), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n481), .A2(new_n653), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n262), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(G169gat), .ZN(G1348gat));
  OR3_X1    g722(.A1(new_n920), .A2(G176gat), .A3(new_n766), .ZN(new_n924));
  OAI21_X1  g723(.A(G176gat), .B1(new_n920), .B2(new_n773), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(new_n351), .B1(new_n920), .B2(new_n840), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n921), .A2(new_n606), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n332), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT60), .Z(G1350gat));
  NOR2_X1   g729(.A1(new_n920), .A2(new_n581), .ZN(new_n931));
  NAND2_X1  g730(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g732(.A(KEYINPUT61), .B(G190gat), .Z(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n931), .B2(new_n934), .ZN(G1351gat));
  AND2_X1   g734(.A1(new_n666), .A2(new_n919), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n902), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(G197gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(new_n263), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n936), .A2(new_n861), .ZN(new_n940));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n262), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n939), .A2(new_n941), .ZN(G1352gat));
  NOR2_X1   g741(.A1(new_n766), .A2(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n936), .A2(new_n861), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n945), .A2(KEYINPUT62), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT62), .B1(new_n945), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n937), .B2(new_n773), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1353gat));
  OAI211_X1 g750(.A(new_n606), .B(new_n936), .C1(new_n899), .C2(new_n901), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G211gat), .ZN(new_n953));
  NOR2_X1   g752(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n952), .B(G211gat), .C1(KEYINPUT127), .C2(KEYINPUT63), .ZN(new_n956));
  NAND2_X1  g755(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n278), .A3(new_n606), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1354gat));
  OAI21_X1  g759(.A(G218gat), .B1(new_n937), .B2(new_n581), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n940), .A2(new_n279), .A3(new_n679), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1355gat));
endmodule


