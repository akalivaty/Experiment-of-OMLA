//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n597,
    new_n599, new_n600, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n451), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n467), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n460), .B1(new_n476), .B2(new_n477), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n474), .B(new_n480), .C1(G124), .C2(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n483), .A2(KEYINPUT68), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n481), .A2(G126), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n460), .A2(G138), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n476), .B2(new_n477), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n460), .A2(G138), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(new_n493), .C1(new_n462), .C2(new_n461), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n485), .B(new_n490), .C1(new_n494), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n506), .A2(new_n509), .ZN(G303));
  INV_X1    g085(.A(G303), .ZN(G166));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(G51), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n504), .B2(new_n514), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT5), .B(G543), .Z(new_n516));
  NAND2_X1  g091(.A1(new_n500), .A2(G89), .ZN(new_n517));
  NAND2_X1  g092(.A1(G63), .A2(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(G168));
  INV_X1    g095(.A(G90), .ZN(new_n521));
  INV_X1    g096(.A(G52), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n502), .A2(new_n521), .B1(new_n504), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n508), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n523), .A2(new_n525), .ZN(G301));
  INV_X1    g101(.A(G301), .ZN(G171));
  AOI22_X1  g102(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n508), .ZN(new_n529));
  INV_X1    g104(.A(new_n502), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G81), .ZN(new_n531));
  INV_X1    g106(.A(new_n504), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G43), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n534), .B1(new_n531), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g115(.A(KEYINPUT70), .B(KEYINPUT8), .Z(new_n541));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(G188));
  INV_X1    g119(.A(G53), .ZN(new_n545));
  OR3_X1    g120(.A1(new_n504), .A2(KEYINPUT9), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT9), .B1(new_n504), .B2(new_n545), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G78), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n516), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G651), .B1(new_n530), .B2(G91), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G299));
  INV_X1    g128(.A(G168), .ZN(G286));
  NAND2_X1  g129(.A1(new_n530), .A2(G87), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n532), .A2(G49), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(G288));
  NAND2_X1  g133(.A1(new_n530), .A2(G86), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n532), .A2(G48), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT71), .ZN(new_n561));
  NAND2_X1  g136(.A1(G73), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G61), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n516), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n561), .B1(new_n564), .B2(G651), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n566), .A2(KEYINPUT71), .A3(new_n508), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n559), .B(new_n560), .C1(new_n565), .C2(new_n567), .ZN(G305));
  AOI22_X1  g143(.A1(G85), .A2(new_n530), .B1(new_n532), .B2(G47), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n508), .B2(new_n570), .ZN(G290));
  INV_X1    g146(.A(G868), .ZN(new_n572));
  NOR2_X1   g147(.A1(G301), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT10), .ZN(new_n575));
  INV_X1    g150(.A(G92), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n502), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n574), .A2(new_n577), .B1(G54), .B2(new_n532), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G66), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n516), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT73), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n584), .A2(new_n585), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n588), .A2(new_n589), .A3(new_n578), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n573), .B1(new_n591), .B2(new_n572), .ZN(G284));
  AOI21_X1  g167(.A(new_n573), .B1(new_n591), .B2(new_n572), .ZN(G321));
  NAND2_X1  g168(.A1(G299), .A2(new_n572), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n572), .B2(G168), .ZN(G297));
  OAI21_X1  g170(.A(new_n594), .B1(new_n572), .B2(G168), .ZN(G280));
  XNOR2_X1  g171(.A(KEYINPUT74), .B(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n591), .B1(G860), .B2(new_n597), .ZN(G148));
  NAND2_X1  g173(.A1(new_n537), .A2(new_n572), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n591), .A2(new_n597), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n572), .ZN(G323));
  XOR2_X1   g176(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n602));
  XNOR2_X1  g177(.A(G323), .B(new_n602), .ZN(G282));
  NAND2_X1  g178(.A1(new_n476), .A2(new_n477), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(new_n468), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G2100), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT77), .ZN(new_n610));
  AOI22_X1  g185(.A1(G123), .A2(new_n481), .B1(new_n478), .B2(G135), .ZN(new_n611));
  NOR3_X1   g186(.A1(new_n460), .A2(KEYINPUT78), .A3(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT78), .B1(new_n460), .B2(G111), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n613), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2096), .Z(new_n616));
  OAI211_X1 g191(.A(new_n610), .B(new_n616), .C1(G2100), .C2(new_n608), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT79), .Z(G156));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT81), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2427), .B(G2430), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(G14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT82), .ZN(G401));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT83), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT17), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT84), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n643), .B(new_n645), .C1(new_n642), .C2(new_n638), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n638), .A2(new_n640), .A3(new_n644), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n641), .A2(new_n644), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n648), .C1(new_n639), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2096), .B(G2100), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1981), .B(G1986), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G305), .ZN(new_n673));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(G6), .B2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT32), .B(G1981), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(G22), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n674), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1971), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n674), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(G288), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n674), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT33), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR4_X1   g263(.A1(new_n679), .A2(new_n680), .A3(new_n683), .A4(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n674), .A2(G24), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT90), .Z(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G290), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G25), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n478), .A2(G131), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT88), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n481), .A2(G119), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n460), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT89), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n698), .B1(new_n705), .B2(new_n697), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n696), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n706), .B2(new_n708), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n691), .A2(new_n692), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT36), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n697), .A2(G32), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n481), .A2(G129), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT98), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT99), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT26), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n715), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n713), .B1(new_n720), .B2(G29), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT100), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n674), .A2(G5), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G171), .B2(new_n674), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT103), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n729));
  INV_X1    g304(.A(G34), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n697), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT96), .Z(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G29), .B2(G160), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT97), .Z(new_n735));
  OAI221_X1 g310(.A(new_n725), .B1(G1961), .B2(new_n728), .C1(new_n735), .C2(G2084), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT104), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(G2084), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n538), .A2(new_n674), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n674), .B2(G19), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G1341), .ZN(new_n742));
  INV_X1    g317(.A(G2090), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n697), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n697), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT29), .Z(new_n746));
  OAI211_X1 g321(.A(new_n738), .B(new_n742), .C1(new_n743), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n674), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n591), .B2(new_n674), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(G1348), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n749), .A2(G1348), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n747), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n746), .A2(new_n743), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g330(.A1(G164), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G27), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT105), .B(G2078), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n697), .A2(G26), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n478), .A2(G140), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n481), .A2(G128), .ZN(new_n765));
  OR2_X1    g340(.A1(G104), .A2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n766), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n763), .B1(new_n769), .B2(new_n697), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n758), .B2(new_n759), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n754), .A2(new_n755), .A3(new_n760), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n728), .A2(G1961), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT93), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT25), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n478), .A2(G139), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n604), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n777), .B(new_n778), .C1(new_n460), .C2(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G2072), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(KEYINPUT94), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n721), .A2(new_n724), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n674), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n774), .A2(new_n783), .A3(new_n784), .A4(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT31), .B(G11), .Z(new_n790));
  INV_X1    g365(.A(G28), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(KEYINPUT30), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT102), .Z(new_n793));
  AOI21_X1  g368(.A(G29), .B1(new_n791), .B2(KEYINPUT30), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n674), .A2(G21), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G168), .B2(new_n674), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n795), .B1(new_n697), .B2(new_n615), .C1(new_n797), .C2(G1966), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n781), .B2(G2072), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n741), .B2(G1341), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(G1966), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT101), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n782), .B2(KEYINPUT94), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n773), .A2(new_n789), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n712), .A2(new_n737), .A3(new_n752), .A4(new_n804), .ZN(G150));
  INV_X1    g380(.A(G150), .ZN(G311));
  INV_X1    g381(.A(G93), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n502), .A2(new_n807), .B1(new_n504), .B2(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n508), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n591), .A2(G559), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n812), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n538), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n537), .A2(new_n812), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n817), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n823), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n814), .B1(new_n824), .B2(new_n826), .ZN(G145));
  INV_X1    g402(.A(G37), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n498), .B(new_n769), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n780), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n720), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n704), .B(new_n606), .ZN(new_n832));
  AOI22_X1  g407(.A1(G130), .A2(new_n481), .B1(new_n478), .B2(G142), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT108), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n834), .A2(new_n460), .A3(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n460), .B2(G118), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n836), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n833), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n832), .B(new_n838), .Z(new_n839));
  OR2_X1    g414(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(G162), .B(G160), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n615), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n831), .A2(new_n839), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n828), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n845), .B(KEYINPUT109), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n840), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n846), .B1(new_n848), .B2(new_n842), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g425(.A(new_n600), .B(new_n821), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n588), .A2(new_n578), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G299), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT110), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n853), .B(KEYINPUT41), .Z(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  XNOR2_X1  g435(.A(G305), .B(G290), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n685), .B(G303), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n863), .B1(new_n859), .B2(new_n860), .ZN(new_n865));
  OAI21_X1  g440(.A(G868), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(G868), .B2(new_n818), .ZN(G295));
  OAI21_X1  g442(.A(new_n866), .B1(G868), .B2(new_n818), .ZN(G331));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n869));
  XNOR2_X1  g444(.A(G301), .B(G168), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n819), .A2(new_n820), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n819), .B2(new_n820), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n856), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT111), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n871), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n873), .B2(new_n876), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n853), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n863), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT112), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n828), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n875), .A2(new_n880), .A3(new_n863), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n881), .B2(new_n828), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n869), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n854), .A2(new_n874), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n878), .A2(new_n879), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(new_n856), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n863), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n828), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n869), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT44), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n885), .B2(new_n886), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(KEYINPUT43), .B2(new_n892), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n898), .ZN(G397));
  INV_X1    g474(.A(G1384), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n498), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(KEYINPUT113), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT45), .B1(new_n901), .B2(KEYINPUT113), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G40), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n465), .A2(new_n470), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(G1996), .A3(new_n720), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT114), .ZN(new_n910));
  INV_X1    g485(.A(G2067), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n768), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n720), .B2(G1996), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n704), .B(new_n708), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n908), .ZN(new_n918));
  XOR2_X1   g493(.A(G290), .B(G1986), .Z(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G8), .ZN(new_n921));
  OAI211_X1 g496(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n922));
  OR2_X1    g497(.A1(G102), .A2(G2105), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n487), .A3(G2104), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n493), .B1(new_n604), .B2(new_n495), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n484), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n483), .A2(KEYINPUT68), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(KEYINPUT4), .A3(new_n496), .ZN(new_n929));
  AOI21_X1  g504(.A(G1384), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n921), .B1(new_n930), .B2(new_n906), .ZN(new_n931));
  NOR2_X1   g506(.A1(G305), .A2(G1981), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G1981), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n564), .A2(new_n561), .A3(G651), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT71), .B1(new_n566), .B2(new_n508), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n935), .A2(new_n936), .B1(G48), .B2(new_n532), .ZN(new_n937));
  XOR2_X1   g512(.A(KEYINPUT119), .B(G86), .Z(new_n938));
  NAND2_X1  g513(.A1(new_n530), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n934), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n933), .A2(new_n941), .A3(KEYINPUT49), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT49), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n932), .B2(new_n940), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n944), .A3(new_n931), .ZN(new_n945));
  INV_X1    g520(.A(G1976), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n945), .A2(new_n946), .A3(new_n685), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n932), .B(KEYINPUT120), .Z(new_n948));
  OAI21_X1  g523(.A(new_n931), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n906), .B1(new_n930), .B2(KEYINPUT45), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  AOI211_X1 g526(.A(new_n951), .B(G1384), .C1(new_n927), .C2(new_n929), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT115), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n907), .B1(new_n901), .B2(new_n951), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT115), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n900), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1971), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT116), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n953), .A2(new_n957), .A3(new_n961), .A4(new_n958), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n963));
  NAND3_X1  g538(.A1(new_n498), .A2(new_n900), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n964), .B(new_n906), .C1(new_n930), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n743), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n960), .A2(new_n962), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(G303), .A2(G8), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT55), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(G8), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n931), .A2(new_n946), .A3(G288), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n685), .A2(G1976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n931), .A2(KEYINPUT118), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n931), .A2(new_n977), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(KEYINPUT118), .A3(new_n974), .A4(new_n975), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n945), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n949), .B1(new_n973), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n494), .A2(new_n497), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n490), .A2(new_n485), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n965), .B(new_n900), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(new_n906), .C1(new_n930), .C2(new_n963), .ZN(new_n987));
  INV_X1    g562(.A(G1956), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n990));
  XNOR2_X1  g565(.A(G299), .B(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT56), .B(G2072), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n954), .A2(new_n956), .A3(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT124), .B1(new_n989), .B2(new_n993), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n991), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n989), .A2(new_n993), .A3(KEYINPUT124), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n907), .B1(new_n930), .B2(new_n963), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n965), .B1(new_n498), .B2(new_n900), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1348), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n498), .A2(new_n900), .A3(new_n906), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT123), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n930), .A2(KEYINPUT123), .A3(new_n906), .ZN(new_n1007));
  AOI21_X1  g582(.A(G2067), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n591), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n994), .B1(new_n999), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT58), .B(G1341), .Z(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n1007), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n901), .A2(new_n951), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n956), .A4(new_n906), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT59), .B1(new_n1016), .B2(new_n538), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n1018), .B(new_n537), .C1(new_n1012), .C2(new_n1015), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT61), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n991), .B1(new_n989), .B2(new_n993), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n994), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT61), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n996), .B2(new_n998), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT60), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT123), .B1(new_n930), .B2(new_n906), .ZN(new_n1030));
  AND4_X1   g605(.A1(KEYINPUT123), .A2(new_n498), .A3(new_n900), .A4(new_n906), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n911), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1348), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n964), .A2(new_n906), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(new_n1001), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1029), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1009), .B1(new_n1036), .B2(new_n591), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1009), .B(new_n1038), .C1(new_n1036), .C2(new_n591), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1010), .B1(new_n1028), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G2078), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n956), .A2(KEYINPUT53), .A3(new_n1044), .A4(new_n906), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1961), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n904), .A2(new_n1046), .B1(new_n1047), .B2(new_n966), .ZN(new_n1048));
  AOI21_X1  g623(.A(G2078), .B1(new_n953), .B2(new_n957), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(G301), .C1(new_n1049), .C2(KEYINPUT53), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n966), .A2(new_n1047), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1013), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(new_n1045), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n950), .A2(KEYINPUT115), .A3(new_n952), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n955), .B1(new_n954), .B2(new_n956), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1044), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1050), .B1(new_n1058), .B2(G301), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1966), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n950), .B2(new_n952), .ZN(new_n1063));
  INV_X1    g638(.A(G2084), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1000), .A2(new_n1002), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(G168), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1066), .A2(new_n1067), .A3(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G286), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(G8), .A3(new_n1066), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1068), .B1(new_n1071), .B2(KEYINPUT51), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1053), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(G301), .C1(new_n1049), .C2(KEYINPUT53), .ZN(new_n1075));
  INV_X1    g650(.A(new_n904), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1051), .B1(new_n1076), .B2(new_n1045), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT54), .B(new_n1075), .C1(new_n1078), .C2(G301), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1061), .A2(new_n1073), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1049), .A2(KEYINPUT53), .ZN(new_n1081));
  OAI21_X1  g656(.A(G171), .B1(new_n1081), .B2(new_n1053), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1066), .A2(G8), .ZN(new_n1084));
  AOI21_X1  g659(.A(G168), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT51), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1066), .A2(new_n1067), .A3(G8), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1087), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1083), .B(new_n1089), .C1(new_n1090), .C2(KEYINPUT126), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT126), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1072), .A2(new_n1092), .A3(new_n1087), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1043), .A2(new_n1080), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n959), .B1(G2090), .B2(new_n987), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G8), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n982), .B1(new_n1096), .B2(new_n971), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n973), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n983), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n921), .B(G286), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n973), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT121), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1097), .A2(new_n973), .A3(new_n1105), .A4(new_n1101), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n972), .B1(new_n969), .B2(G8), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT122), .B1(new_n1108), .B2(new_n982), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  INV_X1    g685(.A(new_n982), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n959), .A2(KEYINPUT116), .B1(new_n743), .B2(new_n967), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n921), .B1(new_n1112), .B2(new_n962), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1110), .B(new_n1111), .C1(new_n1113), .C2(new_n972), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n973), .A2(KEYINPUT63), .A3(new_n1101), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1107), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n920), .B1(new_n1100), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n914), .A2(new_n705), .A3(new_n707), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n768), .A2(G2067), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n918), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n908), .A2(new_n1014), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT46), .ZN(new_n1126));
  INV_X1    g701(.A(new_n912), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n908), .B1(new_n720), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT47), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n918), .A2(G1986), .A3(G290), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT48), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n917), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1124), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT127), .B1(new_n1119), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1130), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n1123), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1106), .A2(new_n1104), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1139), .A2(new_n1103), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n997), .A2(new_n995), .A3(new_n991), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1009), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1025), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1020), .B(new_n1023), .C1(new_n1141), .C2(new_n1026), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1059), .A2(new_n1060), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n1079), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1092), .B1(new_n1072), .B2(new_n1087), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1082), .B1(new_n1072), .B2(new_n1087), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1090), .A2(KEYINPUT126), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1098), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1140), .A2(new_n1153), .A3(new_n983), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1136), .B(new_n1138), .C1(new_n1154), .C2(new_n920), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1135), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g731(.A(G319), .ZN(new_n1158));
  OR3_X1    g732(.A1(G401), .A2(new_n1158), .A3(G227), .ZN(new_n1159));
  NOR3_X1   g733(.A1(new_n849), .A2(G229), .A3(new_n1159), .ZN(new_n1160));
  AND2_X1   g734(.A1(new_n1160), .A2(new_n896), .ZN(G308));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n896), .ZN(G225));
endmodule


