//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n203), .A2(KEYINPUT65), .A3(G131), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT65), .B1(new_n203), .B2(G131), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n199), .A2(new_n201), .A3(new_n207), .A4(new_n202), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT80), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT78), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT67), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  AND4_X1   g034(.A1(KEYINPUT67), .A2(new_n215), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n212), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n218), .A3(new_n220), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n213), .A2(KEYINPUT67), .A3(new_n215), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT78), .ZN(new_n227));
  INV_X1    g041(.A(new_n213), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n214), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n222), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G101), .ZN(new_n232));
  INV_X1    g046(.A(G104), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G107), .ZN(new_n234));
  INV_X1    g048(.A(G107), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n235), .A2(KEYINPUT3), .A3(G104), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT3), .B1(new_n235), .B2(G104), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n232), .B(new_n234), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT77), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n235), .A2(G104), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n233), .B2(G107), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n235), .A2(KEYINPUT3), .A3(G104), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT77), .A3(new_n232), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n235), .A2(G104), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n234), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n240), .A2(new_n246), .B1(G101), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n231), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n219), .C2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G128), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT68), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n228), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT69), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(new_n228), .C1(new_n252), .C2(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n248), .A2(G101), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n243), .A2(new_n244), .ZN(new_n260));
  AND4_X1   g074(.A1(KEYINPUT77), .A2(new_n260), .A3(new_n232), .A4(new_n234), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT77), .B1(new_n245), .B2(new_n232), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n225), .A2(new_n226), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n258), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI211_X1 g079(.A(KEYINPUT12), .B(new_n211), .C1(new_n250), .C2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT12), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n250), .ZN(new_n268));
  INV_X1    g082(.A(new_n211), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT10), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n232), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n240), .A2(new_n246), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n260), .A2(new_n234), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G101), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n273), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  OR2_X1    g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n213), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n213), .A2(new_n280), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n250), .A2(new_n272), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n255), .A2(new_n257), .B1(new_n225), .B2(new_n226), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT10), .A3(new_n249), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT79), .B1(new_n206), .B2(new_n210), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n203), .A2(G131), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n203), .A2(KEYINPUT65), .A3(G131), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n208), .B(KEYINPUT64), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT79), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n285), .A2(new_n288), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n196), .B1(new_n271), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n285), .A2(new_n288), .A3(new_n298), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n294), .A2(new_n295), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(new_n285), .B2(new_n288), .ZN(new_n304));
  INV_X1    g118(.A(new_n196), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT81), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n268), .A2(new_n269), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT12), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n268), .A2(new_n267), .A3(new_n269), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n299), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n305), .ZN(new_n312));
  INV_X1    g126(.A(new_n304), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n299), .A3(new_n196), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n192), .B1(new_n307), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n305), .B1(new_n301), .B2(new_n304), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n309), .A2(new_n299), .A3(new_n196), .A4(new_n310), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n192), .A3(new_n189), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n192), .A2(new_n189), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n191), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n277), .B1(new_n261), .B2(new_n262), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT71), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n329));
  INV_X1    g143(.A(G113), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(KEYINPUT71), .A2(KEYINPUT2), .A3(G113), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT70), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(KEYINPUT2), .B2(G113), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n331), .A2(new_n332), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G116), .B(G119), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n273), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(KEYINPUT5), .ZN(new_n343));
  INV_X1    g157(.A(G116), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n344), .A2(KEYINPUT5), .A3(G119), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n330), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n336), .A2(new_n337), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n249), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g163(.A(G110), .B(G122), .Z(new_n350));
  AOI21_X1  g164(.A(new_n326), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n278), .A2(new_n340), .B1(new_n249), .B2(new_n347), .ZN(new_n353));
  INV_X1    g167(.A(new_n350), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n352), .A2(new_n342), .A3(new_n348), .A4(new_n354), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n284), .A2(G125), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n286), .B2(G125), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT84), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n363), .B(new_n360), .C1(new_n286), .C2(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT85), .B(G224), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G953), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n362), .A2(new_n368), .A3(new_n364), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(KEYINPUT83), .B(new_n351), .C1(new_n355), .C2(new_n356), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n349), .A2(new_n326), .A3(new_n350), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n359), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n355), .A2(new_n356), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n350), .B(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n249), .A2(new_n347), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(new_n348), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n369), .A2(KEYINPUT7), .ZN(new_n381));
  OR2_X1    g195(.A1(new_n361), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n361), .A2(new_n381), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(G902), .B1(new_n376), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G210), .B1(G237), .B2(G902), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n387), .B(KEYINPUT87), .Z(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G214), .B1(G237), .B2(G902), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n375), .A2(new_n385), .A3(new_n388), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n325), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G125), .ZN(new_n396));
  INV_X1    g210(.A(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT16), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT74), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G125), .B(G140), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n217), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n401), .A2(new_n403), .A3(G146), .A4(new_n404), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT23), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(G119), .B2(new_n214), .ZN(new_n410));
  INV_X1    g224(.A(G119), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n411), .A2(KEYINPUT23), .A3(G128), .ZN(new_n412));
  OAI22_X1  g226(.A1(new_n410), .A2(new_n412), .B1(G119), .B2(new_n214), .ZN(new_n413));
  XNOR2_X1  g227(.A(G119), .B(G128), .ZN(new_n414));
  XOR2_X1   g228(.A(KEYINPUT24), .B(G110), .Z(new_n415));
  AOI22_X1  g229(.A1(new_n413), .A2(G110), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n408), .A2(new_n416), .ZN(new_n417));
  OAI22_X1  g231(.A1(new_n413), .A2(G110), .B1(new_n414), .B2(new_n415), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT75), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n402), .A2(new_n217), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n418), .A2(new_n407), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n407), .A3(new_n420), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G137), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n417), .A2(new_n421), .A3(new_n423), .A4(new_n427), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G217), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(G234), .B2(new_n189), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(new_n189), .A3(new_n430), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT25), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n429), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n430), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(KEYINPUT76), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT76), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n442), .A3(new_n437), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n433), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n435), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT30), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT66), .ZN(new_n447));
  XNOR2_X1  g261(.A(G134), .B(G137), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n448), .B2(new_n207), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n200), .A2(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n202), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT66), .A3(G131), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n258), .B2(new_n264), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n283), .B1(new_n294), .B2(new_n295), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n446), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n284), .B1(new_n206), .B2(new_n210), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(KEYINPUT30), .C1(new_n286), .C2(new_n456), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n340), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n457), .A2(new_n458), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT72), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n340), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT72), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(G237), .A2(G953), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G210), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n232), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n462), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT31), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n463), .A2(new_n467), .A3(KEYINPUT28), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n460), .B1(new_n286), .B2(new_n456), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n465), .A2(new_n466), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n340), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n477), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n473), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT31), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n462), .A2(new_n485), .A3(new_n468), .A4(new_n474), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n476), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(G472), .A2(G902), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n487), .A2(KEYINPUT32), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT32), .B1(new_n487), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n462), .A2(new_n468), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n473), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n477), .A2(new_n481), .A3(new_n482), .A4(new_n474), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n493), .A2(KEYINPUT73), .A3(new_n494), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n479), .A2(new_n480), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n473), .A2(new_n494), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n477), .A2(new_n481), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n189), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G472), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n445), .B1(new_n491), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n469), .A2(G143), .A3(G214), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(G143), .B1(new_n469), .B2(G214), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n194), .A3(G214), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n219), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n207), .A3(new_n510), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n396), .A2(new_n398), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT19), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT19), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n402), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n522), .A3(new_n217), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n407), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n516), .B(new_n510), .C1(new_n525), .C2(new_n207), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n519), .A2(G146), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n420), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n526), .B(new_n528), .C1(new_n513), .C2(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(G113), .B(G122), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(new_n233), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT88), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n535), .B(new_n532), .C1(new_n524), .C2(new_n529), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n513), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT17), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n513), .A2(new_n541), .A3(new_n517), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT89), .B1(new_n513), .B2(new_n541), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n532), .B(new_n529), .C1(new_n544), .C2(new_n408), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n509), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT90), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n530), .A2(new_n533), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n535), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n530), .A2(KEYINPUT88), .A3(new_n533), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n545), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n508), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT90), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n546), .A2(new_n547), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT91), .B1(new_n214), .B2(G143), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n219), .A3(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT13), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n558), .A2(new_n560), .A3(KEYINPUT13), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n214), .A2(G143), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(KEYINPUT92), .A3(G134), .ZN(new_n567));
  XOR2_X1   g381(.A(G116), .B(G122), .Z(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G107), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n198), .A3(new_n565), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n561), .A2(new_n562), .B1(new_n214), .B2(G143), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n198), .B1(new_n572), .B2(new_n564), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n567), .B(new_n569), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n188), .A2(G217), .A3(new_n194), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n344), .A2(G122), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n235), .B1(new_n577), .B2(KEYINPUT14), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n578), .A2(new_n568), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n568), .ZN(new_n580));
  INV_X1    g394(.A(new_n570), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n198), .B1(new_n561), .B2(new_n565), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n574), .A2(new_n576), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n576), .B1(new_n574), .B2(new_n583), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n189), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n567), .A2(new_n569), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n573), .A2(new_n571), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n583), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n575), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n574), .A2(new_n576), .A3(new_n583), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT93), .A3(new_n189), .ZN(new_n595));
  INV_X1    g409(.A(G478), .ZN(new_n596));
  AOI211_X1 g410(.A(KEYINPUT15), .B(new_n596), .C1(new_n587), .C2(KEYINPUT94), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n588), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  OAI22_X1  g412(.A1(new_n586), .A2(KEYINPUT94), .B1(KEYINPUT15), .B2(new_n596), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(G234), .A2(G237), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(G952), .A3(new_n194), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT21), .B(G898), .Z(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(G902), .A3(G953), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n603), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n529), .B1(new_n544), .B2(new_n408), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n533), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n545), .ZN(new_n612));
  OAI21_X1  g426(.A(G475), .B1(new_n612), .B2(G902), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n557), .A2(new_n600), .A3(new_n609), .A4(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n394), .A2(new_n507), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G101), .ZN(G3));
  NOR3_X1   g431(.A1(new_n300), .A2(new_n306), .A3(KEYINPUT81), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n315), .B1(new_n312), .B2(new_n314), .ZN(new_n619));
  OAI21_X1  g433(.A(G469), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI211_X1 g434(.A(G469), .B(G902), .C1(new_n318), .C2(new_n319), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n322), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n190), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n443), .A2(new_n433), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n624), .A2(new_n440), .B1(new_n431), .B2(new_n434), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n487), .A2(new_n488), .ZN(new_n626));
  INV_X1    g440(.A(G472), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n487), .B2(new_n189), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n623), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n594), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n632), .A2(KEYINPUT33), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(KEYINPUT33), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n633), .A2(G478), .A3(new_n189), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n588), .A2(new_n595), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT95), .B1(new_n636), .B2(new_n596), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n638), .B(G478), .C1(new_n588), .C2(new_n595), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n557), .A2(new_n613), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n609), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n393), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n631), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  XOR2_X1   g460(.A(new_n608), .B(KEYINPUT96), .Z(new_n647));
  AND4_X1   g461(.A1(new_n391), .A2(new_n390), .A3(new_n392), .A4(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT97), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n641), .A2(new_n600), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n390), .A2(new_n391), .A3(new_n392), .A4(new_n647), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n557), .A2(new_n613), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n598), .A2(new_n599), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT97), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n631), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NOR2_X1   g474(.A1(new_n428), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n424), .B(new_n661), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n624), .A2(new_n440), .B1(new_n434), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n614), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n664), .A2(new_n629), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n394), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n603), .B1(new_n607), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n654), .A2(new_n613), .A3(new_n557), .A4(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n663), .B1(new_n491), .B2(new_n506), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n394), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  INV_X1    g491(.A(new_n392), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n388), .B1(new_n375), .B2(new_n385), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n600), .B1(new_n557), .B2(new_n613), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n391), .A3(new_n663), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n670), .B(KEYINPUT39), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n623), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n685), .B1(new_n688), .B2(KEYINPUT40), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n683), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n492), .A2(new_n474), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n474), .B1(new_n463), .B2(new_n467), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n694), .B2(new_n500), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n627), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n692), .B1(new_n491), .B2(new_n697), .ZN(new_n698));
  NOR4_X1   g512(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT100), .A4(new_n696), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n691), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n219), .ZN(G45));
  NAND2_X1  g516(.A1(new_n640), .A2(new_n641), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n670), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n394), .A2(new_n675), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  AOI21_X1  g520(.A(new_n192), .B1(new_n320), .B2(new_n189), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n707), .A2(new_n621), .A3(new_n190), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n643), .A2(new_n507), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND2_X1  g525(.A1(new_n491), .A2(new_n506), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n625), .A3(new_n708), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n651), .B2(new_n656), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n344), .ZN(G18));
  INV_X1    g529(.A(new_n393), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n712), .A2(new_n716), .A3(new_n664), .A4(new_n708), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT101), .B(G119), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G21));
  AND3_X1   g533(.A1(new_n477), .A2(new_n481), .A3(new_n500), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n476), .B(new_n486), .C1(new_n474), .C2(new_n720), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n721), .A2(new_n488), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n445), .A3(new_n628), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n648), .A2(new_n684), .A3(new_n708), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NOR3_X1   g539(.A1(new_n722), .A2(new_n663), .A3(new_n628), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n704), .A2(new_n716), .A3(new_n708), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  OAI21_X1  g542(.A(new_n391), .B1(new_n678), .B2(new_n679), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n312), .A2(new_n314), .A3(G469), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n321), .A2(new_n323), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n191), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n507), .A3(new_n704), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n507), .A3(KEYINPUT42), .A4(new_n704), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  AND3_X1   g553(.A1(new_n674), .A2(new_n733), .A3(new_n507), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT102), .B(G134), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G36));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n640), .A2(new_n653), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n653), .A2(KEYINPUT103), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n641), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n640), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n744), .B1(new_n748), .B2(KEYINPUT43), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  AOI211_X1 g564(.A(new_n629), .B(new_n663), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT105), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n751), .A2(new_n756), .A3(KEYINPUT44), .A4(new_n752), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT45), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n300), .A2(new_n306), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n192), .B1(new_n760), .B2(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n322), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT46), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n621), .B1(new_n762), .B2(KEYINPUT46), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n190), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n687), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n729), .B(new_n766), .C1(new_n753), .C2(new_n754), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  NAND2_X1  g583(.A1(new_n763), .A2(new_n764), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n191), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(KEYINPUT47), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n765), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n704), .A2(new_n445), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n712), .A3(new_n729), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT106), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT107), .B(G140), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G42));
  NAND3_X1  g595(.A1(new_n625), .A2(new_n391), .A3(new_n191), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT108), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n707), .A2(new_n621), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n748), .B(new_n783), .C1(KEYINPUT49), .C2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT109), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n785), .A2(KEYINPUT49), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n700), .A3(new_n682), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n616), .A2(new_n666), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n625), .B(new_n191), .C1(new_n317), .C2(new_n324), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n703), .A2(new_n655), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n648), .A3(new_n629), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n790), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n325), .A2(new_n393), .A3(new_n614), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n798), .A2(new_n507), .B1(new_n394), .B2(new_n665), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(KEYINPUT110), .A3(new_n795), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n663), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n489), .A2(new_n490), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n503), .B1(new_n496), .B2(new_n497), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n627), .B1(new_n804), .B2(new_n499), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n391), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n390), .B2(new_n392), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n641), .A2(new_n654), .A3(new_n670), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n623), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n636), .A2(new_n596), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n638), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n636), .A2(KEYINPUT95), .A3(new_n596), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n814), .A2(new_n635), .B1(new_n613), .B2(new_n557), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n726), .A2(new_n815), .A3(new_n671), .ZN(new_n816));
  INV_X1    g630(.A(new_n732), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n808), .ZN(new_n818));
  OAI22_X1  g632(.A1(new_n806), .A2(new_n810), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n740), .B1(new_n736), .B2(new_n737), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n801), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n714), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n709), .A2(new_n717), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n724), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n709), .A2(new_n717), .A3(new_n724), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT115), .B1(new_n829), .B2(new_n714), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n676), .A2(new_n727), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n390), .A2(new_n684), .A3(new_n391), .A4(new_n392), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n732), .A2(new_n802), .A3(new_n670), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n835), .B(new_n836), .C1(new_n698), .C2(new_n699), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n832), .A2(new_n833), .A3(new_n705), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n676), .A3(new_n705), .A4(new_n727), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n824), .A2(new_n831), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n839), .A2(KEYINPUT52), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n839), .A2(KEYINPUT52), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT112), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n838), .A2(new_n846), .A3(new_n840), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n740), .B(new_n819), .C1(new_n736), .C2(new_n737), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n829), .A2(new_n714), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n801), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT110), .B1(new_n799), .B2(new_n795), .ZN(new_n853));
  AND4_X1   g667(.A1(KEYINPUT110), .A2(new_n616), .A3(new_n795), .A4(new_n666), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n823), .A2(new_n820), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT111), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n848), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AOI211_X1 g674(.A(KEYINPUT54), .B(new_n842), .C1(new_n858), .C2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n857), .A2(new_n852), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n859), .A4(new_n848), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n848), .A2(new_n859), .A3(new_n852), .A4(new_n857), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT114), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n857), .A2(new_n852), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n868), .B2(new_n841), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n861), .B1(new_n870), .B2(KEYINPUT54), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n784), .A2(KEYINPUT116), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n784), .A2(KEYINPUT116), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n190), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT118), .B1(new_n775), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n874), .C1(new_n772), .C2(new_n774), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n749), .A2(new_n603), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n723), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n876), .A2(new_n808), .A3(new_n878), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n723), .A2(new_n708), .ZN(new_n883));
  NOR2_X1   g697(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n391), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n880), .A2(new_n682), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n808), .A2(new_n708), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n889), .A2(new_n445), .A3(new_n602), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n700), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n891), .A2(new_n641), .A3(new_n640), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n879), .A2(new_n889), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n726), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n888), .A2(KEYINPUT51), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n882), .A2(new_n895), .A3(KEYINPUT119), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT119), .B1(new_n882), .B2(new_n895), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n893), .A2(new_n507), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n893), .A2(KEYINPUT120), .A3(new_n507), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT48), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT48), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n881), .A2(new_n716), .A3(new_n708), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n890), .A2(new_n815), .A3(new_n700), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n907), .A2(G952), .A3(new_n194), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n903), .A2(new_n905), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n775), .A2(new_n875), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n881), .A2(new_n808), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n888), .B(new_n894), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n871), .A2(new_n898), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(G952), .A2(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n789), .B1(new_n915), .B2(new_n916), .ZN(G75));
  AND3_X1   g731(.A1(new_n838), .A2(new_n846), .A3(new_n840), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n846), .B1(new_n838), .B2(new_n840), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n860), .B1(new_n868), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n842), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n189), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT56), .B1(new_n923), .B2(new_n388), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n359), .A2(new_n373), .A3(new_n374), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n372), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT55), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n924), .A2(new_n927), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n194), .A2(G952), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT121), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n928), .A2(new_n929), .A3(new_n932), .ZN(G51));
  INV_X1    g747(.A(KEYINPUT54), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n921), .B2(new_n922), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n861), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n323), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n320), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n923), .A2(new_n759), .A3(new_n761), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n932), .B1(new_n939), .B2(new_n940), .ZN(G54));
  AND2_X1   g755(.A1(KEYINPUT58), .A2(G475), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n923), .A2(new_n552), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n552), .B1(new_n923), .B2(new_n942), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n944), .A3(new_n932), .ZN(G60));
  NAND2_X1  g759(.A1(new_n633), .A2(new_n634), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n871), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n946), .A2(new_n948), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n861), .B2(new_n935), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n932), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT123), .B(new_n950), .C1(new_n861), .C2(new_n935), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(new_n921), .A2(new_n922), .ZN(new_n956));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT124), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n431), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n662), .B(KEYINPUT125), .Z(new_n963));
  NAND3_X1  g777(.A1(new_n956), .A2(new_n959), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n931), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n931), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(G66));
  OAI21_X1  g783(.A(G953), .B1(new_n605), .B2(new_n367), .ZN(new_n970));
  INV_X1    g784(.A(new_n855), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n925), .B1(G898), .B2(new_n194), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G69));
  NAND2_X1  g788(.A1(new_n459), .A2(new_n461), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT126), .Z(new_n976));
  AND2_X1   g790(.A1(new_n520), .A2(new_n522), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n976), .B(new_n977), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n832), .A2(new_n705), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n701), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT62), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n778), .A2(KEYINPUT106), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT106), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n775), .B2(new_n777), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n794), .A2(new_n623), .A3(new_n687), .A4(new_n808), .ZN(new_n988));
  INV_X1    g802(.A(new_n507), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n987), .B1(new_n768), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n768), .A2(new_n987), .A3(new_n991), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n986), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n979), .B1(new_n995), .B2(G953), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n766), .A2(new_n989), .A3(new_n834), .ZN(new_n999));
  INV_X1    g813(.A(new_n738), .ZN(new_n1000));
  NOR4_X1   g814(.A1(new_n999), .A2(new_n1000), .A3(new_n740), .A4(new_n980), .ZN(new_n1001));
  AND4_X1   g815(.A1(new_n194), .A2(new_n779), .A3(new_n768), .A4(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n978), .B1(new_n669), .B2(new_n194), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n996), .B(new_n998), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g818(.A(KEYINPUT127), .B(new_n990), .C1(new_n758), .C2(new_n767), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n779), .B(new_n982), .C1(new_n992), .C2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n978), .B1(new_n1006), .B2(new_n194), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n997), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1004), .A2(new_n1009), .ZN(G72));
  NAND4_X1  g824(.A1(new_n779), .A2(new_n768), .A3(new_n971), .A4(new_n1001), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n492), .A2(new_n474), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n932), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1013), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n995), .B2(new_n971), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n1018), .B2(new_n693), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(new_n493), .B2(new_n475), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n870), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1019), .A2(new_n1021), .ZN(G57));
endmodule


