//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT93), .ZN(new_n205));
  INV_X1    g004(.A(G15gat), .ZN(new_n206));
  INV_X1    g005(.A(G22gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G15gat), .A2(G22gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(new_n212), .A3(G8gat), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n204), .B(new_n211), .C1(KEYINPUT93), .C2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218));
  INV_X1    g017(.A(G71gat), .ZN(new_n219));
  INV_X1    g018(.A(G78gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT96), .ZN(new_n222));
  XOR2_X1   g021(.A(G57gat), .B(G64gat), .Z(new_n223));
  XNOR2_X1  g022(.A(G71gat), .B(G78gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT96), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n225), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n224), .ZN(new_n228));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n218), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n216), .B1(new_n217), .B2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(G183gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(G183gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(G231gat), .A2(G233gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n233), .B2(new_n234), .ZN(new_n238));
  XOR2_X1   g037(.A(G127gat), .B(G155gat), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT97), .ZN(new_n240));
  OR3_X1    g039(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n237), .B2(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n231), .A2(new_n217), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n244));
  INV_X1    g043(.A(G211gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n243), .B(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n241), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n241), .B2(new_n242), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT92), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT15), .ZN(new_n253));
  INV_X1    g052(.A(G43gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(G50gat), .ZN(new_n255));
  INV_X1    g054(.A(G50gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G43gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n253), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(G43gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(G50gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT15), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G29gat), .ZN(new_n263));
  INV_X1    g062(.A(G36gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT14), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT14), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(G29gat), .B2(G36gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G29gat), .A2(G36gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT91), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT91), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n258), .A4(new_n261), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT90), .B1(new_n271), .B2(new_n261), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT15), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT90), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n270), .A2(new_n273), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n252), .B1(new_n278), .B2(KEYINPUT17), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n277), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT15), .B1(new_n259), .B2(new_n260), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n272), .B1(new_n282), .B2(new_n271), .ZN(new_n283));
  AND4_X1   g082(.A1(new_n272), .A2(new_n271), .A3(new_n261), .A4(new_n258), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT17), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT92), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT17), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(G99gat), .A2(G106gat), .ZN(new_n290));
  INV_X1    g089(.A(G85gat), .ZN(new_n291));
  INV_X1    g090(.A(G92gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(KEYINPUT8), .A2(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n291), .B2(new_n292), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G99gat), .B(G106gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT98), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(G99gat), .A2(G106gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT98), .A3(new_n290), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n297), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n300), .A3(new_n302), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n288), .B(new_n289), .C1(new_n303), .C2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G134gat), .B(G162gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n305), .A2(new_n303), .ZN(new_n309));
  AND2_X1   g108(.A1(G232gat), .A2(G233gat), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n285), .A2(new_n309), .B1(KEYINPUT41), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n310), .A2(KEYINPUT41), .ZN(new_n314));
  XNOR2_X1  g113(.A(G190gat), .B(G218gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n308), .B1(new_n306), .B2(new_n311), .ZN(new_n318));
  OR3_X1    g117(.A1(new_n313), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n313), .B2(new_n318), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n251), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n227), .A2(new_n230), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n300), .A2(new_n302), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n324), .A2(new_n293), .A3(new_n295), .A4(new_n296), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT99), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n300), .A2(new_n326), .A3(new_n302), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n323), .A2(new_n325), .A3(new_n304), .A4(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT10), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n227), .A3(new_n230), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n305), .B2(new_n303), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n309), .A2(KEYINPUT10), .A3(new_n323), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n328), .A2(new_n331), .ZN(new_n337));
  INV_X1    g136(.A(new_n335), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G120gat), .B(G148gat), .ZN(new_n340));
  INV_X1    g139(.A(G176gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(G204gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n343), .ZN(new_n345));
  INV_X1    g144(.A(new_n339), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n335), .B(KEYINPUT100), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n332), .B2(new_n333), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n322), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT38), .ZN(new_n353));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G169gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n341), .A3(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT26), .ZN(new_n358));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT26), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(KEYINPUT67), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n366));
  INV_X1    g165(.A(G190gat), .ZN(new_n367));
  AND2_X1   g166(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n365), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n370), .B(KEYINPUT28), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n363), .A2(new_n364), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT68), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379));
  INV_X1    g178(.A(new_n364), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT24), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT65), .B1(new_n360), .B2(KEYINPUT23), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n360), .A2(KEYINPUT23), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n388), .B(new_n389), .C1(G169gat), .C2(G176gat), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n386), .A2(new_n359), .A3(new_n387), .A4(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n379), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT24), .B1(new_n380), .B2(KEYINPUT66), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(new_n384), .C1(KEYINPUT66), .C2(new_n383), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT25), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n392), .B1(new_n395), .B2(new_n391), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n377), .A2(new_n378), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n378), .B1(new_n377), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n355), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n365), .A2(new_n372), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n354), .B1(new_n401), .B2(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT76), .ZN(new_n403));
  XOR2_X1   g202(.A(KEYINPUT73), .B(G204gat), .Z(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G197gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT73), .B(G204gat), .ZN(new_n406));
  INV_X1    g205(.A(G197gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(G211gat), .A2(G218gat), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n405), .B(new_n408), .C1(KEYINPUT22), .C2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(G211gat), .A2(G218gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n410), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n414), .B(new_n354), .C1(new_n401), .C2(KEYINPUT29), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n399), .A2(new_n403), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT37), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(new_n355), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n397), .B2(new_n398), .ZN(new_n420));
  INV_X1    g219(.A(new_n412), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n410), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n401), .A2(new_n355), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n417), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT77), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G8gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(new_n264), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n423), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n377), .A2(new_n396), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT74), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n377), .A2(new_n378), .A3(new_n396), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n431), .B1(new_n435), .B2(new_n419), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT86), .B1(new_n436), .B2(new_n422), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n399), .A2(new_n403), .A3(new_n415), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n422), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n423), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n413), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n437), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n353), .B(new_n430), .C1(new_n443), .C2(new_n417), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT0), .B(G57gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(G85gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G113gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G120gat), .ZN(new_n451));
  INV_X1    g250(.A(G120gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(G113gat), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT1), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455));
  XNOR2_X1  g254(.A(G127gat), .B(G134gat), .ZN(new_n456));
  OR3_X1    g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n454), .B2(new_n456), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT70), .B(G120gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(G113gat), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT1), .B1(new_n461), .B2(new_n451), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n456), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT2), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(G155gat), .B2(G162gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT81), .ZN(new_n467));
  INV_X1    g266(.A(G148gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G141gat), .ZN(new_n469));
  XOR2_X1   g268(.A(KEYINPUT79), .B(G141gat), .Z(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(new_n468), .ZN(new_n471));
  XNOR2_X1  g270(.A(G155gat), .B(G162gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT80), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n472), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT80), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n467), .A2(new_n471), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G141gat), .B(G148gat), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n478), .B2(new_n466), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT83), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n459), .A2(new_n477), .A3(new_n479), .A4(new_n463), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n464), .A2(new_n480), .A3(KEYINPUT83), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n480), .A2(KEYINPUT3), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n477), .A2(new_n490), .A3(new_n479), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n464), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n464), .ZN(new_n493));
  INV_X1    g292(.A(new_n480), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT4), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n486), .B1(new_n483), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n488), .A2(new_n498), .A3(KEYINPUT5), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n483), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n449), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n498), .A3(KEYINPUT5), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n502), .A2(new_n503), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n507), .B(new_n448), .C1(new_n508), .C2(new_n501), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n416), .A2(new_n424), .ZN(new_n511));
  INV_X1    g310(.A(new_n429), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT6), .B(new_n449), .C1(new_n499), .C2(new_n504), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n444), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n430), .B1(new_n417), .B2(new_n511), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT38), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n444), .A2(new_n515), .A3(KEYINPUT87), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n490), .B1(new_n422), .B2(new_n418), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n523), .A2(new_n480), .B1(G228gat), .B2(G233gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n418), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n491), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n413), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n413), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n494), .B1(new_n529), .B2(new_n490), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n526), .A2(new_n413), .ZN(new_n531));
  OAI211_X1 g330(.A(G228gat), .B(G233gat), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G78gat), .B(G106gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(new_n256), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n533), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(new_n207), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n537), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n513), .A2(KEYINPUT78), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT30), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n511), .A2(new_n512), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n513), .A2(KEYINPUT78), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n502), .A2(new_n486), .A3(new_n503), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n484), .A2(new_n487), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n485), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT85), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n548), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT39), .B1(new_n550), .B2(new_n551), .ZN(new_n554));
  OAI221_X1 g353(.A(new_n448), .B1(KEYINPUT39), .B2(new_n548), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT40), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n547), .A2(new_n505), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n522), .A2(new_n541), .A3(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n510), .A2(new_n514), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n540), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT71), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n432), .A2(new_n464), .ZN(new_n564));
  NAND2_X1  g363(.A1(G227gat), .A2(G233gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n377), .A2(new_n493), .A3(new_n396), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT34), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n565), .B(KEYINPUT64), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT34), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n564), .A2(new_n566), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n564), .A2(new_n566), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n570), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT32), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G15gat), .B(G43gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G71gat), .B(G99gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n569), .B1(new_n564), .B2(new_n566), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n584), .B2(KEYINPUT33), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT32), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI211_X1 g387(.A(new_n563), .B(new_n574), .C1(new_n583), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n588), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n573), .B1(new_n590), .B2(KEYINPUT71), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT72), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n573), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n583), .A2(new_n588), .A3(new_n574), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT36), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598));
  INV_X1    g397(.A(new_n595), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n574), .B1(new_n583), .B2(new_n588), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n593), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n558), .A2(new_n562), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n541), .A2(new_n592), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT35), .B1(new_n604), .B2(new_n561), .ZN(new_n605));
  INV_X1    g404(.A(new_n560), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n540), .A2(new_n606), .A3(KEYINPUT35), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT88), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n599), .B2(new_n600), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT88), .A3(new_n595), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(new_n547), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n603), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n216), .A2(new_n278), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n213), .A2(new_n215), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n278), .B2(KEYINPUT17), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n288), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT18), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n289), .A2(new_n216), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n279), .B2(new_n287), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  INV_X1    g423(.A(new_n620), .ZN(new_n625));
  NOR4_X1   g424(.A1(new_n623), .A2(new_n624), .A3(new_n616), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT11), .B(G169gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G197gat), .ZN(new_n629));
  XOR2_X1   g428(.A(G113gat), .B(G141gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n285), .B(new_n617), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n620), .B(KEYINPUT13), .Z(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n627), .A2(KEYINPUT94), .A3(new_n632), .A4(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n278), .A2(new_n252), .A3(KEYINPUT17), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT92), .B1(new_n285), .B2(new_n286), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n618), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n616), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n640), .A3(new_n620), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n624), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n639), .A2(KEYINPUT18), .A3(new_n640), .A4(new_n620), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n642), .A2(new_n632), .A3(new_n635), .A4(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n635), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT89), .Z(new_n648));
  AOI22_X1  g447(.A1(new_n636), .A2(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n615), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n615), .A2(KEYINPUT95), .A3(new_n650), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n352), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n606), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n547), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n214), .B1(new_n655), .B2(new_n547), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(G1325gat));
  INV_X1    g466(.A(new_n611), .ZN(new_n668));
  AOI21_X1  g467(.A(G15gat), .B1(new_n655), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n597), .A2(new_n670), .A3(new_n601), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n585), .A2(new_n587), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n585), .A2(new_n587), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT71), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n574), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n590), .A2(new_n573), .A3(KEYINPUT71), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT72), .B1(new_n599), .B2(new_n600), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n598), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n601), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT103), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n671), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n206), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT104), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n669), .B1(new_n655), .B2(new_n684), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n655), .A2(new_n540), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NAND3_X1  g487(.A1(new_n615), .A2(KEYINPUT44), .A3(new_n321), .ZN(new_n689));
  INV_X1    g488(.A(new_n351), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n250), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n649), .ZN(new_n693));
  INV_X1    g492(.A(new_n321), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n682), .A2(new_n558), .A3(new_n562), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n614), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n689), .B(new_n693), .C1(KEYINPUT44), .C2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n560), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n653), .A2(new_n654), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n692), .A2(new_n694), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n263), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n699), .B1(new_n703), .B2(new_n606), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n702), .A2(KEYINPUT45), .A3(new_n560), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n698), .B1(new_n704), .B2(new_n705), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n559), .A2(G36gat), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n700), .A2(new_n707), .A3(new_n701), .A4(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G36gat), .B1(new_n697), .B2(new_n559), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT95), .B1(new_n615), .B2(new_n650), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n652), .B(new_n649), .C1(new_n603), .C2(new_n614), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n701), .B(new_n708), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT46), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n709), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT105), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n709), .A2(new_n710), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1329gat));
  OAI21_X1  g518(.A(G43gat), .B1(new_n697), .B2(new_n682), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n611), .A2(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n700), .A2(new_n701), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT47), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  AOI211_X1 g525(.A(KEYINPUT106), .B(new_n726), .C1(new_n720), .C2(new_n722), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(G1330gat));
  OAI21_X1  g527(.A(G50gat), .B1(new_n697), .B2(new_n541), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n541), .A2(G50gat), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n701), .B(new_n730), .C1(new_n711), .C2(new_n712), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(KEYINPUT48), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n700), .A2(new_n733), .A3(new_n701), .A4(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(KEYINPUT108), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n734), .A2(new_n729), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n732), .B1(new_n736), .B2(new_n737), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n695), .A2(new_n614), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n650), .A2(new_n351), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n322), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n560), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT109), .B(G57gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n559), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  OAI21_X1  g548(.A(new_n219), .B1(new_n741), .B2(new_n611), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n741), .A2(new_n219), .A3(new_n682), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT110), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n752), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(new_n750), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n753), .A2(new_n756), .A3(KEYINPUT50), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n741), .A2(new_n541), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT111), .B(G78gat), .Z(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT112), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n762), .B(new_n764), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n650), .A2(new_n250), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n696), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n696), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(KEYINPUT113), .A3(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n775), .A2(new_n291), .A3(new_n606), .A4(new_n690), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n766), .A2(new_n690), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n689), .B(new_n778), .C1(KEYINPUT44), .C2(new_n696), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n560), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(G1336gat));
  AND3_X1   g580(.A1(new_n696), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT51), .B1(new_n696), .B2(new_n766), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n547), .B(new_n690), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n779), .A2(new_n559), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n292), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT52), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n790));
  AOI211_X1 g589(.A(new_n790), .B(new_n694), .C1(new_n603), .C2(new_n614), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n547), .A4(new_n778), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT114), .B1(new_n779), .B2(new_n559), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(G92gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n771), .A2(new_n292), .A3(new_n547), .A4(new_n690), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n788), .A2(new_n799), .ZN(G1337gat));
  INV_X1    g599(.A(G99gat), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n775), .A2(new_n801), .A3(new_n668), .A4(new_n690), .ZN(new_n802));
  OAI21_X1  g601(.A(G99gat), .B1(new_n779), .B2(new_n682), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1338gat));
  OAI21_X1  g603(.A(G106gat), .B1(new_n779), .B2(new_n541), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n541), .A2(G106gat), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n690), .B(new_n806), .C1(new_n782), .C2(new_n783), .ZN(new_n807));
  NAND2_X1  g606(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OR2_X1    g608(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(new_n810), .ZN(G1339gat));
  AOI21_X1  g610(.A(new_n620), .B1(new_n639), .B2(new_n640), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n633), .A2(new_n634), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n631), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT116), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n816), .B(new_n631), .C1(new_n812), .C2(new_n813), .ZN(new_n817));
  AOI221_X4 g616(.A(new_n351), .B1(new_n815), .B2(new_n817), .C1(new_n636), .C2(new_n646), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n332), .A2(new_n333), .A3(new_n348), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n336), .A2(KEYINPUT54), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n343), .B1(new_n349), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n821), .B1(new_n820), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n344), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n636), .A2(new_n646), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n647), .A2(new_n648), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n694), .B1(new_n818), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n826), .B1(new_n319), .B2(new_n320), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n817), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n827), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n250), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n250), .A2(new_n694), .A3(new_n649), .A4(new_n351), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT117), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n827), .A2(new_n690), .A3(new_n832), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n649), .B2(new_n826), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n827), .A2(new_n832), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n840), .A2(new_n694), .B1(new_n841), .B2(new_n831), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n838), .B(new_n835), .C1(new_n842), .C2(new_n250), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n560), .B(new_n540), .C1(new_n837), .C2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n844), .A2(new_n559), .A3(new_n592), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT118), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n450), .A3(new_n650), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n612), .ZN(new_n848));
  OAI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n649), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1340gat));
  NAND3_X1  g649(.A1(new_n846), .A2(new_n460), .A3(new_n690), .ZN(new_n851));
  OAI21_X1  g650(.A(G120gat), .B1(new_n848), .B2(new_n351), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n848), .A2(new_n854), .A3(new_n251), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n845), .A2(new_n250), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n854), .ZN(G1342gat));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  INV_X1    g658(.A(G134gat), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n859), .A3(new_n860), .A4(new_n321), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n844), .A2(new_n860), .A3(new_n559), .A4(new_n592), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT119), .B1(new_n862), .B2(new_n694), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n858), .B1(new_n864), .B2(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n848), .B2(new_n694), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n861), .A2(KEYINPUT120), .A3(new_n863), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n869), .ZN(G1343gat));
  AOI21_X1  g669(.A(new_n541), .B1(new_n837), .B2(new_n843), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n682), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n560), .A3(new_n547), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n834), .A2(new_n836), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n541), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n873), .B(new_n875), .C1(new_n872), .C2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n470), .B1(new_n878), .B2(new_n649), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n871), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n649), .A2(G141gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g682(.A(new_n880), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n468), .A3(new_n690), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n878), .A2(new_n351), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n886), .A2(KEYINPUT59), .A3(new_n468), .ZN(new_n887));
  XNOR2_X1  g686(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n872), .B(new_n541), .C1(new_n837), .C2(new_n843), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n877), .A2(KEYINPUT57), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n690), .A3(new_n875), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n888), .B1(new_n892), .B2(G148gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n885), .B1(new_n887), .B2(new_n893), .ZN(G1345gat));
  AOI21_X1  g693(.A(G155gat), .B1(new_n884), .B2(new_n250), .ZN(new_n895));
  INV_X1    g694(.A(G155gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n878), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n250), .ZN(G1346gat));
  AOI21_X1  g697(.A(G162gat), .B1(new_n884), .B2(new_n321), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n878), .A2(new_n694), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(G162gat), .ZN(G1347gat));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n837), .A2(new_n843), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n560), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT122), .B(new_n606), .C1(new_n837), .C2(new_n843), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n604), .A2(new_n559), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n356), .A3(new_n650), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n606), .B1(new_n837), .B2(new_n843), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n559), .A2(new_n611), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n541), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n649), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n913), .ZN(G1348gat));
  INV_X1    g713(.A(new_n912), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(G176gat), .A3(new_n690), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n690), .B(new_n907), .C1(new_n904), .C2(new_n905), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n917), .A2(new_n918), .A3(new_n341), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n917), .B2(new_n341), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT124), .B(new_n916), .C1(new_n919), .C2(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1349gat));
  OR2_X1    g724(.A1(new_n368), .A2(new_n369), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n906), .A2(new_n926), .A3(new_n250), .A4(new_n907), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n929));
  OAI21_X1  g728(.A(G183gat), .B1(new_n912), .B2(new_n251), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n908), .A2(new_n367), .A3(new_n321), .ZN(new_n934));
  OAI21_X1  g733(.A(G190gat), .B1(new_n912), .B2(new_n694), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1351gat));
  NAND2_X1  g737(.A1(new_n891), .A2(KEYINPUT126), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n874), .A2(new_n606), .A3(new_n559), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT126), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n649), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n874), .A2(new_n559), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n540), .B(new_n944), .C1(new_n904), .C2(new_n905), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(new_n407), .A3(new_n650), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n947), .ZN(G1352gat));
  OR3_X1    g747(.A1(new_n945), .A2(G204gat), .A3(new_n351), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n950));
  OAI21_X1  g749(.A(G204gat), .B1(new_n942), .B2(new_n351), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n946), .A2(new_n245), .A3(new_n250), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n891), .A2(new_n250), .A3(new_n940), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  AOI21_X1  g757(.A(G218gat), .B1(new_n946), .B2(new_n321), .ZN(new_n959));
  INV_X1    g758(.A(new_n942), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n321), .A2(G218gat), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(G1355gat));
endmodule


