//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G120gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(G127gat), .A2(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT69), .B(G127gat), .Z(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT70), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(new_n203), .B2(G120gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n205), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n213), .B(new_n214), .C1(G113gat), .C2(new_n205), .ZN(new_n215));
  NAND2_X1  g014(.A1(G127gat), .A2(G134gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT1), .B1(new_n208), .B2(new_n216), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n215), .A2(KEYINPUT71), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT71), .B1(new_n215), .B2(new_n217), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G141gat), .B(G148gat), .Z(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n221), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G141gat), .B(G148gat), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n225), .B(new_n224), .C1(new_n229), .C2(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n220), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n215), .A2(KEYINPUT71), .A3(new_n217), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n228), .A2(new_n230), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n211), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n232), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G225gat), .A2(G233gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n220), .A2(KEYINPUT80), .A3(new_n231), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n241), .A2(KEYINPUT81), .A3(new_n243), .A4(new_n244), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(KEYINPUT5), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT82), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n247), .A2(KEYINPUT82), .A3(KEYINPUT5), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n239), .A2(KEYINPUT4), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n237), .A2(new_n254), .A3(new_n211), .A4(new_n238), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n237), .A2(new_n211), .B1(KEYINPUT3), .B2(new_n231), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT78), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT78), .B1(new_n231), .B2(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n253), .A2(new_n255), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n262), .A2(KEYINPUT79), .A3(new_n242), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT79), .B1(new_n262), .B2(new_n242), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n251), .A2(new_n252), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT5), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(new_n267), .A3(new_n242), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270));
  INV_X1    g069(.A(G85gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT0), .B(G57gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  XOR2_X1   g073(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n275));
  NAND3_X1  g074(.A1(new_n269), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n274), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n266), .A2(new_n268), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n275), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n266), .B2(new_n268), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G92gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT75), .B(G64gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT27), .B(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n290));
  AOI22_X1  g089(.A1(new_n289), .A2(new_n290), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G169gat), .ZN(new_n295));
  INV_X1    g094(.A(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT26), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n298), .A2(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(KEYINPUT67), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT65), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT68), .B(KEYINPUT26), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n291), .B(new_n294), .C1(new_n300), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n297), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n312), .A2(KEYINPUT25), .A3(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n310), .B(new_n314), .C1(new_n311), .C2(new_n302), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT23), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n318), .B2(new_n309), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G226gat), .ZN(new_n321));
  INV_X1    g120(.A(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G211gat), .B(G218gat), .Z(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  INV_X1    g126(.A(G211gat), .ZN(new_n328));
  INV_X1    g127(.A(G218gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(KEYINPUT22), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n326), .B(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n305), .A2(new_n320), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n321), .B2(new_n322), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n324), .B(new_n332), .C1(new_n334), .C2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n332), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n305), .A2(new_n320), .A3(new_n323), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n305), .B2(new_n320), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n339), .A2(new_n340), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT74), .A3(new_n332), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n286), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(KEYINPUT77), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n345), .A3(new_n286), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT76), .A4(new_n286), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT30), .B1(new_n346), .B2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n349), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n220), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n333), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G227gat), .A2(G233gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G15gat), .B(G43gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G71gat), .B(G99gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  NOR2_X1   g163(.A1(new_n359), .A2(new_n360), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n361), .B(new_n364), .C1(new_n365), .C2(KEYINPUT33), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT33), .ZN(new_n367));
  INV_X1    g166(.A(new_n364), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n359), .B(new_n360), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT32), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT34), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT34), .ZN(new_n373));
  OAI211_X1 g172(.A(KEYINPUT32), .B(new_n373), .C1(new_n359), .C2(new_n360), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n366), .A2(new_n372), .A3(new_n374), .A4(new_n369), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n338), .B1(new_n261), .B2(new_n335), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n380), .ZN(new_n382));
  INV_X1    g181(.A(G228gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n258), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n384));
  AOI211_X1 g183(.A(new_n383), .B(new_n322), .C1(new_n384), .C2(new_n231), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n325), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n331), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n387), .B2(new_n331), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n238), .B1(new_n389), .B2(new_n258), .ZN(new_n390));
  OAI22_X1  g189(.A1(new_n379), .A2(new_n390), .B1(new_n383), .B2(new_n322), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT31), .B(G50gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(G106gat), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT84), .B(G78gat), .Z(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G22gat), .ZN(new_n396));
  INV_X1    g195(.A(G22gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(KEYINPUT86), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n398), .B2(new_n395), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n386), .A2(new_n391), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n386), .B2(new_n391), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n378), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n282), .A2(new_n357), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT35), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n349), .A2(new_n354), .A3(new_n356), .ZN(new_n407));
  NOR4_X1   g206(.A1(new_n378), .A2(new_n407), .A3(new_n403), .A4(KEYINPUT35), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n277), .B1(new_n269), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n266), .A2(KEYINPUT88), .A3(new_n268), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n280), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n276), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n406), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n266), .A2(KEYINPUT88), .A3(new_n268), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT88), .B1(new_n266), .B2(new_n268), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n416), .A2(new_n417), .A3(new_n277), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT40), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n253), .A2(new_n255), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n256), .A2(new_n261), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n242), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT39), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n277), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n243), .B1(new_n241), .B2(new_n244), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n422), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n419), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT87), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n430), .B(new_n419), .C1(new_n425), .C2(new_n427), .ZN(new_n431));
  OR3_X1    g230(.A1(new_n425), .A2(new_n427), .A3(new_n419), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n407), .A2(new_n429), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n402), .B1(new_n418), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n412), .A2(new_n413), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n337), .A2(new_n341), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT37), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n286), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT37), .B1(new_n343), .B2(new_n345), .ZN(new_n440));
  OR3_X1    g239(.A1(new_n439), .A2(KEYINPUT89), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT89), .B1(new_n439), .B2(new_n440), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n347), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT37), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n286), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT90), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n447), .A3(new_n286), .ZN(new_n448));
  INV_X1    g247(.A(new_n440), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT38), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT91), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(KEYINPUT91), .A3(KEYINPUT38), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n443), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n434), .B1(new_n435), .B2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n457));
  NOR2_X1   g256(.A1(new_n378), .A2(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n376), .A2(new_n377), .B1(KEYINPUT72), .B2(KEYINPUT36), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n281), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n278), .A3(new_n279), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n407), .B1(new_n463), .B2(new_n276), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n464), .B2(new_n402), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n415), .B1(new_n456), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G50gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G43gat), .ZN(new_n468));
  INV_X1    g267(.A(G43gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G50gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT15), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT95), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n470), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT15), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(KEYINPUT93), .A2(G36gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n478));
  NAND2_X1  g277(.A1(KEYINPUT93), .A2(G36gat), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n477), .A2(new_n478), .A3(G29gat), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(G29gat), .A3(new_n479), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n483));
  INV_X1    g282(.A(G29gat), .ZN(new_n484));
  INV_X1    g283(.A(G36gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n481), .A2(KEYINPUT94), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n473), .A2(KEYINPUT95), .A3(new_n474), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n476), .A2(new_n480), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT96), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n471), .B1(new_n487), .B2(new_n480), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT15), .B1(new_n468), .B2(new_n470), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(KEYINPUT95), .B2(new_n471), .ZN(new_n494));
  INV_X1    g293(.A(new_n488), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT94), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n486), .A2(new_n482), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n480), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n492), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(KEYINPUT17), .B(new_n491), .C1(new_n501), .C2(new_n490), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n503));
  INV_X1    g302(.A(new_n471), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n490), .B1(new_n489), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT96), .B1(new_n496), .B2(new_n500), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G15gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n397), .ZN(new_n510));
  INV_X1    g309(.A(G1gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(G15gat), .A2(G22gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n510), .A2(new_n512), .B1(KEYINPUT16), .B2(new_n511), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n516), .A2(KEYINPUT98), .ZN(new_n517));
  INV_X1    g316(.A(new_n515), .ZN(new_n518));
  AOI21_X1  g317(.A(G8gat), .B1(new_n518), .B2(KEYINPUT98), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT97), .ZN(new_n520));
  INV_X1    g319(.A(G8gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(KEYINPUT97), .B(G8gat), .C1(new_n514), .C2(new_n515), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n517), .A2(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n502), .A2(new_n508), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n491), .B1(new_n501), .B2(new_n490), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n517), .A2(new_n519), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(new_n523), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n525), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n526), .B(KEYINPUT13), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n506), .A2(new_n507), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(new_n524), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n530), .A2(new_n506), .A3(new_n507), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n526), .A4(new_n531), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n534), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT12), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT100), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n532), .A2(new_n552), .A3(new_n533), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(new_n532), .B2(new_n533), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n541), .A2(new_n540), .A3(new_n548), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n534), .A2(KEYINPUT99), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n532), .A2(new_n552), .A3(new_n533), .ZN(new_n559));
  AND4_X1   g358(.A1(new_n551), .A2(new_n556), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n550), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n271), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n563), .A2(new_n566), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n271), .B2(new_n567), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(new_n571), .A3(new_n566), .A4(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n527), .A2(new_n577), .B1(KEYINPUT41), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n502), .A2(new_n508), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G190gat), .B(G218gat), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT106), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n588));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n585), .B1(KEYINPUT106), .B2(new_n590), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n584), .A2(KEYINPUT107), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n584), .B2(KEYINPUT107), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n592), .A2(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G57gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT102), .B1(new_n598), .B2(G64gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT101), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(G57gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n601), .A3(G57gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(KEYINPUT101), .A3(G64gat), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n599), .A2(new_n602), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G71gat), .A2(G78gat), .ZN(new_n607));
  OR2_X1    g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT9), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n601), .A2(G57gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n598), .A2(G64gat), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT9), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n608), .A2(new_n607), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n606), .A2(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n524), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT105), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT105), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n524), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT104), .B(KEYINPUT19), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n618), .A3(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n631), .A3(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G183gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G211gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n630), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n630), .B2(new_n632), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n597), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT109), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT108), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n570), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n615), .A2(new_n575), .A3(new_n573), .A4(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n606), .A2(new_n610), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n613), .A2(new_n614), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n576), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n642), .B(new_n644), .C1(new_n648), .C2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n644), .B1(new_n648), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT109), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n647), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n577), .A2(KEYINPUT10), .A3(new_n615), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n644), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n654), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT110), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n662), .B(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n641), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n466), .A2(new_n561), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n282), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g471(.A1(new_n669), .A2(new_n407), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n673), .B2(new_n521), .ZN(new_n674));
  NAND2_X1  g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  OR2_X1    g474(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  MUX2_X1   g476(.A(KEYINPUT42), .B(new_n674), .S(new_n677), .Z(G1325gat));
  INV_X1    g477(.A(new_n378), .ZN(new_n679));
  AOI21_X1  g478(.A(G15gat), .B1(new_n669), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n461), .A2(new_n509), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n669), .B2(new_n681), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n669), .A2(new_n403), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT43), .B(G22gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n357), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n410), .A2(new_n411), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n403), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n276), .B1(new_n418), .B2(new_n280), .ZN(new_n691));
  INV_X1    g490(.A(new_n443), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n450), .A2(KEYINPUT91), .A3(KEYINPUT38), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT91), .B1(new_n450), .B2(KEYINPUT38), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n690), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n282), .A2(new_n357), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n460), .B1(new_n697), .B2(new_n403), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n696), .A2(new_n698), .B1(new_n406), .B2(new_n414), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n686), .B1(new_n699), .B2(new_n597), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n466), .A2(KEYINPUT44), .A3(new_n596), .ZN(new_n701));
  INV_X1    g500(.A(new_n640), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n555), .A2(new_n551), .A3(new_n556), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n704), .A2(new_n705), .B1(new_n542), .B2(new_n549), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n667), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n282), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n699), .A2(new_n597), .A3(new_n640), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(new_n707), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n670), .A2(new_n484), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n710), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AND4_X1   g514(.A1(new_n710), .A2(new_n711), .A3(new_n707), .A4(new_n714), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n709), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1328gat));
  NAND2_X1  g518(.A1(new_n477), .A2(new_n479), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n712), .A2(new_n407), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT46), .Z(new_n722));
  NOR2_X1   g521(.A1(new_n708), .A2(new_n357), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(G1329gat));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725));
  OAI21_X1  g524(.A(G43gat), .B1(new_n708), .B2(new_n461), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n712), .A2(new_n469), .A3(new_n679), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1330gat));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n708), .A2(new_n731), .A3(new_n402), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n708), .B2(new_n402), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n732), .A2(G50gat), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n712), .A2(new_n467), .A3(new_n403), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT48), .ZN(new_n736));
  OAI21_X1  g535(.A(G50gat), .B1(new_n708), .B2(new_n402), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n735), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n734), .A2(new_n736), .B1(KEYINPUT48), .B2(new_n738), .ZN(G1331gat));
  INV_X1    g538(.A(new_n667), .ZN(new_n740));
  NOR4_X1   g539(.A1(new_n699), .A2(new_n561), .A3(new_n641), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n670), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g542(.A(new_n357), .B(KEYINPUT114), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT115), .Z(new_n748));
  NOR2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1333gat));
  AOI21_X1  g549(.A(G71gat), .B1(new_n741), .B2(new_n679), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n460), .A2(G71gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n741), .B2(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g553(.A1(new_n741), .A2(new_n403), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n561), .A2(new_n740), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n758), .A2(new_n271), .A3(new_n282), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n699), .A2(new_n597), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n706), .A4(new_n702), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n466), .A2(new_n706), .A3(new_n596), .A4(new_n702), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n740), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n670), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n759), .B1(new_n766), .B2(new_n271), .ZN(G1336gat));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n567), .A3(new_n744), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  OAI21_X1  g568(.A(G92gat), .B1(new_n758), .B2(new_n745), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G92gat), .B1(new_n758), .B2(new_n357), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT116), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(G92gat), .C1(new_n758), .C2(new_n357), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n773), .A2(new_n768), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n771), .B1(new_n776), .B2(new_n769), .ZN(G1337gat));
  INV_X1    g576(.A(G99gat), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n758), .A2(new_n778), .A3(new_n461), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n765), .A2(new_n679), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n778), .ZN(G1338gat));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n758), .B2(new_n402), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT117), .B1(new_n758), .B2(new_n402), .ZN(new_n785));
  INV_X1    g584(.A(G106gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI211_X1 g586(.A(new_n402), .B(new_n740), .C1(new_n761), .C2(new_n764), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(KEYINPUT53), .B(new_n784), .C1(new_n787), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1339gat));
  NAND2_X1  g592(.A1(new_n668), .A2(new_n706), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n704), .A2(new_n705), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n661), .A2(new_n666), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n658), .A2(new_n659), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n643), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n658), .A2(new_n644), .A3(new_n659), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n666), .B1(new_n660), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT55), .B1(new_n801), .B2(new_n803), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n797), .B(new_n804), .C1(new_n805), .C2(KEYINPUT118), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n658), .A2(new_n644), .A3(new_n659), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(new_n660), .A3(new_n802), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n798), .A2(new_n802), .A3(new_n643), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n665), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n796), .B1(new_n806), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n797), .A2(new_n804), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n805), .A2(KEYINPUT118), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT119), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n547), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n538), .A2(new_n539), .A3(new_n536), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n526), .B1(new_n525), .B2(new_n531), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND4_X1   g623(.A1(new_n795), .A2(new_n820), .A3(new_n596), .A4(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n667), .B(new_n824), .C1(new_n557), .C2(new_n560), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n815), .A2(new_n819), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n706), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n825), .B1(new_n828), .B2(new_n597), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n794), .B1(new_n829), .B2(new_n640), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n404), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n831), .A2(new_n282), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n745), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n706), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(new_n203), .ZN(G1340gat));
  NOR2_X1   g635(.A1(new_n834), .A2(new_n740), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(new_n205), .ZN(G1341gat));
  NOR2_X1   g637(.A1(new_n834), .A2(new_n702), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(new_n210), .ZN(G1342gat));
  NOR2_X1   g639(.A1(new_n597), .A2(new_n407), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n833), .A2(new_n209), .A3(new_n841), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n842), .B(KEYINPUT56), .Z(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n834), .B2(new_n597), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1343gat));
  AND2_X1   g644(.A1(new_n795), .A2(new_n824), .ZN(new_n846));
  INV_X1    g645(.A(new_n816), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n801), .A2(KEYINPUT120), .A3(new_n803), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT120), .B1(new_n801), .B2(new_n803), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(KEYINPUT55), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n846), .A2(new_n667), .B1(new_n561), .B2(new_n851), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(new_n596), .ZN(new_n853));
  INV_X1    g652(.A(new_n825), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n855), .A2(new_n702), .B1(new_n706), .B2(new_n668), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n402), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n831), .A2(new_n402), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n461), .A2(new_n670), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n744), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G141gat), .B1(new_n863), .B2(new_n706), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n858), .A2(new_n862), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n865), .A2(G141gat), .A3(new_n706), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n864), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1344gat));
  OR3_X1    g670(.A1(new_n865), .A2(G148gat), .A3(new_n740), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n806), .A2(new_n814), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n846), .A2(new_n596), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n853), .A2(KEYINPUT121), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n702), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT121), .B1(new_n853), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n794), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n859), .A3(new_n403), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT57), .B1(new_n831), .B2(new_n402), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n667), .A3(new_n862), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n873), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n873), .A2(G148gat), .ZN(new_n884));
  INV_X1    g683(.A(new_n863), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n667), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n872), .B1(new_n883), .B2(new_n886), .ZN(G1345gat));
  INV_X1    g686(.A(new_n865), .ZN(new_n888));
  AOI21_X1  g687(.A(G155gat), .B1(new_n888), .B2(new_n640), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n702), .A2(new_n222), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n885), .B2(new_n890), .ZN(G1346gat));
  OAI21_X1  g690(.A(G162gat), .B1(new_n863), .B2(new_n597), .ZN(new_n892));
  INV_X1    g691(.A(new_n861), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n858), .A2(new_n223), .A3(new_n841), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n892), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1347gat));
  NAND2_X1  g698(.A1(new_n561), .A2(new_n820), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n596), .B1(new_n900), .B2(new_n826), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n702), .B1(new_n901), .B2(new_n825), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n670), .B1(new_n902), .B2(new_n794), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n404), .A3(new_n744), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n295), .A3(new_n561), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n830), .A2(new_n282), .A3(new_n407), .A4(new_n404), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT123), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n903), .A2(new_n909), .A3(new_n407), .A4(new_n404), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(new_n561), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n906), .B1(new_n912), .B2(new_n295), .ZN(G1348gat));
  AOI21_X1  g712(.A(G176gat), .B1(new_n905), .B2(new_n667), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n740), .A2(new_n296), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n911), .B2(new_n915), .ZN(G1349gat));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n908), .A2(new_n640), .A3(new_n910), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G183gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n830), .A2(new_n282), .A3(new_n404), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n640), .A2(new_n287), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n921), .A2(new_n745), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT125), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n920), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n918), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n920), .B2(new_n924), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT125), .B(new_n923), .C1(new_n919), .C2(G183gat), .ZN(new_n931));
  INV_X1    g730(.A(new_n918), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n929), .A2(new_n933), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n905), .A2(new_n288), .A3(new_n596), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n911), .A2(new_n596), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(G190gat), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT61), .B(new_n288), .C1(new_n911), .C2(new_n596), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1351gat));
  NAND4_X1  g739(.A1(new_n903), .A2(new_n403), .A3(new_n461), .A4(new_n744), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT126), .ZN(new_n942));
  XOR2_X1   g741(.A(KEYINPUT127), .B(G197gat), .Z(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n561), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n880), .A2(new_n881), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n670), .A2(new_n460), .A3(new_n357), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n946), .A2(new_n706), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n949), .B2(new_n944), .ZN(G1352gat));
  NOR3_X1   g749(.A1(new_n941), .A2(G204gat), .A3(new_n740), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n946), .A2(new_n740), .A3(new_n948), .ZN(new_n953));
  INV_X1    g752(.A(G204gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n942), .A2(new_n328), .A3(new_n640), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n880), .A2(new_n640), .A3(new_n881), .A4(new_n947), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  NOR4_X1   g759(.A1(new_n946), .A2(new_n329), .A3(new_n597), .A4(new_n948), .ZN(new_n961));
  AOI21_X1  g760(.A(G218gat), .B1(new_n942), .B2(new_n596), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(G1355gat));
endmodule


