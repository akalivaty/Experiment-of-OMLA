

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779;

  AND2_X1 U375 ( .A1(n437), .A2(n356), .ZN(n435) );
  OR2_X1 U376 ( .A1(n657), .A2(n438), .ZN(n437) );
  XNOR2_X1 U377 ( .A(n476), .B(n475), .ZN(n497) );
  NOR2_X1 U378 ( .A1(n694), .A2(n682), .ZN(n431) );
  XNOR2_X1 U379 ( .A(n431), .B(KEYINPUT100), .ZN(n563) );
  XNOR2_X2 U380 ( .A(n386), .B(n365), .ZN(n368) );
  XNOR2_X2 U381 ( .A(n494), .B(n493), .ZN(n708) );
  XNOR2_X2 U382 ( .A(n715), .B(KEYINPUT6), .ZN(n583) );
  AND2_X1 U383 ( .A1(n736), .A2(KEYINPUT2), .ZN(n637) );
  INV_X1 U384 ( .A(G953), .ZN(n769) );
  XNOR2_X1 U385 ( .A(G140), .B(G131), .ZN(n522) );
  NAND2_X1 U386 ( .A1(n385), .A2(n631), .ZN(n739) );
  NOR2_X1 U387 ( .A1(n613), .A2(n612), .ZN(n370) );
  NAND2_X1 U388 ( .A1(n399), .A2(n395), .ZN(n647) );
  XNOR2_X1 U389 ( .A(n430), .B(n429), .ZN(n778) );
  AND2_X1 U390 ( .A1(n417), .A2(n414), .ZN(n413) );
  OR2_X1 U391 ( .A1(n630), .A2(n618), .ZN(n430) );
  NOR2_X1 U392 ( .A1(n620), .A2(n595), .ZN(n689) );
  AND2_X1 U393 ( .A1(n409), .A2(n408), .ZN(n407) );
  XNOR2_X1 U394 ( .A(n664), .B(n663), .ZN(n665) );
  OR2_X1 U395 ( .A1(n523), .A2(n359), .ZN(n422) );
  XNOR2_X1 U396 ( .A(n448), .B(G146), .ZN(n503) );
  XNOR2_X1 U397 ( .A(G101), .B(KEYINPUT79), .ZN(n475) );
  NAND2_X1 U398 ( .A1(n413), .A2(n411), .ZN(n367) );
  XNOR2_X2 U399 ( .A(n353), .B(n489), .ZN(n672) );
  AND2_X2 U400 ( .A1(n432), .A2(n715), .ZN(n682) );
  BUF_X1 U401 ( .A(n650), .Z(n352) );
  BUF_X1 U402 ( .A(n384), .Z(n353) );
  INV_X1 U403 ( .A(n572), .ZN(n354) );
  XNOR2_X1 U404 ( .A(n384), .B(n478), .ZN(n650) );
  XNOR2_X1 U405 ( .A(n767), .B(G146), .ZN(n384) );
  XNOR2_X2 U406 ( .A(n592), .B(n480), .ZN(n547) );
  XNOR2_X1 U407 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U408 ( .A(n503), .B(n449), .ZN(n523) );
  INV_X1 U409 ( .A(KEYINPUT10), .ZN(n449) );
  NAND2_X1 U410 ( .A1(n439), .A2(n507), .ZN(n438) );
  INV_X1 U411 ( .A(n510), .ZN(n439) );
  XNOR2_X1 U412 ( .A(G478), .B(n537), .ZN(n560) );
  NOR2_X1 U413 ( .A1(n750), .A2(G902), .ZN(n537) );
  XNOR2_X1 U414 ( .A(n705), .B(n374), .ZN(n597) );
  INV_X1 U415 ( .A(KEYINPUT86), .ZN(n374) );
  OR2_X1 U416 ( .A1(n647), .A2(n646), .ZN(n574) );
  INV_X1 U417 ( .A(KEYINPUT96), .ZN(n428) );
  NAND2_X1 U418 ( .A1(KEYINPUT23), .A2(n428), .ZN(n426) );
  NAND2_X1 U419 ( .A1(n425), .A2(n424), .ZN(n423) );
  NAND2_X1 U420 ( .A1(KEYINPUT96), .A2(KEYINPUT23), .ZN(n425) );
  NAND2_X1 U421 ( .A1(n428), .A2(n450), .ZN(n424) );
  XNOR2_X1 U422 ( .A(n394), .B(n392), .ZN(n532) );
  XNOR2_X1 U423 ( .A(KEYINPUT8), .B(KEYINPUT72), .ZN(n394) );
  NOR2_X1 U424 ( .A1(n393), .A2(G953), .ZN(n392) );
  INV_X1 U425 ( .A(G234), .ZN(n393) );
  NOR2_X1 U426 ( .A1(G953), .A2(G237), .ZN(n526) );
  NAND2_X1 U427 ( .A1(n371), .A2(n369), .ZN(n419) );
  AND2_X1 U428 ( .A1(n420), .A2(n697), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n370), .B(KEYINPUT76), .ZN(n369) );
  NAND2_X1 U430 ( .A1(n558), .A2(n416), .ZN(n415) );
  INV_X1 U431 ( .A(n443), .ZN(n416) );
  NAND2_X1 U432 ( .A1(n479), .A2(n509), .ZN(n406) );
  INV_X1 U433 ( .A(G134), .ZN(n433) );
  XNOR2_X1 U434 ( .A(n536), .B(n404), .ZN(n403) );
  INV_X1 U435 ( .A(KEYINPUT9), .ZN(n404) );
  XNOR2_X1 U436 ( .A(G116), .B(G107), .ZN(n536) );
  NOR2_X1 U437 ( .A1(n739), .A2(n507), .ZN(n379) );
  XNOR2_X1 U438 ( .A(G104), .B(G122), .ZN(n524) );
  XNOR2_X1 U439 ( .A(G113), .B(G143), .ZN(n528) );
  INV_X1 U440 ( .A(G125), .ZN(n448) );
  XNOR2_X1 U441 ( .A(n496), .B(n495), .ZN(n376) );
  XNOR2_X1 U442 ( .A(KEYINPUT16), .B(G122), .ZN(n495) );
  XNOR2_X1 U443 ( .A(n619), .B(n366), .ZN(n724) );
  INV_X1 U444 ( .A(KEYINPUT41), .ZN(n366) );
  INV_X1 U445 ( .A(n691), .ZN(n618) );
  NAND2_X1 U446 ( .A1(n398), .A2(n397), .ZN(n396) );
  NAND2_X1 U447 ( .A1(n355), .A2(n363), .ZN(n400) );
  XNOR2_X1 U448 ( .A(n373), .B(n372), .ZN(n562) );
  XNOR2_X1 U449 ( .A(KEYINPUT13), .B(G475), .ZN(n372) );
  OR2_X1 U450 ( .A1(n664), .A2(G902), .ZN(n373) );
  NOR2_X1 U451 ( .A1(n558), .A2(n544), .ZN(n546) );
  INV_X1 U452 ( .A(G237), .ZN(n508) );
  NAND2_X1 U453 ( .A1(n410), .A2(G902), .ZN(n408) );
  XNOR2_X1 U454 ( .A(n502), .B(n469), .ZN(n470) );
  XNOR2_X1 U455 ( .A(G137), .B(KEYINPUT73), .ZN(n469) );
  NAND2_X1 U456 ( .A1(G237), .A2(G234), .ZN(n514) );
  OR2_X1 U457 ( .A1(n691), .A2(n693), .ZN(n705) );
  AND2_X1 U458 ( .A1(n562), .A2(n560), .ZN(n703) );
  NAND2_X1 U459 ( .A1(n510), .A2(n632), .ZN(n440) );
  XNOR2_X1 U460 ( .A(G101), .B(G131), .ZN(n485) );
  XOR2_X1 U461 ( .A(KEYINPUT5), .B(KEYINPUT78), .Z(n483) );
  XOR2_X1 U462 ( .A(KEYINPUT24), .B(G140), .Z(n456) );
  XNOR2_X1 U463 ( .A(G119), .B(G110), .ZN(n455) );
  NAND2_X1 U464 ( .A1(n523), .A2(n423), .ZN(n421) );
  INV_X1 U465 ( .A(KEYINPUT81), .ZN(n451) );
  XNOR2_X1 U466 ( .A(n389), .B(G137), .ZN(n452) );
  XNOR2_X1 U467 ( .A(n633), .B(KEYINPUT70), .ZN(n634) );
  XNOR2_X1 U468 ( .A(n419), .B(n364), .ZN(n385) );
  AND2_X1 U469 ( .A1(n415), .A2(n540), .ZN(n414) );
  NAND2_X1 U470 ( .A1(n412), .A2(n416), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n535), .B(n402), .ZN(n750) );
  XOR2_X1 U472 ( .A(G122), .B(KEYINPUT7), .Z(n534) );
  XNOR2_X1 U473 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U474 ( .A(n754), .B(n506), .ZN(n657) );
  AND2_X1 U475 ( .A1(n641), .A2(G953), .ZN(n753) );
  NOR2_X1 U476 ( .A1(n724), .A2(n620), .ZN(n622) );
  XNOR2_X1 U477 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n429) );
  OR2_X1 U478 ( .A1(n551), .A2(n362), .ZN(n395) );
  AND2_X1 U479 ( .A1(n401), .A2(n400), .ZN(n399) );
  BUF_X1 U480 ( .A(G128), .Z(n389) );
  NOR2_X1 U481 ( .A1(n562), .A2(n561), .ZN(n691) );
  OR2_X1 U482 ( .A1(n549), .A2(n583), .ZN(n355) );
  AND2_X1 U483 ( .A1(n440), .A2(n436), .ZN(n356) );
  NOR2_X1 U484 ( .A1(n702), .A2(n701), .ZN(n357) );
  AND2_X1 U485 ( .A1(n556), .A2(n443), .ZN(n358) );
  AND2_X1 U486 ( .A1(n427), .A2(n426), .ZN(n359) );
  OR2_X1 U487 ( .A1(n576), .A2(n575), .ZN(n360) );
  AND2_X1 U488 ( .A1(n437), .A2(n440), .ZN(n361) );
  OR2_X1 U489 ( .A1(n549), .A2(n396), .ZN(n362) );
  XOR2_X1 U490 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n363) );
  XOR2_X1 U491 ( .A(KEYINPUT74), .B(KEYINPUT48), .Z(n364) );
  XNOR2_X1 U492 ( .A(n376), .B(n497), .ZN(n754) );
  INV_X1 U493 ( .A(n507), .ZN(n632) );
  XNOR2_X1 U494 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n365) );
  NAND2_X2 U495 ( .A1(n407), .A2(n405), .ZN(n592) );
  OR2_X1 U496 ( .A1(n650), .A2(n406), .ZN(n405) );
  NAND2_X1 U497 ( .A1(n368), .A2(n379), .ZN(n635) );
  OR2_X2 U498 ( .A1(n669), .A2(KEYINPUT89), .ZN(n391) );
  XNOR2_X2 U499 ( .A(n367), .B(n542), .ZN(n669) );
  INV_X1 U500 ( .A(n368), .ZN(n738) );
  AND2_X1 U501 ( .A1(n368), .A2(n375), .ZN(n736) );
  INV_X1 U502 ( .A(n693), .ZN(n629) );
  NOR2_X1 U503 ( .A1(n597), .A2(KEYINPUT47), .ZN(n598) );
  INV_X1 U504 ( .A(n739), .ZN(n375) );
  XNOR2_X2 U505 ( .A(G107), .B(G104), .ZN(n474) );
  XNOR2_X2 U506 ( .A(n377), .B(KEYINPUT0), .ZN(n558) );
  NAND2_X1 U507 ( .A1(n594), .A2(n521), .ZN(n377) );
  XNOR2_X2 U508 ( .A(n378), .B(n513), .ZN(n594) );
  NAND2_X1 U509 ( .A1(n435), .A2(n441), .ZN(n378) );
  XNOR2_X2 U510 ( .A(n380), .B(n470), .ZN(n767) );
  XNOR2_X1 U511 ( .A(n380), .B(n403), .ZN(n402) );
  XNOR2_X2 U512 ( .A(n498), .B(n433), .ZN(n380) );
  XNOR2_X2 U513 ( .A(n382), .B(n381), .ZN(n496) );
  XNOR2_X2 U514 ( .A(KEYINPUT3), .B(G119), .ZN(n381) );
  XNOR2_X2 U515 ( .A(G116), .B(G113), .ZN(n382) );
  AND2_X1 U516 ( .A1(n383), .A2(n590), .ZN(n722) );
  XNOR2_X2 U517 ( .A(n481), .B(KEYINPUT77), .ZN(n383) );
  NAND2_X1 U518 ( .A1(n383), .A2(n583), .ZN(n494) );
  NAND2_X1 U519 ( .A1(n387), .A2(n360), .ZN(n386) );
  XNOR2_X1 U520 ( .A(n571), .B(n388), .ZN(n387) );
  INV_X1 U521 ( .A(KEYINPUT88), .ZN(n388) );
  INV_X2 U522 ( .A(G128), .ZN(n434) );
  NAND2_X1 U523 ( .A1(n669), .A2(n447), .ZN(n390) );
  NOR2_X2 U524 ( .A1(n563), .A2(n597), .ZN(n564) );
  XNOR2_X2 U525 ( .A(n557), .B(KEYINPUT31), .ZN(n694) );
  NAND2_X1 U526 ( .A1(n391), .A2(n390), .ZN(n442) );
  INV_X1 U527 ( .A(n363), .ZN(n397) );
  INV_X1 U528 ( .A(n583), .ZN(n398) );
  NAND2_X1 U529 ( .A1(n551), .A2(n363), .ZN(n401) );
  OR2_X1 U530 ( .A1(n551), .A2(n583), .ZN(n567) );
  NAND2_X1 U531 ( .A1(n650), .A2(n410), .ZN(n409) );
  NAND2_X1 U532 ( .A1(n547), .A2(n418), .ZN(n481) );
  INV_X1 U533 ( .A(n479), .ZN(n410) );
  INV_X1 U534 ( .A(n708), .ZN(n412) );
  NAND2_X1 U535 ( .A1(n708), .A2(n358), .ZN(n417) );
  NAND2_X1 U536 ( .A1(n418), .A2(n592), .ZN(n602) );
  NOR2_X1 U537 ( .A1(n716), .A2(n418), .ZN(n717) );
  NOR2_X2 U538 ( .A1(n548), .A2(n543), .ZN(n418) );
  XNOR2_X1 U539 ( .A(n623), .B(KEYINPUT46), .ZN(n420) );
  NAND2_X1 U540 ( .A1(n422), .A2(n421), .ZN(n454) );
  NAND2_X1 U541 ( .A1(n450), .A2(KEYINPUT96), .ZN(n427) );
  XNOR2_X1 U542 ( .A(n559), .B(KEYINPUT98), .ZN(n432) );
  XNOR2_X2 U543 ( .A(n434), .B(G143), .ZN(n498) );
  NAND2_X1 U544 ( .A1(n441), .A2(n361), .ZN(n615) );
  INV_X1 U545 ( .A(n701), .ZN(n436) );
  NAND2_X1 U546 ( .A1(n657), .A2(n510), .ZN(n441) );
  BUF_X1 U547 ( .A(n547), .Z(n716) );
  XNOR2_X1 U548 ( .A(n454), .B(n453), .ZN(n460) );
  AND2_X1 U549 ( .A1(n548), .A2(n582), .ZN(n589) );
  NOR2_X4 U550 ( .A1(n638), .A2(n637), .ZN(n748) );
  XNOR2_X2 U551 ( .A(n636), .B(KEYINPUT65), .ZN(n638) );
  XOR2_X1 U552 ( .A(KEYINPUT84), .B(KEYINPUT34), .Z(n443) );
  XOR2_X1 U553 ( .A(n545), .B(KEYINPUT22), .Z(n444) );
  AND2_X1 U554 ( .A1(n526), .A2(G214), .ZN(n445) );
  OR2_X1 U555 ( .A1(KEYINPUT44), .A2(KEYINPUT89), .ZN(n446) );
  AND2_X1 U556 ( .A1(KEYINPUT44), .A2(KEYINPUT89), .ZN(n447) );
  INV_X1 U557 ( .A(n574), .ZN(n554) );
  INV_X1 U558 ( .A(KEYINPUT99), .ZN(n484) );
  XNOR2_X1 U559 ( .A(n485), .B(n484), .ZN(n486) );
  NOR2_X1 U560 ( .A1(n603), .A2(n543), .ZN(n582) );
  XNOR2_X1 U561 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U562 ( .A(n527), .B(n445), .ZN(n530) );
  XNOR2_X1 U563 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U564 ( .A1(n616), .A2(n702), .ZN(n617) );
  INV_X1 U565 ( .A(KEYINPUT23), .ZN(n450) );
  NAND2_X1 U566 ( .A1(n532), .A2(G221), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U568 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U569 ( .A(n460), .B(n459), .ZN(n639) );
  INV_X1 U570 ( .A(G902), .ZN(n509) );
  NAND2_X1 U571 ( .A1(n639), .A2(n509), .ZN(n465) );
  XOR2_X1 U572 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n463) );
  XNOR2_X1 U573 ( .A(G902), .B(KEYINPUT15), .ZN(n507) );
  NAND2_X1 U574 ( .A1(n507), .A2(G234), .ZN(n461) );
  XNOR2_X1 U575 ( .A(n461), .B(KEYINPUT20), .ZN(n466) );
  NAND2_X1 U576 ( .A1(n466), .A2(G217), .ZN(n462) );
  XNOR2_X1 U577 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X2 U578 ( .A(n465), .B(n464), .ZN(n548) );
  AND2_X1 U579 ( .A1(n466), .A2(G221), .ZN(n468) );
  INV_X1 U580 ( .A(KEYINPUT21), .ZN(n467) );
  XNOR2_X1 U581 ( .A(n468), .B(n467), .ZN(n543) );
  XNOR2_X2 U582 ( .A(KEYINPUT71), .B(KEYINPUT4), .ZN(n502) );
  INV_X1 U583 ( .A(n522), .ZN(n471) );
  XOR2_X1 U584 ( .A(n471), .B(KEYINPUT82), .Z(n473) );
  NAND2_X1 U585 ( .A1(G227), .A2(n769), .ZN(n472) );
  XNOR2_X1 U586 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U587 ( .A(n474), .B(G110), .ZN(n476) );
  XNOR2_X1 U588 ( .A(n477), .B(n497), .ZN(n478) );
  XNOR2_X1 U589 ( .A(KEYINPUT75), .B(G469), .ZN(n479) );
  XNOR2_X1 U590 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n480) );
  NAND2_X1 U591 ( .A1(n526), .A2(G210), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n483), .B(n482), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n496), .B(n488), .ZN(n489) );
  NAND2_X1 U594 ( .A1(n672), .A2(n509), .ZN(n491) );
  INV_X1 U595 ( .A(G472), .ZN(n490) );
  XNOR2_X2 U596 ( .A(n491), .B(n490), .ZN(n715) );
  INV_X1 U597 ( .A(KEYINPUT103), .ZN(n492) );
  XNOR2_X1 U598 ( .A(n492), .B(KEYINPUT33), .ZN(n493) );
  XNOR2_X1 U599 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n500) );
  NAND2_X1 U600 ( .A1(n769), .A2(G224), .ZN(n499) );
  XNOR2_X1 U601 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U602 ( .A(n498), .B(n501), .ZN(n505) );
  XNOR2_X1 U603 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U604 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U605 ( .A1(n509), .A2(n508), .ZN(n511) );
  NAND2_X1 U606 ( .A1(n511), .A2(G210), .ZN(n510) );
  NAND2_X1 U607 ( .A1(n511), .A2(G214), .ZN(n512) );
  XNOR2_X1 U608 ( .A(n512), .B(KEYINPUT93), .ZN(n701) );
  XNOR2_X1 U609 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n513) );
  XNOR2_X1 U610 ( .A(n514), .B(KEYINPUT14), .ZN(n516) );
  NAND2_X1 U611 ( .A1(G952), .A2(n516), .ZN(n515) );
  XNOR2_X1 U612 ( .A(KEYINPUT94), .B(n515), .ZN(n731) );
  NOR2_X1 U613 ( .A1(G953), .A2(n731), .ZN(n581) );
  NAND2_X1 U614 ( .A1(G902), .A2(n516), .ZN(n577) );
  INV_X1 U615 ( .A(n577), .ZN(n517) );
  NOR2_X1 U616 ( .A1(G898), .A2(n769), .ZN(n755) );
  AND2_X1 U617 ( .A1(n517), .A2(n755), .ZN(n518) );
  OR2_X1 U618 ( .A1(n581), .A2(n518), .ZN(n520) );
  INV_X1 U619 ( .A(KEYINPUT95), .ZN(n519) );
  XNOR2_X1 U620 ( .A(n520), .B(n519), .ZN(n521) );
  INV_X1 U621 ( .A(n558), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n523), .B(n522), .ZN(n766) );
  XOR2_X1 U623 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n525) );
  XNOR2_X1 U624 ( .A(n525), .B(n524), .ZN(n527) );
  XNOR2_X1 U625 ( .A(n528), .B(KEYINPUT11), .ZN(n529) );
  XNOR2_X1 U626 ( .A(n766), .B(n531), .ZN(n664) );
  NAND2_X1 U627 ( .A1(G217), .A2(n532), .ZN(n533) );
  XNOR2_X1 U628 ( .A(n534), .B(n533), .ZN(n535) );
  NOR2_X1 U629 ( .A1(n562), .A2(n560), .ZN(n539) );
  INV_X1 U630 ( .A(KEYINPUT104), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n539), .B(n538), .ZN(n608) );
  INV_X1 U632 ( .A(n608), .ZN(n540) );
  INV_X1 U633 ( .A(KEYINPUT83), .ZN(n541) );
  XNOR2_X1 U634 ( .A(n541), .B(KEYINPUT35), .ZN(n542) );
  INV_X1 U635 ( .A(n543), .ZN(n712) );
  NAND2_X1 U636 ( .A1(n703), .A2(n712), .ZN(n544) );
  INV_X1 U637 ( .A(KEYINPUT67), .ZN(n545) );
  XNOR2_X1 U638 ( .A(n546), .B(n444), .ZN(n551) );
  NAND2_X1 U639 ( .A1(n716), .A2(n548), .ZN(n549) );
  INV_X1 U640 ( .A(n548), .ZN(n711) );
  OR2_X1 U641 ( .A1(n716), .A2(n711), .ZN(n550) );
  INV_X1 U642 ( .A(n715), .ZN(n590) );
  NOR2_X1 U643 ( .A1(n550), .A2(n590), .ZN(n553) );
  INV_X1 U644 ( .A(n551), .ZN(n552) );
  AND2_X1 U645 ( .A1(n553), .A2(n552), .ZN(n646) );
  NAND2_X1 U646 ( .A1(n442), .A2(n554), .ZN(n555) );
  NAND2_X1 U647 ( .A1(n555), .A2(n446), .ZN(n570) );
  NAND2_X1 U648 ( .A1(n722), .A2(n556), .ZN(n557) );
  NOR2_X1 U649 ( .A1(n602), .A2(n558), .ZN(n559) );
  INV_X1 U650 ( .A(n560), .ZN(n561) );
  AND2_X1 U651 ( .A1(n562), .A2(n561), .ZN(n693) );
  XNOR2_X1 U652 ( .A(n564), .B(KEYINPUT102), .ZN(n568) );
  INV_X1 U653 ( .A(n716), .ZN(n565) );
  NAND2_X1 U654 ( .A1(n565), .A2(n711), .ZN(n566) );
  NOR2_X1 U655 ( .A1(n567), .A2(n566), .ZN(n678) );
  NOR2_X1 U656 ( .A1(n568), .A2(n678), .ZN(n569) );
  NAND2_X1 U657 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U658 ( .A(n669), .ZN(n572) );
  INV_X1 U659 ( .A(KEYINPUT44), .ZN(n573) );
  NAND2_X1 U660 ( .A1(n572), .A2(n573), .ZN(n576) );
  XNOR2_X1 U661 ( .A(n574), .B(KEYINPUT90), .ZN(n575) );
  NOR2_X1 U662 ( .A1(G900), .A2(n577), .ZN(n578) );
  NAND2_X1 U663 ( .A1(G953), .A2(n578), .ZN(n579) );
  XNOR2_X1 U664 ( .A(KEYINPUT105), .B(n579), .ZN(n580) );
  NOR2_X1 U665 ( .A1(n581), .A2(n580), .ZN(n603) );
  NAND2_X1 U666 ( .A1(n583), .A2(n589), .ZN(n584) );
  NOR2_X1 U667 ( .A1(n618), .A2(n584), .ZN(n585) );
  XNOR2_X1 U668 ( .A(n585), .B(KEYINPUT106), .ZN(n586) );
  NAND2_X1 U669 ( .A1(n586), .A2(n436), .ZN(n624) );
  NOR2_X1 U670 ( .A1(n624), .A2(n615), .ZN(n587) );
  XNOR2_X1 U671 ( .A(n587), .B(KEYINPUT36), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n588), .A2(n716), .ZN(n697) );
  AND2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U674 ( .A(KEYINPUT28), .B(n591), .ZN(n593) );
  NAND2_X1 U675 ( .A1(n593), .A2(n592), .ZN(n620) );
  INV_X1 U676 ( .A(n594), .ZN(n595) );
  INV_X1 U677 ( .A(KEYINPUT47), .ZN(n610) );
  NOR2_X1 U678 ( .A1(n689), .A2(n610), .ZN(n596) );
  XNOR2_X1 U679 ( .A(n596), .B(KEYINPUT85), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n689), .A2(n598), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n613) );
  INV_X1 U682 ( .A(n615), .ZN(n626) );
  NOR2_X1 U683 ( .A1(n701), .A2(n715), .ZN(n601) );
  XNOR2_X1 U684 ( .A(KEYINPUT30), .B(n601), .ZN(n605) );
  NOR2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n616) );
  INV_X1 U687 ( .A(n616), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n626), .A2(n606), .ZN(n607) );
  OR2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U690 ( .A(KEYINPUT108), .B(n609), .ZN(n779) );
  OR2_X1 U691 ( .A1(n705), .A2(n610), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n779), .A2(n611), .ZN(n612) );
  INV_X1 U693 ( .A(KEYINPUT38), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n615), .B(n614), .ZN(n702) );
  XNOR2_X1 U695 ( .A(n617), .B(KEYINPUT39), .ZN(n630) );
  NAND2_X1 U696 ( .A1(n357), .A2(n703), .ZN(n619) );
  XNOR2_X1 U697 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n622), .B(n621), .ZN(n776) );
  NOR2_X1 U699 ( .A1(n778), .A2(n776), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n716), .A2(n624), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n625), .B(KEYINPUT43), .ZN(n627) );
  NOR2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT107), .ZN(n777) );
  OR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n698) );
  AND2_X1 U705 ( .A1(n777), .A2(n698), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n748), .A2(G217), .ZN(n640) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n642) );
  INV_X1 U710 ( .A(G952), .ZN(n641) );
  INV_X1 U711 ( .A(n753), .ZN(n675) );
  NAND2_X1 U712 ( .A1(n642), .A2(n675), .ZN(n644) );
  INV_X1 U713 ( .A(KEYINPUT122), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(G66) );
  XNOR2_X1 U715 ( .A(G110), .B(KEYINPUT114), .ZN(n645) );
  XOR2_X1 U716 ( .A(n646), .B(n645), .Z(G12) );
  XOR2_X1 U717 ( .A(G119), .B(KEYINPUT127), .Z(n648) );
  XOR2_X1 U718 ( .A(n648), .B(n647), .Z(G21) );
  NAND2_X1 U719 ( .A1(n748), .A2(G469), .ZN(n652) );
  XOR2_X1 U720 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n649) );
  XNOR2_X1 U721 ( .A(n352), .B(n649), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X2 U723 ( .A1(n653), .A2(n753), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n654), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U725 ( .A1(n748), .A2(G210), .ZN(n659) );
  XNOR2_X1 U726 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n655), .B(KEYINPUT55), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X2 U729 ( .A1(n660), .A2(n753), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U731 ( .A1(n748), .A2(G475), .ZN(n666) );
  XOR2_X1 U732 ( .A(KEYINPUT69), .B(KEYINPUT121), .Z(n662) );
  XNOR2_X1 U733 ( .A(n662), .B(KEYINPUT59), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X2 U735 ( .A1(n667), .A2(n753), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n668), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U737 ( .A(n354), .B(G122), .Z(G24) );
  NAND2_X1 U738 ( .A1(n748), .A2(G472), .ZN(n674) );
  XNOR2_X1 U739 ( .A(KEYINPUT92), .B(KEYINPUT111), .ZN(n670) );
  XOR2_X1 U740 ( .A(n670), .B(KEYINPUT62), .Z(n671) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n677), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U745 ( .A(G101), .B(n678), .Z(n679) );
  XNOR2_X1 U746 ( .A(KEYINPUT112), .B(n679), .ZN(G3) );
  XOR2_X1 U747 ( .A(G104), .B(KEYINPUT113), .Z(n681) );
  NAND2_X1 U748 ( .A1(n682), .A2(n691), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(G6) );
  XOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n684) );
  NAND2_X1 U751 ( .A1(n682), .A2(n693), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U753 ( .A(G107), .B(n685), .ZN(G9) );
  XOR2_X1 U754 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n687) );
  NAND2_X1 U755 ( .A1(n689), .A2(n693), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n687), .B(n686), .ZN(n688) );
  XOR2_X1 U757 ( .A(n389), .B(n688), .Z(G30) );
  NAND2_X1 U758 ( .A1(n689), .A2(n691), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n690), .B(G146), .ZN(G48) );
  NAND2_X1 U760 ( .A1(n694), .A2(n691), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(G113), .ZN(G15) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U763 ( .A(n695), .B(G116), .ZN(G18) );
  XOR2_X1 U764 ( .A(G125), .B(KEYINPUT37), .Z(n696) );
  XNOR2_X1 U765 ( .A(n697), .B(n696), .ZN(G27) );
  INV_X1 U766 ( .A(n698), .ZN(n699) );
  XOR2_X1 U767 ( .A(G134), .B(n699), .Z(n700) );
  XNOR2_X1 U768 ( .A(KEYINPUT116), .B(n700), .ZN(G36) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n357), .A2(n705), .ZN(n706) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n710) );
  BUF_X1 U773 ( .A(n708), .Z(n709) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n727) );
  NOR2_X1 U775 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U776 ( .A(n713), .B(KEYINPUT49), .ZN(n714) );
  NAND2_X1 U777 ( .A1(n715), .A2(n714), .ZN(n719) );
  XNOR2_X1 U778 ( .A(n717), .B(KEYINPUT50), .ZN(n718) );
  NOR2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U780 ( .A(KEYINPUT117), .B(n720), .Z(n721) );
  NOR2_X1 U781 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U782 ( .A(KEYINPUT51), .B(n723), .ZN(n725) );
  INV_X1 U783 ( .A(n724), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n725), .A2(n732), .ZN(n726) );
  NAND2_X1 U785 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U786 ( .A(n728), .B(KEYINPUT52), .ZN(n729) );
  XOR2_X1 U787 ( .A(KEYINPUT118), .B(n729), .Z(n730) );
  NOR2_X1 U788 ( .A1(n731), .A2(n730), .ZN(n735) );
  AND2_X1 U789 ( .A1(n709), .A2(n732), .ZN(n733) );
  XOR2_X1 U790 ( .A(KEYINPUT119), .B(n733), .Z(n734) );
  NOR2_X1 U791 ( .A1(n735), .A2(n734), .ZN(n745) );
  NOR2_X1 U792 ( .A1(n736), .A2(KEYINPUT87), .ZN(n737) );
  XNOR2_X1 U793 ( .A(n737), .B(KEYINPUT2), .ZN(n743) );
  INV_X1 U794 ( .A(n738), .ZN(n740) );
  NAND2_X1 U795 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U796 ( .A1(n741), .A2(KEYINPUT87), .ZN(n742) );
  NAND2_X1 U797 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U798 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n746), .A2(G953), .ZN(n747) );
  XNOR2_X1 U800 ( .A(n747), .B(KEYINPUT53), .ZN(G75) );
  BUF_X1 U801 ( .A(n748), .Z(n749) );
  NAND2_X1 U802 ( .A1(n749), .A2(G478), .ZN(n751) );
  XNOR2_X1 U803 ( .A(n751), .B(n750), .ZN(n752) );
  NOR2_X1 U804 ( .A1(n753), .A2(n752), .ZN(G63) );
  XOR2_X1 U805 ( .A(KEYINPUT126), .B(n754), .Z(n756) );
  NOR2_X1 U806 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U807 ( .A(KEYINPUT125), .B(n757), .Z(n765) );
  NOR2_X1 U808 ( .A1(n738), .A2(G953), .ZN(n758) );
  XOR2_X1 U809 ( .A(KEYINPUT124), .B(n758), .Z(n763) );
  XOR2_X1 U810 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n760) );
  NAND2_X1 U811 ( .A1(G224), .A2(G953), .ZN(n759) );
  XNOR2_X1 U812 ( .A(n760), .B(n759), .ZN(n761) );
  NAND2_X1 U813 ( .A1(n761), .A2(G898), .ZN(n762) );
  NAND2_X1 U814 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U815 ( .A(n765), .B(n764), .ZN(G69) );
  XOR2_X1 U816 ( .A(n767), .B(n766), .Z(n771) );
  INV_X1 U817 ( .A(n771), .ZN(n768) );
  XNOR2_X1 U818 ( .A(n768), .B(n375), .ZN(n770) );
  NAND2_X1 U819 ( .A1(n770), .A2(n769), .ZN(n775) );
  XNOR2_X1 U820 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U821 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U822 ( .A1(n773), .A2(G953), .ZN(n774) );
  NAND2_X1 U823 ( .A1(n775), .A2(n774), .ZN(G72) );
  XOR2_X1 U824 ( .A(G137), .B(n776), .Z(G39) );
  XNOR2_X1 U825 ( .A(G140), .B(n777), .ZN(G42) );
  XOR2_X1 U826 ( .A(G131), .B(n778), .Z(G33) );
  XNOR2_X1 U827 ( .A(G143), .B(n779), .ZN(G45) );
endmodule

