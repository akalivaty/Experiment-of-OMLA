//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  OAI211_X1 g009(.A(G128), .B(new_n192), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n197), .B(new_n198), .C1(KEYINPUT1), .C2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G137), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n203), .A2(G137), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n203), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .A4(new_n204), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n207), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n196), .A2(new_n215), .A3(new_n200), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n202), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n209), .A2(new_n204), .A3(new_n211), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n213), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n197), .A2(new_n198), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n217), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT68), .B1(new_n217), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n190), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT28), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n217), .A2(new_n228), .ZN(new_n234));
  INV_X1    g048(.A(new_n190), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n217), .A2(new_n190), .A3(new_n228), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT28), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G237), .ZN(new_n242));
  INV_X1    g056(.A(G953), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(G210), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n244), .B(KEYINPUT27), .Z(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(G902), .B1(new_n241), .B2(new_n249), .ZN(new_n250));
  AND4_X1   g064(.A1(new_n207), .A2(new_n196), .A3(new_n213), .A4(new_n200), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n222), .B(new_n253), .C1(new_n225), .C2(new_n226), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n252), .A2(new_n254), .B1(new_n213), .B2(new_n219), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n258));
  INV_X1    g072(.A(new_n254), .ZN(new_n259));
  OAI22_X1  g073(.A1(new_n193), .A2(new_n195), .B1(new_n224), .B2(new_n223), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n260), .B2(new_n222), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n220), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n257), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n258), .B1(new_n217), .B2(new_n228), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n190), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n237), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n247), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n190), .B1(new_n257), .B2(new_n263), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT28), .B1(new_n270), .B2(new_n268), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n233), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n269), .B(new_n248), .C1(new_n272), .C2(new_n247), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n250), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n187), .B1(new_n274), .B2(G472), .ZN(new_n275));
  INV_X1    g089(.A(G472), .ZN(new_n276));
  AOI211_X1 g090(.A(KEYINPUT69), .B(new_n276), .C1(new_n250), .C2(new_n273), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n256), .B(new_n220), .C1(new_n259), .C2(new_n261), .ZN(new_n279));
  INV_X1    g093(.A(new_n251), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n252), .A2(new_n254), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n256), .B1(new_n282), .B2(new_n220), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n281), .A2(new_n283), .A3(KEYINPUT30), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n235), .B1(new_n284), .B2(new_n265), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  INV_X1    g100(.A(new_n247), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .A4(new_n237), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT67), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n264), .A2(new_n266), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n268), .B1(new_n291), .B2(new_n235), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n292), .A2(KEYINPUT67), .A3(new_n286), .A4(new_n287), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n285), .A2(new_n287), .A3(new_n237), .ZN(new_n295));
  AOI22_X1  g109(.A1(KEYINPUT31), .A2(new_n295), .B1(new_n272), .B2(new_n247), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n276), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n298), .B1(new_n297), .B2(new_n276), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n278), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G119), .ZN(new_n303));
  OR3_X1    g117(.A1(new_n303), .A2(KEYINPUT23), .A3(G128), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT23), .B1(new_n303), .B2(G128), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n199), .A2(G119), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G110), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n199), .A2(KEYINPUT72), .A3(G119), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT72), .B1(new_n199), .B2(G119), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n310), .A2(new_n311), .B1(G119), .B2(new_n199), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT24), .B(G110), .Z(new_n313));
  OAI21_X1  g127(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n319), .A2(KEYINPUT16), .A3(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(G146), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(new_n315), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n194), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n316), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n320), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(G146), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n312), .A2(new_n313), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n308), .B2(new_n307), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n243), .A2(G221), .A3(G234), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT74), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G137), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n334), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n324), .A2(new_n329), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G217), .ZN(new_n339));
  INV_X1    g153(.A(G902), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(G234), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n341), .B(KEYINPUT70), .Z(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n340), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n342), .B(KEYINPUT71), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n338), .A2(G902), .ZN(new_n346));
  NOR2_X1   g160(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n338), .A2(G902), .B1(KEYINPUT75), .B2(KEYINPUT25), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G110), .B(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n243), .A2(G227), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g171(.A(G104), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G107), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  INV_X1    g176(.A(G107), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT76), .A4(G104), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n358), .A2(G107), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n361), .A2(new_n366), .A3(KEYINPUT77), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n363), .A2(G104), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n359), .B2(new_n357), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n362), .A2(KEYINPUT76), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n362), .A2(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n363), .A2(G104), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n368), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(G101), .B(new_n355), .C1(new_n367), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G101), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT77), .B1(new_n361), .B2(new_n366), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n370), .A2(new_n368), .A3(new_n374), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n370), .A2(new_n377), .A3(new_n374), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n376), .B(new_n227), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n220), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n196), .A2(new_n215), .A3(new_n200), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n215), .B1(new_n196), .B2(new_n200), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G101), .B1(new_n359), .B2(new_n369), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n381), .A2(KEYINPUT10), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n381), .A2(new_n200), .A3(new_n196), .A4(new_n388), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n391));
  AOI22_X1  g205(.A1(new_n387), .A2(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n383), .A2(new_n384), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n384), .B1(new_n383), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n354), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(KEYINPUT81), .A3(new_n353), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n381), .A2(new_n388), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n201), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n384), .B1(new_n399), .B2(new_n390), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(KEYINPUT12), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT81), .B1(new_n393), .B2(new_n353), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n396), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G469), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n340), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n394), .A2(new_n395), .A3(new_n354), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n353), .B1(new_n401), .B2(new_n393), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n340), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n408), .B1(new_n411), .B2(G469), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n408), .A3(G469), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n191), .A2(G128), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n199), .A2(G143), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n203), .ZN(new_n419));
  INV_X1    g233(.A(G116), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G122), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(G122), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(KEYINPUT14), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(KEYINPUT14), .B2(new_n421), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G107), .ZN(new_n425));
  XNOR2_X1  g239(.A(G116), .B(G122), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n363), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n416), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(KEYINPUT13), .B2(new_n417), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n429), .A2(KEYINPUT13), .ZN(new_n431));
  OAI21_X1  g245(.A(G134), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n418), .A2(new_n203), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n426), .B(new_n363), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT9), .B(G234), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n437), .A2(new_n339), .A3(G953), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT90), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(new_n441), .A3(new_n438), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n436), .A2(new_n438), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n340), .ZN(new_n445));
  INV_X1    g259(.A(G478), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n445), .B(new_n451), .Z(new_n452));
  NAND2_X1  g266(.A1(new_n243), .A2(G952), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(G234), .B2(G237), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n340), .B(new_n243), .C1(G234), .C2(G237), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(G898), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n242), .A2(new_n243), .A3(G214), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(G143), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT89), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n460), .A2(new_n212), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n317), .A2(new_n194), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n464), .A2(KEYINPUT18), .B1(new_n323), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G113), .B(G122), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n358), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(KEYINPUT17), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n460), .B(new_n212), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n326), .B(new_n470), .C1(new_n471), .C2(KEYINPUT17), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n317), .B(KEYINPUT19), .Z(new_n474));
  MUX2_X1   g288(.A(new_n325), .B(new_n474), .S(new_n194), .Z(new_n475));
  AOI22_X1  g289(.A1(new_n463), .A2(new_n466), .B1(new_n475), .B2(new_n471), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n476), .B2(new_n469), .ZN(new_n477));
  NOR2_X1   g291(.A1(G475), .A2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT20), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n473), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n469), .B1(new_n467), .B2(new_n472), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n340), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G475), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n452), .A2(new_n458), .A3(new_n483), .A4(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n437), .B2(G902), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n415), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G214), .B1(G237), .B2(G902), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT82), .Z(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n227), .A2(G125), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(G125), .B2(new_n201), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT86), .Z(new_n498));
  INV_X1    g312(.A(G224), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(G953), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n498), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(G110), .B(G122), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n398), .ZN(new_n504));
  INV_X1    g318(.A(new_n188), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(new_n189), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n188), .A2(KEYINPUT5), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n420), .A2(KEYINPUT5), .A3(G119), .ZN(new_n508));
  INV_X1    g322(.A(G113), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n506), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n376), .B(new_n235), .C1(new_n380), .C2(new_n382), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(KEYINPUT83), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT83), .ZN(new_n515));
  OAI21_X1  g329(.A(G101), .B1(new_n367), .B2(new_n375), .ZN(new_n516));
  INV_X1    g330(.A(new_n382), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n190), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n515), .B1(new_n518), .B2(new_n376), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT85), .B(new_n503), .C1(new_n514), .C2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n515), .A3(new_n376), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n512), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n525), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n503), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT84), .B1(new_n525), .B2(new_n503), .ZN(new_n528));
  INV_X1    g342(.A(new_n514), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT84), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n523), .A4(new_n502), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(new_n503), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n501), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n528), .A2(new_n531), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT7), .B1(new_n499), .B2(G953), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n497), .B(new_n536), .Z(new_n537));
  NOR2_X1   g351(.A1(new_n504), .A2(new_n511), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT87), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n510), .B1(new_n507), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n539), .B2(new_n507), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n541), .A2(new_n506), .A3(new_n398), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n538), .B1(new_n542), .B2(KEYINPUT88), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(KEYINPUT88), .B2(new_n542), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n502), .B(KEYINPUT8), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n537), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n340), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n495), .B1(new_n534), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n501), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n522), .A2(new_n526), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n535), .B2(new_n546), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n494), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n493), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n302), .A2(new_n350), .A3(new_n491), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT92), .B(G101), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(G3));
  INV_X1    g373(.A(new_n493), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n534), .A2(new_n548), .A3(new_n495), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n494), .B1(new_n553), .B2(new_n554), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n560), .B(new_n458), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n482), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n481), .B1(new_n477), .B2(new_n478), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n487), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n445), .A2(new_n446), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n444), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n443), .A2(KEYINPUT33), .A3(new_n439), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n446), .A2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n568), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n567), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n563), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n294), .A2(new_n296), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n340), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n297), .A2(new_n276), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n411), .A2(new_n408), .A3(G469), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n406), .B1(new_n585), .B2(new_n412), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n350), .A3(new_n489), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT93), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT34), .B(G104), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  NOR2_X1   g406(.A1(new_n452), .A2(new_n566), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n563), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n588), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G107), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT94), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(G9));
  INV_X1    g413(.A(new_n584), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n330), .A2(KEYINPUT36), .A3(new_n334), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n334), .A2(KEYINPUT36), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n324), .B2(new_n329), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n601), .A2(new_n343), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n348), .B2(new_n349), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n600), .A2(new_n491), .A3(new_n556), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT95), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT37), .B(G110), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G12));
  XNOR2_X1  g424(.A(new_n445), .B(new_n451), .ZN(new_n611));
  INV_X1    g425(.A(new_n454), .ZN(new_n612));
  INV_X1    g426(.A(new_n455), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(G900), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n611), .A2(new_n483), .A3(new_n487), .A4(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n415), .A2(new_n490), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n302), .A2(new_n556), .A3(new_n616), .A4(new_n606), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT96), .B(G128), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G30));
  XNOR2_X1  g433(.A(new_n614), .B(KEYINPUT39), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n586), .A2(new_n489), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT99), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n623), .A2(KEYINPUT40), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(KEYINPUT40), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n549), .A2(new_n555), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n566), .A2(new_n560), .A3(new_n611), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n628), .A2(new_n606), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n624), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n583), .A2(KEYINPUT32), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n299), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n238), .A2(new_n247), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n295), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n276), .B1(new_n635), .B2(new_n340), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT98), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n639), .B(new_n636), .C1(new_n632), .C2(new_n299), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n191), .ZN(G45));
  NAND3_X1  g457(.A1(new_n566), .A2(new_n575), .A3(new_n614), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n415), .A2(new_n490), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n302), .A2(new_n556), .A3(new_n645), .A4(new_n606), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G146), .ZN(G48));
  INV_X1    g461(.A(new_n350), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n633), .B2(new_n278), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n404), .A2(new_n340), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G469), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n489), .A3(new_n406), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n649), .A2(new_n579), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT41), .B(G113), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G15));
  NAND3_X1  g470(.A1(new_n649), .A2(new_n595), .A3(new_n653), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G116), .ZN(G18));
  AOI21_X1  g472(.A(new_n605), .B1(new_n633), .B2(new_n278), .ZN(new_n659));
  NOR4_X1   g473(.A1(new_n652), .A2(new_n457), .A3(new_n566), .A4(new_n611), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n556), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G119), .ZN(G21));
  AOI21_X1  g476(.A(new_n276), .B1(new_n580), .B2(new_n340), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n276), .A2(new_n340), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n295), .A2(KEYINPUT31), .B1(new_n240), .B2(new_n247), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n664), .B1(new_n294), .B2(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n663), .A2(new_n648), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n629), .B1(new_n549), .B2(new_n555), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n667), .A2(new_n458), .A3(new_n653), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G122), .ZN(G24));
  AOI211_X1 g484(.A(new_n493), .B(new_n652), .C1(new_n549), .C2(new_n555), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n644), .B(KEYINPUT101), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n666), .B1(new_n581), .B2(G472), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT100), .B1(new_n673), .B2(new_n606), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n663), .A2(new_n605), .A3(new_n675), .A4(new_n666), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n671), .B(new_n672), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G125), .ZN(G27));
  NAND4_X1  g492(.A1(new_n549), .A2(new_n560), .A3(new_n555), .A4(new_n489), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n407), .B1(G469), .B2(new_n411), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n649), .A2(new_n672), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n649), .A2(KEYINPUT42), .A3(new_n672), .A4(new_n681), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G131), .ZN(G33));
  INV_X1    g501(.A(new_n615), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n681), .A2(new_n350), .A3(new_n302), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G134), .ZN(G36));
  NAND4_X1  g504(.A1(new_n575), .A2(new_n483), .A3(KEYINPUT43), .A4(new_n487), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n576), .B2(new_n566), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n692), .B(new_n694), .C1(new_n576), .C2(new_n566), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n584), .A3(new_n606), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n401), .A2(new_n393), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n354), .ZN(new_n705));
  INV_X1    g519(.A(new_n395), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n353), .A3(new_n393), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n705), .A2(KEYINPUT45), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT102), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT45), .B1(new_n705), .B2(new_n707), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n405), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n405), .A2(new_n340), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(KEYINPUT46), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n406), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT46), .B1(new_n712), .B2(new_n714), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n490), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n626), .A2(new_n493), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n699), .B2(new_n700), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n703), .A2(new_n620), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G137), .ZN(G39));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n725), .B(new_n726), .C1(new_n718), .C2(new_n490), .ZN(new_n727));
  INV_X1    g541(.A(new_n717), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n406), .A3(new_n715), .ZN(new_n729));
  NAND2_X1  g543(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n725), .A2(new_n726), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n729), .A2(new_n489), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n721), .A2(new_n302), .A3(new_n350), .A4(new_n644), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  NOR2_X1   g550(.A1(new_n652), .A2(new_n560), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n628), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT111), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n628), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n612), .B1(new_n696), .B2(new_n697), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n667), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT50), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n747), .B(new_n744), .C1(new_n739), .C2(new_n741), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n651), .A2(new_n406), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n727), .B(new_n732), .C1(new_n489), .C2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n745), .A2(new_n753), .A3(new_n720), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT110), .B1(new_n744), .B2(new_n721), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n673), .A2(new_n606), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n675), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n673), .A2(KEYINPUT100), .A3(new_n606), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n679), .A2(new_n751), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n743), .A2(new_n762), .A3(KEYINPUT112), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT112), .B1(new_n743), .B2(new_n762), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n350), .A2(new_n454), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n566), .A2(new_n575), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n641), .A2(new_n762), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n757), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT51), .B1(new_n750), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n757), .A2(new_n765), .A3(new_n769), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n749), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n453), .B1(new_n745), .B2(new_n671), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n641), .A2(new_n577), .A3(new_n762), .A4(new_n767), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n649), .B1(new_n763), .B2(new_n764), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT48), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n781), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(KEYINPUT48), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n779), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n771), .A2(new_n774), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n654), .A2(new_n657), .A3(new_n661), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n493), .B(new_n457), .C1(new_n549), .C2(new_n555), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n588), .B(new_n790), .C1(new_n577), .C2(new_n593), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n557), .A3(new_n669), .A4(new_n607), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n761), .A2(new_n672), .A3(new_n681), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT107), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT107), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n761), .A2(new_n796), .A3(new_n672), .A4(new_n681), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n452), .A2(new_n487), .A3(new_n483), .A4(new_n614), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n415), .A2(new_n799), .A3(new_n490), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n302), .A2(new_n720), .A3(new_n606), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n689), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n684), .B2(new_n685), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n793), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n677), .A2(new_n617), .A3(new_n646), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n605), .A2(new_n489), .A3(new_n614), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n680), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n668), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n637), .B1(new_n300), .B2(new_n301), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n639), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n633), .A2(KEYINPUT98), .A3(new_n637), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT108), .B1(new_n805), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n659), .B(new_n556), .C1(new_n616), .C2(new_n645), .ZN(new_n814));
  INV_X1    g628(.A(new_n808), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n638), .B2(new_n640), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT108), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n814), .A2(new_n816), .A3(new_n817), .A4(new_n677), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n813), .A2(KEYINPUT52), .A3(new_n818), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  INV_X1    g640(.A(new_n805), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n816), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n804), .A2(new_n819), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(new_n824), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n793), .A2(new_n798), .A3(new_n803), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n813), .A2(new_n818), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n826), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n834), .A3(KEYINPUT53), .A4(new_n821), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT109), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n820), .A2(new_n837), .A3(KEYINPUT53), .A4(new_n821), .ZN(new_n838));
  INV_X1    g652(.A(new_n828), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n820), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n836), .A2(new_n838), .B1(new_n825), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n788), .B(new_n831), .C1(new_n841), .C2(new_n824), .ZN(new_n842));
  NOR2_X1   g656(.A1(G952), .A2(G953), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT115), .Z(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n751), .B(KEYINPUT49), .Z(new_n846));
  NAND2_X1  g660(.A1(new_n560), .A2(new_n489), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n648), .A2(new_n566), .A3(new_n576), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n641), .A2(new_n628), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n845), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(G75));
  NOR2_X1   g668(.A1(new_n243), .A2(G952), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(G902), .B1(new_n822), .B2(new_n829), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT56), .B1(new_n858), .B2(G210), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n551), .A2(new_n552), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(new_n550), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT55), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n856), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(KEYINPUT117), .B(G902), .C1(new_n822), .C2(new_n829), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n495), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT118), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(KEYINPUT118), .B2(new_n862), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n863), .B1(new_n867), .B2(new_n870), .ZN(G51));
  INV_X1    g685(.A(new_n712), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n865), .A2(new_n872), .A3(new_n866), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT120), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n865), .A2(new_n875), .A3(new_n872), .A4(new_n866), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n822), .A2(new_n829), .A3(KEYINPUT119), .A4(KEYINPUT54), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n822), .B2(new_n829), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n831), .B2(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n713), .B(KEYINPUT57), .Z(new_n883));
  OAI21_X1  g697(.A(new_n404), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n855), .B1(new_n877), .B2(new_n884), .ZN(G54));
  NAND4_X1  g699(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .A4(new_n866), .ZN(new_n886));
  INV_X1    g700(.A(new_n477), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(new_n855), .ZN(G60));
  INV_X1    g704(.A(new_n572), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n446), .A2(new_n340), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n856), .B1(new_n882), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n831), .B1(new_n841), .B2(new_n824), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n891), .B1(new_n897), .B2(new_n894), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(G63));
  NAND2_X1  g713(.A1(new_n823), .A2(new_n830), .ZN(new_n900));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT60), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n338), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n601), .A2(new_n603), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n900), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n856), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(G66));
  INV_X1    g723(.A(new_n793), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(KEYINPUT122), .A3(new_n243), .ZN(new_n911));
  OAI21_X1  g725(.A(G953), .B1(new_n456), .B2(new_n499), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT122), .B1(new_n910), .B2(new_n243), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n860), .B1(G898), .B2(new_n243), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n915), .B(new_n916), .Z(G69));
  XNOR2_X1  g731(.A(new_n474), .B(KEYINPUT123), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n291), .B(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n719), .A2(new_n649), .A3(new_n620), .A4(new_n668), .ZN(new_n920));
  AND4_X1   g734(.A1(new_n689), .A2(new_n723), .A3(new_n735), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n805), .B1(new_n684), .B2(new_n685), .ZN(new_n922));
  AOI21_X1  g736(.A(G953), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n243), .A2(G900), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT125), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n919), .B(KEYINPUT124), .Z(new_n927));
  AOI21_X1  g741(.A(new_n621), .B1(new_n578), .B2(new_n594), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n649), .A2(new_n720), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n723), .A2(new_n735), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n642), .B2(new_n805), .ZN(new_n932));
  OAI211_X1 g746(.A(KEYINPUT62), .B(new_n827), .C1(new_n631), .C2(new_n641), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n934), .B2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n243), .B1(G227), .B2(G900), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G72));
  NAND3_X1  g752(.A1(new_n921), .A2(new_n793), .A3(new_n922), .ZN(new_n939));
  NAND2_X1  g753(.A1(G472), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT63), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n267), .A2(new_n287), .A3(new_n268), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n855), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n941), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n934), .B2(new_n793), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n292), .A2(new_n247), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n946), .B2(new_n947), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n944), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n841), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n945), .B1(new_n269), .B2(new_n295), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT127), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(G57));
endmodule


