

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  NOR2_X2 U326 ( .A1(n544), .A2(n490), .ZN(n571) );
  XNOR2_X1 U327 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U328 ( .A(KEYINPUT73), .B(n564), .ZN(n570) );
  XOR2_X1 U329 ( .A(n487), .B(KEYINPUT28), .Z(n536) );
  XOR2_X1 U330 ( .A(n460), .B(KEYINPUT107), .Z(n294) );
  XOR2_X1 U331 ( .A(n443), .B(n361), .Z(n295) );
  XOR2_X1 U332 ( .A(n359), .B(n358), .Z(n296) );
  XNOR2_X1 U333 ( .A(n483), .B(KEYINPUT54), .ZN(n484) );
  XNOR2_X1 U334 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U335 ( .A(n326), .B(n325), .ZN(n331) );
  XNOR2_X1 U336 ( .A(n360), .B(n296), .ZN(n364) );
  XNOR2_X1 U337 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n488) );
  NOR2_X1 U338 ( .A1(n465), .A2(n425), .ZN(n426) );
  XNOR2_X1 U339 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U340 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U341 ( .A(n334), .B(n333), .Z(n564) );
  XOR2_X1 U342 ( .A(n383), .B(n382), .Z(n534) );
  INV_X1 U343 ( .A(G29GAT), .ZN(n461) );
  XNOR2_X1 U344 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U345 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U346 ( .A(n495), .B(n494), .ZN(G1349GAT) );
  XNOR2_X1 U347 ( .A(n464), .B(n463), .ZN(G1328GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT6), .B(G57GAT), .Z(n298) );
  XNOR2_X1 U349 ( .A(KEYINPUT1), .B(KEYINPUT93), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n318) );
  XOR2_X1 U351 ( .A(KEYINPUT5), .B(G127GAT), .Z(n300) );
  XNOR2_X1 U352 ( .A(G1GAT), .B(G120GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U354 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n302) );
  XNOR2_X1 U355 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U357 ( .A(n304), .B(n303), .Z(n316) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n305), .B(KEYINPUT2), .ZN(n358) );
  XOR2_X1 U360 ( .A(n358), .B(KEYINPUT89), .Z(n307) );
  NAND2_X1 U361 ( .A1(G225GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n314) );
  XOR2_X1 U363 ( .A(G155GAT), .B(G148GAT), .Z(n309) );
  XNOR2_X1 U364 ( .A(G134GAT), .B(G162GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U366 ( .A(n310), .B(G85GAT), .Z(n312) );
  XOR2_X1 U367 ( .A(G113GAT), .B(KEYINPUT0), .Z(n369) );
  XNOR2_X1 U368 ( .A(G29GAT), .B(n369), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n395) );
  INV_X1 U373 ( .A(n395), .ZN(n529) );
  XOR2_X1 U374 ( .A(KEYINPUT36), .B(KEYINPUT106), .Z(n335) );
  XOR2_X1 U375 ( .A(G162GAT), .B(KEYINPUT70), .Z(n320) );
  XNOR2_X1 U376 ( .A(G50GAT), .B(G218GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n359) );
  XNOR2_X1 U378 ( .A(n359), .B(KEYINPUT10), .ZN(n326) );
  XOR2_X1 U379 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n322) );
  XNOR2_X1 U380 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n324) );
  AND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U383 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n327), .B(KEYINPUT7), .ZN(n429) );
  XOR2_X1 U385 ( .A(G92GAT), .B(G85GAT), .Z(n329) );
  XNOR2_X1 U386 ( .A(G99GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n456) );
  XOR2_X1 U388 ( .A(n429), .B(n456), .Z(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(G43GAT), .B(G134GAT), .Z(n372) );
  XNOR2_X1 U391 ( .A(n332), .B(n372), .ZN(n334) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(G190GAT), .ZN(n344) );
  INV_X1 U393 ( .A(n344), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n335), .B(n570), .ZN(n465) );
  XOR2_X1 U395 ( .A(G8GAT), .B(G183GAT), .Z(n405) );
  XOR2_X1 U396 ( .A(G204GAT), .B(G64GAT), .Z(n449) );
  XOR2_X1 U397 ( .A(n405), .B(n449), .Z(n340) );
  XOR2_X1 U398 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n337) );
  XNOR2_X1 U399 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n337), .B(n336), .ZN(n368) );
  XNOR2_X1 U401 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n338), .B(G211GAT), .ZN(n361) );
  XNOR2_X1 U403 ( .A(n368), .B(n361), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n348) );
  XOR2_X1 U405 ( .A(KEYINPUT94), .B(G92GAT), .Z(n342) );
  XNOR2_X1 U406 ( .A(G176GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n346) );
  NAND2_X1 U409 ( .A1(G226GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U411 ( .A(n348), .B(n347), .Z(n532) );
  XOR2_X1 U412 ( .A(n532), .B(KEYINPUT95), .Z(n349) );
  XNOR2_X1 U413 ( .A(KEYINPUT27), .B(n349), .ZN(n389) );
  NAND2_X1 U414 ( .A1(n389), .A2(n529), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n350), .B(KEYINPUT96), .ZN(n541) );
  XOR2_X1 U416 ( .A(KEYINPUT24), .B(KEYINPUT84), .Z(n352) );
  XNOR2_X1 U417 ( .A(KEYINPUT85), .B(KEYINPUT23), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n366) );
  XOR2_X1 U419 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n354) );
  XNOR2_X1 U420 ( .A(KEYINPUT88), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U422 ( .A(n355), .B(KEYINPUT87), .Z(n357) );
  XOR2_X1 U423 ( .A(G22GAT), .B(G155GAT), .Z(n411) );
  XNOR2_X1 U424 ( .A(n411), .B(G106GAT), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n360) );
  XOR2_X1 U426 ( .A(G148GAT), .B(G78GAT), .Z(n443) );
  NAND2_X1 U427 ( .A1(G228GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n295), .B(n362), .ZN(n363) );
  XOR2_X1 U429 ( .A(n366), .B(n365), .Z(n487) );
  INV_X1 U430 ( .A(n536), .ZN(n542) );
  XNOR2_X1 U431 ( .A(G71GAT), .B(G176GAT), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n367), .B(G120GAT), .ZN(n457) );
  XNOR2_X1 U433 ( .A(n368), .B(n457), .ZN(n383) );
  XOR2_X1 U434 ( .A(G15GAT), .B(G127GAT), .Z(n412) );
  XOR2_X1 U435 ( .A(n369), .B(n412), .Z(n371) );
  NAND2_X1 U436 ( .A1(G227GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n371), .B(n370), .ZN(n373) );
  XOR2_X1 U438 ( .A(n373), .B(n372), .Z(n381) );
  XOR2_X1 U439 ( .A(KEYINPUT81), .B(G183GAT), .Z(n375) );
  XNOR2_X1 U440 ( .A(G99GAT), .B(G190GAT), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U442 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n377) );
  XNOR2_X1 U443 ( .A(KEYINPUT82), .B(KEYINPUT79), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n382) );
  INV_X1 U447 ( .A(n534), .ZN(n544) );
  XOR2_X1 U448 ( .A(KEYINPUT83), .B(n544), .Z(n384) );
  NAND2_X1 U449 ( .A1(n542), .A2(n384), .ZN(n385) );
  NOR2_X1 U450 ( .A1(n541), .A2(n385), .ZN(n386) );
  XNOR2_X1 U451 ( .A(KEYINPUT97), .B(n386), .ZN(n398) );
  NOR2_X1 U452 ( .A1(n487), .A2(n534), .ZN(n388) );
  XNOR2_X1 U453 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n576) );
  NAND2_X1 U455 ( .A1(n389), .A2(n576), .ZN(n394) );
  NAND2_X1 U456 ( .A1(n532), .A2(n534), .ZN(n390) );
  XOR2_X1 U457 ( .A(KEYINPUT99), .B(n390), .Z(n391) );
  NAND2_X1 U458 ( .A1(n487), .A2(n391), .ZN(n392) );
  XOR2_X1 U459 ( .A(KEYINPUT25), .B(n392), .Z(n393) );
  NAND2_X1 U460 ( .A1(n394), .A2(n393), .ZN(n396) );
  NAND2_X1 U461 ( .A1(n396), .A2(n395), .ZN(n397) );
  NAND2_X1 U462 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n399), .B(KEYINPUT100), .ZN(n500) );
  XOR2_X1 U464 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n401) );
  XNOR2_X1 U465 ( .A(KEYINPUT15), .B(KEYINPUT77), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n402), .B(KEYINPUT75), .ZN(n424) );
  XOR2_X1 U468 ( .A(KEYINPUT14), .B(G64GAT), .Z(n404) );
  XNOR2_X1 U469 ( .A(G78GAT), .B(G211GAT), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U472 ( .A(G1GAT), .B(G71GAT), .Z(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U474 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n409), .B(KEYINPUT66), .ZN(n444) );
  XNOR2_X1 U476 ( .A(n410), .B(n444), .ZN(n413) );
  XOR2_X1 U477 ( .A(n412), .B(n411), .Z(n414) );
  NAND2_X1 U478 ( .A1(n413), .A2(n414), .ZN(n418) );
  INV_X1 U479 ( .A(n413), .ZN(n416) );
  INV_X1 U480 ( .A(n414), .ZN(n415) );
  NAND2_X1 U481 ( .A1(n416), .A2(n415), .ZN(n417) );
  NAND2_X1 U482 ( .A1(n418), .A2(n417), .ZN(n422) );
  XOR2_X1 U483 ( .A(KEYINPUT74), .B(KEYINPUT78), .Z(n420) );
  NAND2_X1 U484 ( .A1(G231GAT), .A2(G233GAT), .ZN(n419) );
  XOR2_X1 U485 ( .A(n420), .B(n419), .Z(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U487 ( .A(n424), .B(n423), .Z(n473) );
  NAND2_X1 U488 ( .A1(n500), .A2(n473), .ZN(n425) );
  XNOR2_X1 U489 ( .A(KEYINPUT37), .B(n426), .ZN(n528) );
  XOR2_X1 U490 ( .A(G197GAT), .B(G141GAT), .Z(n428) );
  XNOR2_X1 U491 ( .A(G36GAT), .B(G22GAT), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n442) );
  XOR2_X1 U493 ( .A(G43GAT), .B(n429), .Z(n431) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U496 ( .A(n432), .B(G50GAT), .Z(n440) );
  XOR2_X1 U497 ( .A(G1GAT), .B(G15GAT), .Z(n434) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(G113GAT), .ZN(n433) );
  XNOR2_X1 U499 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U500 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n436) );
  XNOR2_X1 U501 ( .A(G8GAT), .B(KEYINPUT65), .ZN(n435) );
  XNOR2_X1 U502 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n578) );
  INV_X1 U506 ( .A(n578), .ZN(n566) );
  XNOR2_X1 U507 ( .A(n444), .B(n443), .ZN(n446) );
  AND2_X1 U508 ( .A1(G230GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n446), .B(n445), .ZN(n448) );
  INV_X1 U510 ( .A(KEYINPUT67), .ZN(n447) );
  XNOR2_X1 U511 ( .A(n448), .B(n447), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n449), .B(KEYINPUT68), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n451), .B(n450), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n453) );
  XNOR2_X1 U515 ( .A(KEYINPUT33), .B(KEYINPUT69), .ZN(n452) );
  XNOR2_X1 U516 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U517 ( .A(n455), .B(n454), .ZN(n459) );
  XOR2_X1 U518 ( .A(n457), .B(n456), .Z(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n470) );
  NAND2_X1 U520 ( .A1(n566), .A2(n470), .ZN(n502) );
  NOR2_X1 U521 ( .A1(n528), .A2(n502), .ZN(n460) );
  XNOR2_X1 U522 ( .A(KEYINPUT38), .B(n294), .ZN(n516) );
  NAND2_X1 U523 ( .A1(n529), .A2(n516), .ZN(n464) );
  XOR2_X1 U524 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n462) );
  NOR2_X1 U525 ( .A1(n465), .A2(n473), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT45), .ZN(n468) );
  AND2_X1 U527 ( .A1(n470), .A2(n578), .ZN(n467) );
  AND2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n480) );
  XOR2_X1 U529 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n472) );
  XNOR2_X1 U530 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(n491) );
  AND2_X1 U532 ( .A1(n566), .A2(n491), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n472), .B(n471), .ZN(n474) );
  XOR2_X1 U534 ( .A(n473), .B(KEYINPUT112), .Z(n568) );
  NOR2_X1 U535 ( .A1(n474), .A2(n568), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n475), .A2(n564), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(KEYINPUT47), .ZN(n479) );
  NOR2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT48), .ZN(n540) );
  INV_X1 U542 ( .A(n540), .ZN(n482) );
  NAND2_X1 U543 ( .A1(n482), .A2(n532), .ZN(n485) );
  XOR2_X1 U544 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n483) );
  NOR2_X1 U545 ( .A1(n529), .A2(n486), .ZN(n575) );
  NAND2_X1 U546 ( .A1(n575), .A2(n487), .ZN(n489) );
  NAND2_X1 U547 ( .A1(n571), .A2(n491), .ZN(n495) );
  XOR2_X1 U548 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n493) );
  XNOR2_X1 U549 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n492) );
  XOR2_X1 U550 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n497) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n496) );
  XNOR2_X1 U552 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U553 ( .A(KEYINPUT101), .B(n498), .Z(n504) );
  NOR2_X1 U554 ( .A1(n570), .A2(n473), .ZN(n499) );
  XNOR2_X1 U555 ( .A(KEYINPUT16), .B(n499), .ZN(n501) );
  NAND2_X1 U556 ( .A1(n501), .A2(n500), .ZN(n518) );
  NOR2_X1 U557 ( .A1(n502), .A2(n518), .ZN(n509) );
  NAND2_X1 U558 ( .A1(n509), .A2(n529), .ZN(n503) );
  XNOR2_X1 U559 ( .A(n504), .B(n503), .ZN(G1324GAT) );
  NAND2_X1 U560 ( .A1(n509), .A2(n532), .ZN(n505) );
  XNOR2_X1 U561 ( .A(n505), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n507) );
  NAND2_X1 U563 ( .A1(n509), .A2(n534), .ZN(n506) );
  XNOR2_X1 U564 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(n508), .ZN(G1326GAT) );
  NAND2_X1 U566 ( .A1(n509), .A2(n536), .ZN(n510) );
  XNOR2_X1 U567 ( .A(n510), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U568 ( .A1(n516), .A2(n532), .ZN(n511) );
  XNOR2_X1 U569 ( .A(n511), .B(KEYINPUT108), .ZN(n512) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n512), .ZN(G1329GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n514) );
  NAND2_X1 U572 ( .A1(n516), .A2(n534), .ZN(n513) );
  XNOR2_X1 U573 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n515), .ZN(G1330GAT) );
  NAND2_X1 U575 ( .A1(n536), .A2(n516), .ZN(n517) );
  XNOR2_X1 U576 ( .A(G50GAT), .B(n517), .ZN(G1331GAT) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n491), .A2(n578), .ZN(n527) );
  NOR2_X1 U579 ( .A1(n527), .A2(n518), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n529), .A2(n523), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n520), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U582 ( .A1(n523), .A2(n532), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n521), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n534), .A2(n523), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U587 ( .A1(n523), .A2(n536), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(n526), .ZN(G1335GAT) );
  XOR2_X1 U590 ( .A(G85GAT), .B(KEYINPUT111), .Z(n531) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n537), .A2(n529), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n531), .B(n530), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n537), .A2(n532), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n533), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n534), .A2(n537), .ZN(n535) );
  XNOR2_X1 U597 ( .A(n535), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U599 ( .A(n538), .B(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n546) );
  NOR2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n555) );
  NAND2_X1 U603 ( .A1(n555), .A2(n542), .ZN(n543) );
  NOR2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n566), .A2(n552), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n546), .B(n545), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U608 ( .A1(n552), .A2(n491), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n549), .Z(G1341GAT) );
  NAND2_X1 U611 ( .A1(n568), .A2(n552), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n550), .B(KEYINPUT50), .ZN(n551) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U615 ( .A1(n552), .A2(n570), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n554), .B(n553), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n576), .A2(n555), .ZN(n563) );
  NOR2_X1 U618 ( .A1(n578), .A2(n563), .ZN(n556) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n556), .Z(G1344GAT) );
  INV_X1 U620 ( .A(n491), .ZN(n557) );
  NOR2_X1 U621 ( .A1(n557), .A2(n563), .ZN(n559) );
  XNOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n473), .A2(n563), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT118), .B(n561), .Z(n562) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n562), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n571), .A2(n566), .ZN(n567) );
  XNOR2_X1 U631 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n571), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n572) );
  XNOR2_X1 U636 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n574), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT124), .B(n577), .ZN(n587) );
  OR2_X1 U641 ( .A1(n578), .A2(n587), .ZN(n579) );
  XNOR2_X1 U642 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n583) );
  OR2_X1 U645 ( .A1(n587), .A2(n470), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U647 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  OR2_X1 U648 ( .A1(n587), .A2(n473), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT126), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n465), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

