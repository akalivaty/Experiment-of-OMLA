//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n461), .A2(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n454), .A2(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(KEYINPUT68), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n470), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n468), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT69), .B1(new_n470), .B2(KEYINPUT3), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(G137), .A3(new_n467), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n470), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(G160));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(new_n468), .A3(G2104), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n479), .A2(new_n485), .A3(new_n467), .A4(new_n471), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(G112), .B2(new_n467), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT70), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n479), .A2(new_n485), .A3(G2105), .A4(new_n471), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n488), .B(new_n492), .C1(G124), .C2(new_n494), .ZN(G162));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(G114), .B2(new_n467), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n486), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n469), .A2(new_n471), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n504));
  OR3_X1    g079(.A1(new_n503), .A2(new_n504), .A3(G2105), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n500), .B1(new_n502), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(G543), .B1(new_n517), .B2(new_n518), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n514), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  XNOR2_X1  g100(.A(KEYINPUT71), .B(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n521), .A2(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n516), .A2(new_n515), .ZN(new_n531));
  OAI21_X1  g106(.A(G89), .B1(new_n517), .B2(new_n518), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n519), .A2(new_n536), .B1(new_n521), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(G64), .B1(new_n516), .B2(new_n515), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n513), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AND2_X1   g117(.A1(G68), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n511), .B2(G56), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n513), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n519), .A2(new_n546), .B1(new_n521), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  OAI211_X1 g129(.A(G53), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n531), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT6), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(new_n513), .ZN(new_n561));
  NAND2_X1  g136(.A1(KEYINPUT6), .A2(G651), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n509), .A2(new_n510), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n559), .A2(G651), .B1(new_n563), .B2(G91), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n556), .A2(new_n564), .A3(KEYINPUT72), .ZN(new_n565));
  AOI21_X1  g140(.A(KEYINPUT72), .B1(new_n556), .B2(new_n564), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  OR2_X1    g143(.A1(new_n530), .A2(new_n534), .ZN(G286));
  OAI21_X1  g144(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n521), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n563), .A2(G87), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  AOI21_X1  g150(.A(new_n508), .B1(new_n561), .B2(new_n562), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n563), .A2(G86), .B1(new_n576), .B2(G48), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n509), .B2(new_n510), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n582), .B(G61), .C1(new_n516), .C2(new_n515), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(G61), .B1(new_n516), .B2(new_n515), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT73), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n590), .A2(new_n584), .A3(new_n579), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(KEYINPUT74), .A3(G651), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n578), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n589), .A2(KEYINPUT73), .B1(G73), .B2(G543), .ZN(new_n596));
  AOI211_X1 g171(.A(new_n587), .B(new_n513), .C1(new_n596), .C2(new_n584), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT74), .B1(new_n591), .B2(G651), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n594), .B(new_n577), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n595), .A2(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n513), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n519), .A2(new_n604), .B1(new_n521), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n603), .A2(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G171), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT76), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n563), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n519), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n531), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n618), .A2(G651), .B1(G54), .B2(new_n576), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT77), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n619), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(KEYINPUT77), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n610), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n610), .B1(new_n626), .B2(G868), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(G299), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G297));
  OAI21_X1  g206(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n633), .B2(G860), .ZN(G148));
  OAI21_X1  g209(.A(new_n608), .B1(new_n545), .B2(new_n548), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n625), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g213(.A(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n467), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI22_X1  g216(.A1(new_n493), .A2(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n487), .B2(G135), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT78), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n651), .B(new_n653), .Z(new_n654));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n654), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT17), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT80), .Z(new_n673));
  OAI21_X1  g248(.A(new_n670), .B1(new_n671), .B2(new_n667), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  AOI22_X1  g250(.A1(new_n675), .A2(KEYINPUT79), .B1(new_n671), .B2(new_n668), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(KEYINPUT79), .B2(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n669), .A2(new_n671), .A3(new_n667), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  NAND3_X1  g254(.A1(new_n673), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT81), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n688), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(KEYINPUT20), .ZN(new_n693));
  OAI221_X1 g268(.A(new_n690), .B1(new_n688), .B2(new_n686), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n702), .A3(new_n700), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n708), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G1971), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(G23), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n574), .B2(new_n708), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G6), .B(G305), .S(G16), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT32), .B(G1981), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n711), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n717), .B2(new_n716), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n708), .A2(G24), .ZN(new_n723));
  INV_X1    g298(.A(G290), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n708), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G1986), .Z(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  OR2_X1    g303(.A1(G95), .A2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n729), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n730));
  INV_X1    g305(.A(G119), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n493), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n487), .B2(G131), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n728), .B1(new_n733), .B2(new_n727), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT35), .B(G1991), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n726), .B1(KEYINPUT82), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(KEYINPUT82), .B2(new_n737), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n721), .A2(new_n722), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n727), .A2(G33), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n487), .A2(G139), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT83), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  INV_X1    g321(.A(G127), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n503), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n749));
  NAND2_X1  g324(.A1(G103), .A2(G2104), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G2105), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n748), .A2(G2105), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n745), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n743), .B1(new_n754), .B2(new_n727), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G2072), .Z(new_n756));
  AND2_X1   g331(.A1(new_n727), .A2(G32), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G105), .B2(new_n481), .ZN(new_n762));
  INV_X1    g337(.A(G129), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n493), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n487), .B2(G141), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT85), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n757), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT27), .B(G1996), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT86), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  NAND2_X1  g346(.A1(G160), .A2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G34), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(KEYINPUT24), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(KEYINPUT24), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(KEYINPUT84), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(KEYINPUT84), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n756), .B(new_n770), .C1(new_n771), .C2(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT87), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n708), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT23), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n630), .B2(new_n708), .ZN(new_n783));
  INV_X1    g358(.A(G1956), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n727), .A2(G35), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G162), .B2(new_n727), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT29), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n785), .B1(new_n769), .B2(new_n767), .C1(new_n788), .C2(G2090), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n727), .A2(G26), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT28), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n467), .A2(G116), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n493), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n487), .B2(G140), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n792), .B1(new_n797), .B2(new_n727), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n708), .A2(G21), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G168), .B2(new_n708), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT88), .ZN(new_n803));
  INV_X1    g378(.A(G1966), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT31), .B(G11), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(G28), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n727), .B1(new_n807), .B2(G28), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n708), .A2(G19), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n549), .B2(new_n708), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n806), .B1(new_n808), .B2(new_n809), .C1(new_n811), .C2(G1341), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n771), .B2(new_n778), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n811), .A2(G1341), .B1(G29), .B2(new_n643), .ZN(new_n814));
  NOR2_X1   g389(.A1(G5), .A2(G16), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G171), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT89), .B(G1961), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n813), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  AOI211_X1 g394(.A(new_n805), .B(new_n819), .C1(new_n788), .C2(G2090), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n626), .A2(new_n708), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G4), .B2(new_n708), .ZN(new_n822));
  INV_X1    g397(.A(G1348), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  AND4_X1   g400(.A1(new_n800), .A2(new_n820), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G27), .A2(G29), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G164), .B2(G29), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT90), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(G2078), .Z(new_n830));
  NAND4_X1  g405(.A1(new_n780), .A2(new_n790), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n742), .A2(new_n831), .ZN(G311));
  OR2_X1    g407(.A1(new_n742), .A2(new_n831), .ZN(G150));
  NOR2_X1   g408(.A1(new_n625), .A2(new_n633), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n511), .A2(G67), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n513), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  INV_X1    g414(.A(G55), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n519), .A2(new_n839), .B1(new_n521), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n545), .A2(new_n548), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G56), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n531), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(G651), .B1(new_n844), .B2(new_n543), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n563), .A2(G81), .B1(new_n576), .B2(G43), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n563), .A2(G93), .B1(new_n576), .B2(G55), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n837), .B1(new_n531), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G651), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n835), .B(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  INV_X1    g430(.A(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n838), .A2(new_n841), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n856), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(G145));
  XOR2_X1   g437(.A(G160), .B(new_n643), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT85), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n754), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(KEYINPUT92), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n765), .B(new_n797), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n502), .A2(new_n505), .ZN(new_n871));
  INV_X1    g446(.A(new_n500), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT91), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n754), .A2(KEYINPUT92), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(new_n874), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n869), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT93), .ZN(new_n880));
  INV_X1    g455(.A(G118), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n879), .A2(new_n880), .B1(new_n881), .B2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n880), .B2(new_n879), .ZN(new_n883));
  INV_X1    g458(.A(G130), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n884), .B2(new_n493), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n487), .B2(G142), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n646), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(new_n733), .Z(new_n888));
  NAND3_X1  g463(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n868), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n878), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n888), .B1(new_n878), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n865), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n878), .A2(new_n890), .ZN(new_n896));
  INV_X1    g471(.A(new_n888), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n864), .A3(new_n891), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g476(.A(new_n636), .B(new_n852), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n623), .B1(new_n565), .B2(new_n566), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT72), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n905));
  INV_X1    g480(.A(G91), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n905), .A2(new_n513), .B1(new_n906), .B2(new_n519), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT9), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n555), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n904), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n556), .A2(new_n564), .A3(KEYINPUT72), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n620), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT94), .B(KEYINPUT41), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n903), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT41), .B1(new_n903), .B2(new_n912), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n902), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n903), .A2(new_n912), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(new_n902), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT95), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n577), .B1(new_n597), .B2(new_n598), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT75), .ZN(new_n923));
  AOI21_X1  g498(.A(G290), .B1(new_n923), .B2(new_n599), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(G288), .B(G303), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n599), .A3(G290), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n925), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT42), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n921), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n919), .A2(new_n920), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n921), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n608), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n859), .A2(G868), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n935), .A2(KEYINPUT96), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT96), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G295));
  INV_X1    g514(.A(KEYINPUT97), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n934), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G868), .ZN(new_n942));
  INV_X1    g517(.A(new_n936), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n935), .A2(KEYINPUT97), .A3(new_n936), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(G331));
  OAI21_X1  g521(.A(KEYINPUT98), .B1(new_n538), .B2(new_n541), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n539), .A2(new_n540), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(G651), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT98), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n576), .A2(G52), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n561), .A2(new_n562), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n511), .A2(new_n952), .A3(G90), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(G286), .A2(new_n947), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(G171), .A2(new_n950), .A3(G168), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n853), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n955), .A2(new_n842), .A3(new_n956), .A4(new_n851), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n918), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(KEYINPUT99), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT99), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n852), .A2(new_n963), .A3(new_n956), .A4(new_n955), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n962), .A2(new_n964), .B1(new_n853), .B2(new_n957), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT100), .B1(new_n916), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT41), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n565), .A2(new_n566), .A3(new_n623), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n620), .B1(new_n910), .B2(new_n911), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n903), .A2(new_n912), .A3(new_n913), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT100), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n962), .A2(new_n964), .ZN(new_n974));
  INV_X1    g549(.A(new_n958), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n972), .B(new_n973), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n961), .B1(new_n966), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n930), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n895), .B1(new_n977), .B2(new_n930), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n928), .A2(new_n929), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n958), .A2(new_n959), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n918), .A2(new_n913), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n983), .B(new_n984), .C1(KEYINPUT41), .C2(new_n918), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n958), .A2(new_n918), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(new_n974), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G37), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n988), .A2(new_n978), .ZN(new_n989));
  OAI221_X1 g564(.A(KEYINPUT44), .B1(new_n980), .B2(new_n981), .C1(new_n989), .C2(new_n979), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n966), .A2(new_n976), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n991), .A2(new_n930), .A3(new_n960), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n981), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n978), .A3(new_n979), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT101), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT101), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(KEYINPUT44), .C1(new_n993), .C2(new_n994), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT102), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT102), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(new_n990), .C1(new_n997), .C2(new_n999), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(G397));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G164), .B2(G1384), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT103), .B(G40), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n475), .A2(new_n480), .A3(new_n482), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n765), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n797), .B(G2067), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1011), .B(new_n1012), .C1(new_n766), .C2(G1996), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n733), .B(new_n736), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT104), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(G290), .B(G1986), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n503), .A2(new_n504), .A3(G2105), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n478), .A2(G138), .A3(new_n467), .A4(new_n479), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1021), .B2(KEYINPUT4), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT45), .B(new_n1019), .C1(new_n1022), .C2(new_n500), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1008), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1006), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n873), .A2(new_n1028), .A3(new_n1019), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1029), .A3(new_n1024), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT105), .B(G2090), .ZN(new_n1031));
  OAI22_X1  g606(.A1(new_n1026), .A2(G1971), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G8), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G303), .A2(G8), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1033), .B(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1384), .B1(new_n871), .B2(new_n872), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1024), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT106), .B1(new_n1043), .B2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT106), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1045), .B(new_n1037), .C1(new_n1042), .C2(new_n1024), .ZN(new_n1046));
  OAI221_X1 g621(.A(new_n1041), .B1(new_n1040), .B2(G288), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  NOR3_X1   g623(.A1(G164), .A2(new_n1008), .A3(G1384), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n1049), .B2(new_n1037), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(KEYINPUT106), .A3(G8), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1050), .A2(new_n1051), .B1(G1976), .B2(new_n574), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1047), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1054));
  INV_X1    g629(.A(G1981), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n586), .B2(new_n577), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1055), .B(new_n577), .C1(new_n597), .C2(new_n598), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT107), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n588), .A2(new_n592), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1060), .A2(KEYINPUT107), .A3(new_n1055), .A4(new_n577), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1056), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1054), .B1(new_n1062), .B2(KEYINPUT49), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1064), .B(new_n1056), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT108), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1056), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT107), .B1(new_n593), .B2(new_n1055), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1064), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT108), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1062), .A2(KEYINPUT49), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1054), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1053), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1039), .B1(new_n1075), .B2(KEYINPUT111), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1077), .B(new_n1053), .C1(new_n1066), .C2(new_n1074), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT122), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT112), .B(KEYINPUT57), .C1(new_n907), .C2(new_n909), .ZN(new_n1080));
  OR2_X1    g655(.A1(KEYINPUT112), .A2(KEYINPUT57), .ZN(new_n1081));
  NAND2_X1  g656(.A1(KEYINPUT112), .A2(KEYINPUT57), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n556), .A2(new_n564), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1030), .A2(new_n784), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1006), .A2(new_n1023), .A3(new_n1024), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT113), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1030), .A2(new_n823), .B1(new_n799), .B2(new_n1049), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(new_n623), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1086), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1030), .A2(new_n823), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1049), .A2(new_n799), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT60), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1098), .B2(new_n623), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT119), .B(new_n620), .C1(new_n1091), .C2(KEYINPUT60), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1093), .A2(KEYINPUT61), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1019), .B1(new_n1022), .B2(new_n500), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1008), .B1(new_n1106), .B2(KEYINPUT50), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1956), .B1(new_n1107), .B2(new_n1029), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1088), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1084), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT113), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1089), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1105), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT58), .B(G1341), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1025), .A2(G1996), .B1(new_n1049), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n549), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT115), .Z(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1116), .A2(new_n549), .A3(new_n1120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1110), .A2(new_n1093), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT116), .B(KEYINPUT61), .Z(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT117), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1127), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1129), .B(new_n1130), .C1(new_n1110), .C2(new_n1093), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1114), .B(new_n1125), .C1(new_n1128), .C2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1104), .B1(new_n1132), .B2(KEYINPUT118), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1110), .B2(new_n1093), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT117), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1124), .B1(new_n1090), .B2(new_n1105), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1094), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1053), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1070), .B2(new_n1064), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1072), .B1(new_n1142), .B2(new_n1073), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1063), .A2(KEYINPUT108), .A3(new_n1065), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1140), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1077), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1075), .A2(KEYINPUT111), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1039), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1025), .B2(G2078), .ZN(new_n1152));
  INV_X1    g727(.A(G1961), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1030), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1151), .A2(G2078), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1026), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1150), .B1(new_n1157), .B2(G301), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1155), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1156), .A2(G40), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1006), .A2(new_n1023), .A3(G160), .A4(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1162), .A2(KEYINPUT123), .ZN(new_n1163));
  OAI21_X1  g738(.A(G171), .B1(new_n1162), .B2(KEYINPUT123), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1158), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(G286), .A2(G8), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT51), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1107), .A2(new_n771), .A3(new_n1029), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1025), .A2(new_n804), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1037), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1030), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1174), .A2(new_n771), .B1(new_n804), .B2(new_n1025), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT121), .B1(new_n1175), .B2(new_n1037), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1166), .B(KEYINPUT120), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT51), .B1(new_n1171), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1175), .A2(new_n1166), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1157), .A2(G301), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1159), .A2(G301), .A3(new_n1161), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1150), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1165), .A2(new_n1184), .A3(new_n1187), .ZN(new_n1188));
  AND4_X1   g763(.A1(new_n1079), .A2(new_n1139), .A3(new_n1149), .A4(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1033), .B(new_n1035), .Z(new_n1190));
  NAND2_X1  g765(.A1(new_n1171), .A2(G168), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1190), .A2(new_n1075), .A3(KEYINPUT63), .A4(new_n1192), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1076), .A2(new_n1078), .A3(new_n1191), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1193), .B1(new_n1194), .B2(KEYINPUT63), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1178), .B1(new_n1175), .B2(new_n1037), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1173), .A2(new_n1176), .B1(new_n1196), .B2(KEYINPUT51), .ZN(new_n1197));
  OAI21_X1  g772(.A(KEYINPUT62), .B1(new_n1197), .B2(new_n1182), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1181), .A2(new_n1199), .A3(new_n1183), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1198), .A2(new_n1200), .A3(new_n1185), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1201), .A2(new_n1079), .A3(new_n1149), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1145), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1203));
  NOR2_X1   g778(.A1(G288), .A2(G1976), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1204), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1141), .B1(new_n1207), .B2(KEYINPUT109), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT109), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1205), .A2(new_n1209), .A3(new_n1206), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1203), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1195), .A2(new_n1202), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1018), .B1(new_n1189), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1214));
  INV_X1    g789(.A(KEYINPUT46), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1216), .B(KEYINPUT125), .Z(new_n1217));
  INV_X1    g792(.A(new_n1009), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1218), .B1(new_n765), .B2(new_n1012), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1219), .B1(new_n1215), .B2(new_n1214), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT126), .ZN(new_n1222));
  OR2_X1    g797(.A1(new_n1222), .A2(KEYINPUT47), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(KEYINPUT47), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n733), .A2(new_n735), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n1225), .B(KEYINPUT124), .ZN(new_n1226));
  OR2_X1    g801(.A1(new_n1013), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n797), .A2(new_n799), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1218), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g804(.A1(new_n1218), .A2(G1986), .A3(G290), .ZN(new_n1230));
  AOI22_X1  g805(.A1(new_n1016), .A2(new_n1009), .B1(KEYINPUT48), .B2(new_n1230), .ZN(new_n1231));
  OR2_X1    g806(.A1(new_n1230), .A2(KEYINPUT48), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1229), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AND3_X1   g808(.A1(new_n1223), .A2(new_n1224), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1213), .A2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g810(.A1(G401), .A2(new_n465), .A3(G227), .ZN(new_n1237));
  AND3_X1   g811(.A1(new_n900), .A2(new_n706), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g812(.A(KEYINPUT127), .B1(new_n1238), .B2(new_n995), .ZN(new_n1239));
  NAND3_X1  g813(.A1(new_n900), .A2(new_n706), .A3(new_n1237), .ZN(new_n1240));
  INV_X1    g814(.A(new_n995), .ZN(new_n1241));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1242));
  NOR3_X1   g816(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NOR2_X1   g817(.A1(new_n1239), .A2(new_n1243), .ZN(G308));
  OR2_X1    g818(.A1(new_n1239), .A2(new_n1243), .ZN(G225));
endmodule


