//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n542, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT64), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n468), .B2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n463), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n468), .A2(G136), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n461), .B1(new_n465), .B2(new_n467), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(new_n461), .A2(G138), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n465), .B2(new_n467), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n470), .A2(new_n471), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n461), .A3(G138), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n461), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n479), .B2(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT65), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT65), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(G166));
  AND2_X1   g087(.A1(new_n506), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(G63), .A2(G651), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n513), .A2(G51), .B1(new_n502), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n502), .A2(new_n506), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(G89), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n517), .A2(new_n518), .A3(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  AOI22_X1  g100(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n504), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n513), .A2(G52), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT67), .B(G90), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  AOI22_X1  g108(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n504), .ZN(new_n535));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n507), .A2(new_n536), .B1(new_n509), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT68), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT69), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  INV_X1    g121(.A(G65), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n499), .B2(new_n501), .ZN(new_n548));
  AND2_X1   g123(.A1(G78), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n552), .B(G651), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n502), .A2(G91), .A3(new_n506), .ZN(new_n555));
  AND2_X1   g130(.A1(KEYINPUT6), .A2(G651), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n559));
  NOR2_X1   g134(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n506), .A2(G53), .A3(G543), .A4(new_n559), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n555), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n554), .A2(new_n565), .ZN(G299));
  OR2_X1    g141(.A1(new_n505), .A2(new_n511), .ZN(G303));
  OAI21_X1  g142(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n502), .A2(G87), .A3(new_n506), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n506), .A2(G49), .A3(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  INV_X1    g147(.A(G48), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n507), .A2(new_n572), .B1(new_n509), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n499), .B2(new_n501), .ZN(new_n576));
  AND2_X1   g151(.A1(G73), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(KEYINPUT72), .B(G651), .C1(new_n576), .C2(new_n577), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n574), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n519), .A2(G85), .B1(new_n513), .B2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n504), .B2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  XNOR2_X1  g162(.A(KEYINPUT73), .B(G66), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n502), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G79), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(new_n498), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n507), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G168), .B2(new_n602), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(G168), .B2(new_n602), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  INV_X1    g182(.A(new_n539), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n602), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n598), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g187(.A(new_n488), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n464), .A2(G2105), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT74), .B(G2100), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n616), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n468), .A2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n479), .A2(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n461), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G2096), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n619), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT75), .Z(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT76), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(G14), .B1(new_n640), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(KEYINPUT77), .B(KEYINPUT18), .Z(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  INV_X1    g228(.A(new_n646), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n653), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2096), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n660), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n660), .B2(new_n666), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1991), .B(G1996), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G229));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G19), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(new_n539), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT83), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1341), .ZN(new_n684));
  INV_X1    g259(.A(G29), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G26), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT86), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n468), .A2(G140), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT84), .ZN(new_n690));
  OAI21_X1  g265(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n691));
  INV_X1    g266(.A(G116), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G2105), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(KEYINPUT85), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(KEYINPUT85), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n694), .A2(new_n695), .B1(G128), .B2(new_n479), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n688), .B1(new_n697), .B2(G29), .ZN(new_n698));
  INV_X1    g273(.A(G2067), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT25), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n468), .A2(G139), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n613), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n702), .B(new_n703), .C1(new_n461), .C2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G33), .B(new_n705), .S(G29), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2072), .ZN(new_n707));
  INV_X1    g282(.A(G1961), .ZN(new_n708));
  NOR2_X1   g283(.A1(G171), .A2(new_n680), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G5), .B2(new_n680), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n707), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n712));
  INV_X1    g287(.A(G34), .ZN(new_n713));
  AOI21_X1  g288(.A(G29), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G160), .B2(new_n685), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2084), .ZN(new_n718));
  OAI22_X1  g293(.A1(new_n706), .A2(G2072), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR4_X1   g294(.A1(new_n684), .A2(new_n700), .A3(new_n711), .A4(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G4), .A2(G16), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n599), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT82), .ZN(new_n723));
  INV_X1    g298(.A(G1348), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n680), .A2(G20), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT23), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n564), .B1(new_n551), .B2(new_n553), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n680), .ZN(new_n730));
  INV_X1    g305(.A(G1956), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G168), .A2(new_n680), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n680), .B2(G21), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G162), .A2(new_n685), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n685), .B2(G35), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT29), .B(G2090), .Z(new_n739));
  AOI22_X1  g314(.A1(new_n738), .A2(new_n739), .B1(new_n718), .B2(new_n717), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n710), .B2(new_n708), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n685), .A2(G32), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n468), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n479), .A2(G129), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n614), .A2(G105), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n743), .B1(new_n751), .B2(new_n685), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT88), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n752), .B(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n736), .A2(new_n740), .A3(new_n742), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n685), .A2(G27), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n685), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2078), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G11), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT89), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(G28), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n685), .B1(new_n762), .B2(G28), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n761), .B1(new_n763), .B2(new_n764), .C1(new_n624), .C2(new_n685), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT90), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n734), .B2(new_n735), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n756), .A2(new_n759), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n726), .A2(new_n732), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n680), .A2(G6), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n582), .B2(new_n680), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT32), .B(G1981), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT80), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n680), .A2(G22), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n680), .ZN(new_n778));
  INV_X1    g353(.A(G1971), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G23), .B(G288), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT81), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n781), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n775), .A2(new_n776), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT79), .B(KEYINPUT34), .Z(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n680), .A2(G24), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G290), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G1986), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(G1986), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n468), .A2(G131), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n479), .A2(G119), .ZN(new_n795));
  OR2_X1    g370(.A1(G95), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G29), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G25), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT35), .B(G1991), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT78), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n801), .A2(new_n804), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n792), .A2(new_n793), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n787), .A2(new_n788), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT36), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT36), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n769), .B1(new_n809), .B2(new_n810), .ZN(G311));
  INV_X1    g386(.A(G311), .ZN(G150));
  AOI22_X1  g387(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n813), .A2(new_n814), .A3(new_n504), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n813), .B2(new_n504), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n519), .A2(G93), .B1(new_n513), .B2(G55), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G860), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  NOR2_X1   g395(.A1(new_n598), .A2(new_n606), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n818), .A2(new_n608), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n539), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n823), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT93), .ZN(new_n830));
  INV_X1    g405(.A(new_n827), .ZN(new_n831));
  AOI21_X1  g406(.A(G860), .B1(new_n831), .B2(KEYINPUT39), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n830), .A2(KEYINPUT94), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT94), .B1(new_n830), .B2(new_n832), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n820), .B1(new_n833), .B2(new_n834), .ZN(G145));
  XNOR2_X1  g410(.A(new_n495), .B(KEYINPUT95), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n705), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n616), .B(new_n798), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n697), .B(new_n750), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n468), .A2(G142), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n461), .A2(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n479), .A2(KEYINPUT96), .A3(G130), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT96), .B1(new_n479), .B2(G130), .ZN(new_n845));
  OAI221_X1 g420(.A(new_n841), .B1(new_n842), .B2(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n840), .B(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n839), .B(new_n847), .Z(new_n848));
  XOR2_X1   g423(.A(new_n624), .B(new_n476), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n839), .B(new_n847), .ZN(new_n852));
  INV_X1    g427(.A(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G37), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT97), .B(KEYINPUT40), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(G395));
  NAND2_X1  g433(.A1(new_n818), .A2(new_n602), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n824), .A2(new_n861), .A3(new_n825), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n824), .B2(new_n825), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n862), .A2(new_n863), .B1(G559), .B2(new_n598), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n826), .A2(KEYINPUT98), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n824), .A2(new_n861), .A3(new_n825), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n610), .A3(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(G299), .A2(new_n598), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n871));
  NAND2_X1  g446(.A1(G299), .A2(new_n598), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT41), .B1(new_n874), .B2(new_n869), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n874), .A2(new_n869), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(KEYINPUT99), .A3(new_n871), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n860), .B1(new_n868), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n868), .A2(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n864), .A2(new_n867), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n884), .A2(KEYINPUT100), .A3(new_n879), .A4(new_n877), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G166), .B(KEYINPUT101), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n887), .A2(new_n582), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(G288), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n582), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n886), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n881), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n883), .A2(new_n885), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT102), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n895), .B(KEYINPUT102), .C1(new_n897), .C2(new_n898), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n859), .B1(new_n902), .B2(new_n602), .ZN(G295));
  OAI21_X1  g478(.A(new_n859), .B1(new_n902), .B2(new_n602), .ZN(G331));
  NAND3_X1  g479(.A1(new_n824), .A2(G301), .A3(new_n825), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G301), .B1(new_n824), .B2(new_n825), .ZN(new_n907));
  OAI21_X1  g482(.A(G286), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n873), .A2(new_n875), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n826), .A2(G171), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(G168), .A3(new_n905), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n878), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(new_n908), .B2(new_n911), .ZN(new_n914));
  OAI22_X1  g489(.A1(new_n912), .A2(new_n914), .B1(new_n891), .B2(new_n892), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n906), .A2(new_n907), .A3(G286), .ZN(new_n916));
  AOI21_X1  g491(.A(G168), .B1(new_n910), .B2(new_n905), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n878), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n877), .A2(new_n908), .A3(new_n911), .A4(new_n879), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n893), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n915), .A2(new_n920), .A3(KEYINPUT43), .A4(new_n855), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n855), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n893), .B1(new_n918), .B2(new_n919), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT44), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n915), .A2(new_n920), .A3(new_n922), .A4(new_n855), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n923), .B2(new_n924), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n928), .A2(new_n929), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n927), .B1(new_n934), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g510(.A(KEYINPUT49), .ZN(new_n936));
  AOI211_X1 g511(.A(G1981), .B(new_n574), .C1(new_n580), .C2(new_n581), .ZN(new_n937));
  INV_X1    g512(.A(G1981), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n519), .A2(G86), .B1(new_n513), .B2(G48), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(new_n578), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n936), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n578), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(G1981), .ZN(new_n943));
  OAI211_X1 g518(.A(KEYINPUT49), .B(new_n943), .C1(G305), .C2(G1981), .ZN(new_n944));
  INV_X1    g519(.A(G8), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n469), .A2(new_n475), .A3(G40), .ZN(new_n946));
  AOI21_X1  g521(.A(G1384), .B1(new_n490), .B2(new_n494), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n941), .A2(new_n944), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G40), .ZN(new_n950));
  AOI211_X1 g525(.A(new_n950), .B(new_n462), .C1(new_n468), .C2(G137), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n495), .A2(new_n951), .A3(new_n952), .A4(new_n475), .ZN(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT107), .B(G1976), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT52), .B1(G288), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n568), .A2(new_n569), .A3(G1976), .A4(new_n570), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n953), .A2(G8), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT108), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n948), .A2(new_n959), .A3(new_n956), .A4(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n948), .A2(new_n956), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT52), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n949), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n946), .B1(new_n947), .B2(KEYINPUT45), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n966), .B(G1384), .C1(new_n490), .C2(new_n494), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n779), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n495), .A2(new_n952), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n970));
  INV_X1    g545(.A(G2090), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n947), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n970), .A2(new_n971), .A3(new_n946), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n976));
  NAND4_X1  g551(.A1(G303), .A2(new_n976), .A3(KEYINPUT55), .A4(G8), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT55), .B(G8), .C1(new_n505), .C2(new_n511), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT105), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G166), .B2(new_n945), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n975), .A2(G8), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT106), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n945), .B1(new_n968), .B2(new_n974), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n982), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n964), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(G288), .A2(G1976), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n937), .B1(new_n949), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n990), .A2(KEYINPUT109), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n948), .B1(new_n990), .B2(KEYINPUT109), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n984), .A2(new_n987), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n951), .A2(new_n475), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n969), .B2(new_n966), .ZN(new_n996));
  INV_X1    g571(.A(G2078), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n947), .A2(KEYINPUT45), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n495), .B2(new_n952), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n995), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n946), .B(KEYINPUT110), .C1(new_n947), .C2(KEYINPUT45), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1000), .A2(G2078), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n998), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n995), .B1(new_n969), .B2(KEYINPUT50), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n973), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n708), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1001), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n528), .A2(new_n1013), .A3(new_n529), .A4(new_n531), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n999), .A2(new_n1000), .B1(new_n1009), .B2(new_n708), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT121), .B1(new_n472), .B2(new_n473), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n1018));
  OAI21_X1  g593(.A(G2105), .B1(new_n474), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n951), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n951), .B(KEYINPUT122), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n998), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT123), .B(G2078), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1003), .A2(new_n1000), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1015), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1011), .A2(new_n1015), .B1(new_n1016), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n985), .A2(new_n982), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n994), .A2(new_n1028), .A3(new_n1029), .A4(new_n964), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n946), .B1(new_n947), .B2(new_n972), .ZN(new_n1031));
  AOI211_X1 g606(.A(KEYINPUT50), .B(G1384), .C1(new_n490), .C2(new_n494), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1031), .A2(G2084), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1004), .A2(new_n1005), .A3(new_n998), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(new_n735), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n945), .B1(new_n1035), .B2(G168), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n967), .B1(new_n965), .B2(new_n1002), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1966), .B1(new_n1039), .B2(new_n1005), .ZN(new_n1040));
  OAI211_X1 g615(.A(G8), .B(G286), .C1(new_n1040), .C2(new_n1033), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(KEYINPUT120), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1041), .B1(new_n1036), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1030), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1048), .A2(KEYINPUT57), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(KEYINPUT57), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n729), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n729), .B2(new_n1049), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(G299), .A2(new_n1048), .A3(KEYINPUT57), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n729), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n731), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n969), .A2(new_n966), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(new_n946), .A3(new_n998), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1062), .A3(KEYINPUT114), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1058), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1348), .B1(new_n1008), .B2(new_n973), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n953), .A2(G2067), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n599), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1059), .A2(new_n1062), .A3(new_n1056), .A4(new_n1054), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1072), .B(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1072), .A2(KEYINPUT61), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1067), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n724), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1069), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n598), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n599), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n965), .A2(G1996), .A3(new_n967), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(G1341), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n946), .B2(new_n947), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1996), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n996), .A2(new_n1092), .A3(new_n998), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1090), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT117), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT119), .B1(new_n1096), .B2(KEYINPUT59), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1091), .A2(new_n1095), .A3(new_n539), .A4(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1091), .A2(new_n539), .A3(new_n1095), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1097), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1077), .A2(new_n1085), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1063), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT61), .B1(new_n1074), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1075), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n993), .B1(new_n1047), .B2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1040), .A2(G286), .A3(new_n1033), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1037), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1107), .A2(new_n945), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT62), .B1(new_n1045), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1043), .B1(new_n1107), .B2(new_n945), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n1038), .A3(new_n1112), .A4(new_n1041), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n985), .A2(new_n986), .A3(new_n982), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n986), .B1(new_n985), .B2(new_n982), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n964), .B(new_n1029), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1011), .A2(G171), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1110), .A2(new_n1118), .A3(new_n1113), .A4(KEYINPUT124), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  OAI211_X1 g698(.A(G8), .B(G168), .C1(new_n1040), .C2(new_n1033), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1123), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n985), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n982), .B1(new_n1126), .B2(KEYINPUT111), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(KEYINPUT111), .B2(new_n1126), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1124), .A2(new_n1123), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(new_n994), .A3(new_n964), .A4(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1106), .A2(new_n1121), .A3(new_n1122), .A4(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1003), .A2(new_n946), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1092), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n750), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n697), .B(new_n699), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1092), .B2(new_n751), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT104), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1133), .B(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n798), .B(new_n804), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1140), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(G290), .B(G1986), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1134), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1132), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1141), .A2(new_n804), .A3(new_n799), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n690), .A2(new_n699), .A3(new_n696), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1150), .A2(KEYINPUT125), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(KEYINPUT125), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1143), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1137), .A2(new_n751), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1140), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT126), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1135), .B(KEYINPUT46), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(KEYINPUT47), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(KEYINPUT47), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1133), .A2(G1986), .A3(G290), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT48), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n1159), .A2(new_n1160), .B1(new_n1144), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1153), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1147), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g740(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1167), .A2(KEYINPUT127), .ZN(new_n1168));
  OR2_X1    g742(.A1(new_n1167), .A2(KEYINPUT127), .ZN(new_n1169));
  NAND4_X1  g743(.A1(new_n856), .A2(new_n678), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1170), .A2(new_n934), .ZN(G308));
  AND3_X1   g745(.A1(new_n678), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n1172), .B(new_n856), .C1(new_n933), .C2(new_n932), .ZN(G225));
endmodule


