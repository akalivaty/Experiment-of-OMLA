//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G101), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n188), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(KEYINPUT4), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G116), .ZN(new_n199));
  INV_X1    g013(.A(G116), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n203), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT4), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n193), .A2(new_n207), .A3(G101), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n197), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n187), .A2(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n190), .A2(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n196), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n199), .B2(KEYINPUT5), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT5), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT5), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n218), .A2(new_n198), .A3(KEYINPUT80), .A4(G116), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n216), .A2(new_n217), .A3(G113), .A4(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n214), .A2(new_n204), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G110), .B(G122), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n209), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n209), .A2(new_n221), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n222), .B(KEYINPUT81), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n223), .A2(KEYINPUT6), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n224), .A2(KEYINPUT6), .A3(new_n225), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n229), .B(G146), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  INV_X1    g045(.A(G125), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n233), .A3(G143), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g050(.A(G143), .B(G146), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n229), .A2(G146), .ZN(new_n241));
  AND4_X1   g055(.A1(new_n236), .A2(new_n238), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n235), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT82), .ZN(new_n244));
  OR2_X1    g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n240), .A2(new_n241), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n237), .B2(new_n251), .ZN(new_n252));
  AND4_X1   g066(.A1(new_n250), .A2(new_n240), .A3(new_n241), .A4(new_n251), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G125), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(new_n235), .C1(new_n239), .C2(new_n242), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n244), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(G224), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(G224), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n244), .A2(new_n255), .A3(new_n257), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(G902), .B1(new_n228), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(G210), .B1(G237), .B2(G902), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n265), .B(KEYINPUT86), .Z(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n222), .B(KEYINPUT8), .ZN(new_n268));
  AND4_X1   g082(.A1(new_n204), .A2(new_n220), .A3(new_n196), .A4(new_n212), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n220), .A2(new_n204), .B1(new_n196), .B2(new_n212), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT7), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n262), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n274), .A2(new_n272), .B1(new_n259), .B2(G224), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n274), .B2(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n258), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n258), .A2(KEYINPUT84), .A3(new_n276), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n273), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n223), .B1(new_n281), .B2(KEYINPUT85), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n262), .A2(new_n272), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n258), .A2(KEYINPUT84), .A3(new_n276), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT84), .B1(new_n258), .B2(new_n276), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n283), .B(new_n271), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n264), .B(new_n267), .C1(new_n282), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT87), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n264), .B1(new_n282), .B2(new_n288), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n266), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n287), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n281), .A2(KEYINPUT85), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n223), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT87), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n264), .A4(new_n267), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G214), .B1(G237), .B2(G902), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(G472), .A2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT32), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT11), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(G137), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(G137), .ZN(new_n310));
  INV_X1    g124(.A(G137), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT11), .A3(G134), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G131), .ZN(new_n314));
  INV_X1    g128(.A(G131), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n309), .A2(new_n312), .A3(new_n315), .A4(new_n310), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n231), .A2(new_n234), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT65), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n237), .A2(new_n236), .A3(new_n238), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n310), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n308), .A2(G137), .ZN(new_n324));
  OAI21_X1  g138(.A(G131), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n316), .ZN(new_n326));
  OAI22_X1  g140(.A1(new_n317), .A2(new_n254), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n206), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT30), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n327), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n318), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n239), .B2(new_n242), .ZN(new_n337));
  INV_X1    g151(.A(new_n326), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n314), .A2(new_n316), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n240), .A2(new_n241), .A3(new_n251), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT64), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n237), .A2(new_n250), .A3(new_n251), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n344), .A3(new_n249), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n339), .A2(new_n345), .A3(new_n329), .A4(new_n330), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n335), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n328), .B1(new_n347), .B2(new_n206), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT26), .B(G101), .Z(new_n349));
  NOR2_X1   g163(.A1(G237), .A2(G953), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G210), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n349), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n306), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n206), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n335), .B2(new_n346), .ZN(new_n357));
  INV_X1    g171(.A(new_n354), .ZN(new_n358));
  NOR4_X1   g172(.A1(new_n357), .A2(KEYINPUT31), .A3(new_n328), .A4(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n342), .A2(new_n343), .B1(new_n248), .B2(new_n247), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n337), .A2(new_n338), .B1(new_n362), .B2(new_n340), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n356), .B1(new_n363), .B2(KEYINPUT68), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n339), .A2(new_n345), .A3(KEYINPUT68), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n363), .A2(new_n356), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT28), .B1(new_n367), .B2(new_n328), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n358), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n305), .B1(new_n360), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g185(.A(new_n331), .B(new_n333), .C1(new_n339), .C2(new_n345), .ZN(new_n372));
  AND4_X1   g186(.A1(new_n329), .A2(new_n339), .A3(new_n330), .A4(new_n345), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n206), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n363), .A2(new_n356), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n354), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT31), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n348), .A2(new_n306), .A3(new_n354), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n377), .A2(new_n370), .A3(new_n305), .A4(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n304), .B1(new_n371), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G902), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n358), .B1(new_n366), .B2(new_n368), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n357), .A2(new_n328), .A3(new_n354), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT72), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n366), .A2(new_n387), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n368), .A2(KEYINPUT71), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n366), .A2(new_n387), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n368), .A2(KEYINPUT71), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n354), .A2(KEYINPUT29), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n382), .B(new_n386), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G472), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n377), .A2(new_n370), .A3(new_n378), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT69), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n302), .B1(new_n397), .B2(new_n379), .ZN(new_n398));
  XOR2_X1   g212(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n399));
  OAI211_X1 g213(.A(new_n381), .B(new_n395), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT9), .B(G234), .ZN(new_n401));
  OAI21_X1  g215(.A(G221), .B1(new_n401), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G469), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n259), .A2(G227), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT77), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G140), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g222(.A(KEYINPUT78), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n344), .A2(new_n249), .A3(new_n208), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n194), .A2(KEYINPUT4), .A3(new_n196), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n362), .A2(new_n197), .A3(KEYINPUT78), .A4(new_n208), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT10), .B1(new_n322), .B2(new_n213), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT10), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n337), .A2(new_n416), .A3(new_n214), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n414), .A2(new_n317), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n317), .B1(new_n414), .B2(new_n418), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT79), .B(new_n408), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n412), .A2(new_n413), .B1(new_n415), .B2(new_n417), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n408), .B1(new_n422), .B2(new_n317), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n337), .A2(new_n214), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n322), .A2(new_n213), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n317), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT12), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n344), .A2(new_n249), .A3(new_n208), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT78), .B1(new_n430), .B2(new_n197), .ZN(new_n431));
  AND4_X1   g245(.A1(KEYINPUT78), .A2(new_n362), .A3(new_n197), .A4(new_n208), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n418), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n340), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n422), .A2(new_n317), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT79), .B1(new_n436), .B2(new_n408), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n404), .B(new_n382), .C1(new_n429), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n427), .A2(new_n435), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n439), .A2(new_n408), .B1(new_n434), .B2(new_n423), .ZN(new_n440));
  OAI21_X1  g254(.A(G469), .B1(new_n440), .B2(G902), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n403), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G217), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n401), .A2(new_n447), .A3(G953), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT95), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n229), .B2(G128), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n230), .A2(KEYINPUT95), .A3(G143), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n230), .B2(G143), .ZN(new_n454));
  INV_X1    g268(.A(G122), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT94), .B1(new_n455), .B2(G116), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n200), .A3(G122), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n456), .A2(new_n458), .B1(G116), .B2(new_n455), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n454), .A2(new_n308), .B1(new_n459), .B2(new_n190), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n451), .A2(new_n452), .B1(G128), .B2(new_n229), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G134), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n456), .A2(new_n458), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n464), .A2(KEYINPUT14), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n464), .A2(KEYINPUT14), .B1(G116), .B2(new_n455), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n190), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT13), .B1(new_n451), .B2(new_n452), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n308), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n461), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n454), .B1(new_n469), .B2(new_n308), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n459), .A2(new_n190), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n459), .A2(new_n190), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n471), .A2(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n449), .B1(new_n468), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n465), .A2(new_n466), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n462), .B(new_n460), .C1(new_n477), .C2(new_n190), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n472), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n474), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n481), .A3(new_n448), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n446), .B1(new_n483), .B2(new_n382), .ZN(new_n484));
  AOI211_X1 g298(.A(G902), .B(new_n445), .C1(new_n476), .C2(new_n482), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n443), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n468), .A2(new_n475), .A3(new_n449), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n448), .B1(new_n478), .B2(new_n481), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n382), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n445), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n483), .A2(new_n382), .A3(new_n446), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT96), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(G234), .A2(G237), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(G952), .A3(new_n259), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT97), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n493), .A2(G902), .A3(G953), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n486), .A2(new_n492), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G475), .ZN(new_n501));
  INV_X1    g315(.A(G140), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G125), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n232), .A2(G140), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT16), .ZN(new_n505));
  OR3_X1    g319(.A1(new_n232), .A2(KEYINPUT16), .A3(G140), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(G146), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(G146), .B1(new_n505), .B2(new_n506), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT92), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n509), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n507), .ZN(new_n513));
  INV_X1    g327(.A(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n259), .A3(G214), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n229), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n350), .A2(G143), .A3(G214), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G131), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n315), .A3(new_n517), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(KEYINPUT17), .A3(G131), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n510), .A2(new_n513), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n503), .A2(new_n504), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n526), .B2(G146), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(G146), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n525), .A3(G146), .ZN(new_n530));
  INV_X1    g344(.A(new_n518), .ZN(new_n531));
  AND2_X1   g345(.A1(KEYINPUT18), .A2(G131), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n532), .B(KEYINPUT90), .Z(new_n533));
  AOI22_X1  g347(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n517), .ZN(new_n535));
  AOI21_X1  g349(.A(G143), .B1(new_n350), .B2(G214), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n518), .A2(KEYINPUT88), .A3(new_n532), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(G113), .B(G122), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(new_n187), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n524), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n524), .B2(new_n542), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n382), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n501), .B1(new_n547), .B2(KEYINPUT93), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n382), .C1(new_n545), .C2(new_n546), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(G475), .A2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n519), .A2(new_n521), .ZN(new_n553));
  XNOR2_X1  g367(.A(G125), .B(G140), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n554), .A2(KEYINPUT91), .A3(KEYINPUT19), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT19), .B1(new_n554), .B2(KEYINPUT91), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n553), .B(new_n507), .C1(new_n557), .C2(G146), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n544), .B1(new_n542), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n552), .B1(new_n545), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n542), .A2(new_n558), .ZN(new_n562));
  INV_X1    g376(.A(new_n544), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n524), .A2(new_n542), .A3(new_n544), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT20), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n552), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n551), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n500), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n442), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n198), .A2(G128), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n230), .A2(KEYINPUT23), .A3(G119), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n198), .A2(G128), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(KEYINPUT23), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n576), .A2(G110), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT73), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n230), .A2(G119), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n573), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT24), .B(G110), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n577), .A2(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n554), .A2(new_n233), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n507), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n511), .A2(new_n507), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n581), .A2(new_n582), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(G110), .B2(new_n576), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT22), .B(G137), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n591), .B(new_n592), .Z(new_n593));
  NAND3_X1  g407(.A1(new_n586), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n593), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n507), .A2(new_n585), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n579), .B2(new_n583), .ZN(new_n597));
  INV_X1    g411(.A(new_n590), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n594), .A2(new_n382), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT74), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n447), .B1(G234), .B2(new_n382), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n594), .A2(new_n599), .A3(KEYINPUT74), .A4(new_n382), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT25), .B1(new_n606), .B2(KEYINPUT75), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n604), .A2(G902), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT76), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n594), .A2(new_n599), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n300), .A2(new_n400), .A3(new_n572), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  OAI21_X1  g428(.A(new_n382), .B1(new_n371), .B2(new_n380), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n398), .B1(new_n615), .B2(G472), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n612), .A2(new_n442), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT98), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n301), .B1(new_n371), .B2(new_n380), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n397), .B2(new_n379), .ZN(new_n621));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n612), .A2(new_n442), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n263), .B1(new_n226), .B2(new_n227), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n382), .ZN(new_n629));
  INV_X1    g443(.A(new_n223), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n286), .B2(new_n287), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n266), .B(new_n629), .C1(new_n631), .C2(new_n294), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n267), .B1(new_n295), .B2(new_n264), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n299), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n489), .A2(new_n444), .ZN(new_n635));
  AND2_X1   g449(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n483), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n476), .B(new_n482), .C1(new_n639), .C2(new_n636), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n382), .A2(G478), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n635), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n570), .A2(new_n643), .A3(new_n499), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n627), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT100), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n567), .B1(new_n566), .B2(new_n552), .ZN(new_n651));
  INV_X1    g465(.A(new_n552), .ZN(new_n652));
  AOI211_X1 g466(.A(KEYINPUT20), .B(new_n652), .C1(new_n564), .C2(new_n565), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n561), .A2(new_n568), .A3(KEYINPUT101), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n486), .A2(new_n492), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n499), .B(KEYINPUT102), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n548), .B2(new_n550), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT103), .ZN(new_n662));
  INV_X1    g476(.A(new_n299), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n292), .B2(new_n289), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n656), .A2(new_n657), .A3(new_n665), .A4(new_n660), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n627), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT104), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NAND2_X1  g485(.A1(new_n586), .A2(new_n590), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n595), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n610), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n605), .B2(new_n607), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n300), .A2(new_n572), .A3(new_n616), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  INV_X1    g493(.A(new_n676), .ZN(new_n680));
  INV_X1    g494(.A(new_n399), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n620), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n397), .A2(new_n379), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n683), .A2(new_n304), .B1(new_n394), .B2(G472), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n656), .A2(new_n657), .ZN(new_n686));
  OR2_X1    g500(.A1(KEYINPUT105), .A2(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(KEYINPUT105), .A2(G900), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n496), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n495), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n548), .B2(new_n550), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n685), .A2(new_n442), .A3(new_n664), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  XNOR2_X1  g509(.A(new_n690), .B(KEYINPUT39), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n442), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT40), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n298), .B(KEYINPUT38), .Z(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n663), .A3(new_n676), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n699), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n354), .B1(new_n357), .B2(new_n328), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n367), .A2(new_n328), .ZN(new_n705));
  AOI21_X1  g519(.A(G902), .B1(new_n705), .B2(new_n358), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n622), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n683), .B2(new_n304), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n682), .A2(new_n708), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n551), .A2(new_n569), .B1(new_n486), .B2(new_n492), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n700), .A2(new_n702), .A3(new_n703), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND3_X1  g527(.A1(new_n570), .A2(new_n643), .A3(new_n690), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n685), .A2(new_n442), .A3(new_n664), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  OAI21_X1  g531(.A(new_n382), .B1(new_n429), .B2(new_n437), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n402), .A3(new_n438), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n400), .A2(new_n645), .A3(new_n612), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n667), .A2(new_n400), .A3(new_n612), .A4(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NOR2_X1   g540(.A1(new_n720), .A2(new_n634), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n400), .A3(new_n571), .A4(new_n676), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND3_X1  g543(.A1(new_n615), .A2(KEYINPUT107), .A3(G472), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n621), .B2(new_n622), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n710), .B(new_n299), .C1(new_n632), .C2(new_n633), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n734), .A2(new_n720), .A3(new_n659), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n392), .A2(new_n358), .ZN(new_n736));
  INV_X1    g550(.A(new_n360), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n301), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n733), .A2(new_n735), .A3(new_n612), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  NOR3_X1   g554(.A1(new_n720), .A2(new_n634), .A3(new_n714), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n733), .A2(new_n741), .A3(new_n676), .A4(new_n738), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NAND2_X1  g557(.A1(new_n381), .A2(new_n395), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n399), .B1(new_n683), .B2(new_n301), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n612), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n290), .A2(new_n297), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n633), .A2(new_n663), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n715), .A3(new_n442), .A4(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT108), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n612), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n682), .B2(new_n684), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n290), .A2(new_n292), .A3(new_n299), .A4(new_n297), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n438), .A2(new_n441), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n402), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n753), .A2(new_n755), .A3(new_n714), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n750), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n620), .A2(new_n303), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n751), .B1(new_n761), .B2(new_n684), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n756), .A3(KEYINPUT42), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(KEYINPUT109), .B(G131), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G33));
  NOR2_X1   g580(.A1(new_n753), .A2(new_n755), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n686), .B2(new_n692), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n768), .A2(new_n656), .A3(new_n657), .A4(new_n692), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n752), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND2_X1  g587(.A1(new_n440), .A2(KEYINPUT45), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n440), .A2(KEYINPUT45), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n404), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(G469), .A2(G902), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n438), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n783), .A2(KEYINPUT112), .B1(new_n782), .B2(new_n781), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(KEYINPUT112), .B2(new_n783), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(new_n402), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n696), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n643), .A2(new_n569), .A3(new_n551), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT43), .Z(new_n791));
  OR3_X1    g605(.A1(new_n791), .A2(new_n616), .A3(new_n680), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n753), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n793), .B2(new_n792), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(new_n311), .ZN(G39));
  NOR4_X1   g611(.A1(new_n400), .A2(new_n612), .A3(new_n714), .A4(new_n753), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  NAND3_X1  g616(.A1(new_n612), .A2(new_n299), .A3(new_n402), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n709), .A2(new_n788), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n719), .A2(new_n438), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT49), .Z(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n701), .A3(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n733), .A2(new_n738), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n791), .A2(new_n495), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n808), .A2(new_n809), .A3(new_n612), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n663), .A3(new_n701), .A4(new_n721), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT50), .Z(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n747), .A3(new_n721), .A4(new_n748), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n808), .A2(new_n676), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n753), .A2(new_n720), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n816), .A2(new_n709), .A3(new_n751), .A4(new_n495), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n570), .A2(new_n643), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n814), .A2(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n812), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n805), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n821), .A2(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(KEYINPUT117), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n822), .A2(new_n403), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n800), .A2(new_n799), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n810), .A2(new_n747), .A3(new_n748), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n820), .B(KEYINPUT51), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n814), .A2(new_n762), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT48), .ZN(new_n832));
  INV_X1    g646(.A(G952), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n570), .A2(new_n643), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n833), .B(G953), .C1(new_n817), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n727), .B2(new_n810), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n829), .A2(new_n830), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n613), .A2(new_n728), .A3(new_n677), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n725), .A2(new_n722), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n490), .A2(KEYINPUT114), .A3(new_n491), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT114), .B1(new_n490), .B2(new_n491), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n656), .A3(new_n692), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n844), .B1(new_n753), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n847), .A2(new_n656), .A3(new_n692), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n747), .A2(new_n850), .A3(KEYINPUT115), .A4(new_n748), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n685), .A2(new_n442), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n733), .A2(new_n756), .A3(new_n676), .A4(new_n738), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n852), .A2(new_n853), .A3(new_n772), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n569), .B(new_n551), .C1(new_n845), .C2(new_n846), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n659), .B1(new_n855), .B2(new_n834), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n856), .A2(new_n299), .A3(new_n298), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n618), .A2(new_n625), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(new_n739), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n764), .A2(new_n843), .A3(new_n854), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n634), .A2(new_n676), .A3(new_n691), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n709), .A2(new_n863), .A3(new_n442), .A4(new_n710), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n694), .A2(new_n716), .A3(new_n742), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n400), .A2(new_n442), .A3(new_n664), .A4(new_n676), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n693), .B2(new_n715), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT52), .A3(new_n742), .A4(new_n864), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n852), .A2(new_n853), .A3(new_n772), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n760), .B2(new_n763), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n858), .A2(new_n739), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n874), .A2(new_n841), .A3(new_n842), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(KEYINPUT116), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n862), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n871), .B1(new_n860), .B2(new_n861), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT116), .B1(new_n873), .B2(new_n875), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n840), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n875), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n867), .A2(new_n870), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n839), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n807), .B1(new_n890), .B2(new_n891), .ZN(G75));
  AOI21_X1  g706(.A(new_n886), .B1(new_n877), .B2(new_n878), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n382), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n894), .B2(new_n266), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n228), .B(KEYINPUT118), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(new_n263), .Z(new_n898));
  AND2_X1   g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n895), .A2(new_n898), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n833), .A2(G953), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT119), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(G51));
  AOI21_X1  g718(.A(KEYINPUT120), .B1(new_n893), .B2(new_n840), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n888), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n780), .B(KEYINPUT57), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n429), .A2(new_n437), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n894), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n779), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(KEYINPUT121), .A3(new_n902), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n910), .B2(new_n911), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n903), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(G54));
  NAND2_X1  g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT122), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n894), .A2(new_n566), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n566), .B1(new_n894), .B2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n903), .ZN(G60));
  INV_X1    g740(.A(new_n641), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT59), .ZN(new_n929));
  AND4_X1   g743(.A1(new_n927), .A2(new_n907), .A3(new_n908), .A4(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n883), .B2(new_n889), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n903), .B(new_n930), .C1(new_n641), .C2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  AND2_X1   g748(.A1(new_n888), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(new_n674), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n902), .B1(new_n935), .B2(new_n611), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT123), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g753(.A(G224), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n497), .A2(new_n940), .A3(new_n259), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n875), .B2(new_n259), .ZN(new_n942));
  INV_X1    g756(.A(new_n896), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(G898), .B2(new_n259), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n942), .B(new_n944), .ZN(G69));
  XNOR2_X1  g759(.A(new_n347), .B(new_n557), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n855), .A2(new_n834), .ZN(new_n948));
  OR4_X1    g762(.A1(new_n746), .A2(new_n948), .A3(new_n697), .A4(new_n753), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n787), .B2(new_n795), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n712), .A2(new_n742), .A3(new_n869), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT124), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n952), .A2(new_n801), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n947), .B1(new_n957), .B2(new_n259), .ZN(new_n958));
  AND2_X1   g772(.A1(G900), .A2(G953), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n946), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n869), .A2(new_n742), .ZN(new_n961));
  INV_X1    g775(.A(new_n787), .ZN(new_n962));
  INV_X1    g776(.A(new_n762), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n795), .B1(new_n734), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n965), .A2(new_n764), .A3(new_n772), .A4(new_n801), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n960), .B1(new_n966), .B2(G953), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n958), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n259), .B1(G227), .B2(G900), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n969), .B(new_n972), .ZN(G72));
  INV_X1    g787(.A(new_n875), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n957), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  AOI21_X1  g791(.A(new_n704), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n385), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n704), .A3(new_n977), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT127), .Z(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n879), .B2(new_n882), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n977), .B1(new_n966), .B2(new_n974), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(new_n385), .ZN(new_n984));
  NOR4_X1   g798(.A1(new_n978), .A2(new_n903), .A3(new_n982), .A4(new_n984), .ZN(G57));
endmodule


