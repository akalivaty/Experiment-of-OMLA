//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G250), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n204), .B1(new_n205), .B2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G13), .ZN(new_n207));
  NAND4_X1  g0007(.A1(new_n207), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n203), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n213), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(KEYINPUT0), .B2(new_n213), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n212), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G97), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n211), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n205), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n220), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(new_n214), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT69), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n261), .A2(G223), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n259), .ZN(new_n268));
  INV_X1    g0068(.A(G222), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n268), .A2(new_n269), .B1(new_n222), .B2(new_n267), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n255), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT68), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G33), .A3(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(new_n252), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n214), .B1(KEYINPUT68), .B2(new_n253), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(new_n274), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n281), .A2(G226), .B1(new_n284), .B2(new_n278), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G200), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n214), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT70), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n207), .A2(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n289), .A2(new_n294), .A3(new_n214), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G1), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(G50), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n291), .A2(new_n295), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n215), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(G150), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G20), .A2(G33), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n301), .A2(new_n302), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G50), .A2(G58), .ZN(new_n307));
  INV_X1    g0107(.A(G68), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n215), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n300), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n293), .ZN(new_n311));
  INV_X1    g0111(.A(G50), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n299), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT9), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n286), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT10), .B1(new_n288), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n271), .A2(new_n285), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G190), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n287), .A4(new_n315), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n286), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n325), .B(new_n314), .C1(G179), .C2(new_n286), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n301), .B1(new_n297), .B2(G20), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n296), .A2(new_n328), .B1(new_n311), .B2(new_n301), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT7), .B1(new_n258), .B2(new_n215), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n266), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n227), .A2(new_n308), .ZN(new_n334));
  NOR2_X1   g0134(.A1(G58), .A2(G68), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n304), .A2(G159), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT16), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n265), .A2(new_n215), .A3(new_n266), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n308), .B1(new_n343), .B2(new_n331), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n336), .A2(KEYINPUT16), .A3(new_n337), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n290), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n340), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n290), .ZN(new_n349));
  INV_X1    g0149(.A(new_n345), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n333), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n344), .B2(new_n338), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT76), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n329), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT18), .ZN(new_n356));
  INV_X1    g0156(.A(G223), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n259), .ZN(new_n358));
  INV_X1    g0158(.A(G226), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n358), .B(new_n360), .C1(new_n256), .C2(new_n257), .ZN(new_n361));
  AND3_X1   g0161(.A1(KEYINPUT77), .A2(G33), .A3(G87), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT77), .B1(G33), .B2(G87), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n255), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n275), .A2(G274), .A3(new_n278), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n275), .A2(G232), .A3(new_n279), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT78), .B1(new_n369), .B2(G179), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n324), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n255), .A2(new_n365), .B1(new_n284), .B2(new_n278), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT78), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .A4(new_n368), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n370), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n355), .A2(new_n356), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(G190), .B2(new_n369), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n329), .B(new_n381), .C1(new_n348), .C2(new_n354), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n329), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n347), .B1(new_n340), .B2(new_n346), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n351), .A2(KEYINPUT76), .A3(new_n353), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT18), .B1(new_n388), .B2(new_n376), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(KEYINPUT17), .A3(new_n381), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n378), .A2(new_n384), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n367), .B1(new_n280), .B2(new_n223), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n268), .A2(new_n228), .B1(new_n224), .B2(new_n267), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n261), .B2(G238), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n393), .B1(new_n395), .B2(new_n254), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G200), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n311), .A2(new_n290), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n222), .B1(new_n297), .B2(G20), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n398), .A2(new_n399), .B1(new_n222), .B2(new_n311), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT15), .B(G87), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n401), .A2(new_n302), .B1(new_n215), .B2(new_n222), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n301), .A2(new_n305), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n290), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT71), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n397), .B(new_n406), .C1(new_n316), .C2(new_n396), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n396), .A2(new_n324), .B1(new_n404), .B2(new_n400), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n374), .B(new_n393), .C1(new_n395), .C2(new_n254), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n327), .A2(new_n391), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n293), .A2(G68), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OR3_X1    g0214(.A1(new_n414), .A2(KEYINPUT74), .A3(KEYINPUT12), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT74), .B1(new_n414), .B2(KEYINPUT12), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(KEYINPUT12), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n305), .A2(new_n312), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n302), .A2(new_n222), .B1(new_n215), .B2(G68), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n300), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT11), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n398), .A2(G68), .A3(new_n298), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n422), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n418), .A2(new_n423), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT72), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n275), .A2(G238), .A3(new_n279), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n264), .A2(new_n229), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G226), .A2(G1698), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n228), .B2(G1698), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n431), .B1(new_n433), .B2(new_n267), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n430), .B(new_n367), .C1(new_n434), .C2(new_n254), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n429), .B1(new_n435), .B2(KEYINPUT13), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n228), .A2(G1698), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(G226), .B2(G1698), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n438), .A2(new_n258), .B1(new_n264), .B2(new_n229), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(new_n255), .B1(new_n284), .B2(new_n278), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT13), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n440), .A2(KEYINPUT72), .A3(new_n441), .A4(new_n430), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n436), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT14), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(G169), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT73), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n435), .B2(KEYINPUT13), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n440), .A2(KEYINPUT73), .A3(new_n441), .A4(new_n430), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(G179), .A4(new_n443), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n445), .B1(new_n444), .B2(G169), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n428), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n452), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT75), .A3(new_n450), .A4(new_n446), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n427), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n448), .A2(new_n449), .A3(G190), .A4(new_n443), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n444), .A2(G200), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n427), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n412), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n297), .B(G45), .C1(new_n276), .C2(KEYINPUT5), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n276), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n466), .B2(KEYINPUT82), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT82), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n276), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n467), .A2(new_n469), .B1(new_n274), .B2(new_n283), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n267), .A2(G250), .A3(new_n259), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G294), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n470), .A2(G264), .B1(new_n255), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n467), .A2(new_n284), .A3(new_n469), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n374), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n463), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT81), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n482));
  AOI21_X1  g0282(.A(G41), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n478), .B1(new_n483), .B2(new_n468), .ZN(new_n484));
  INV_X1    g0284(.A(new_n469), .ZN(new_n485));
  OAI211_X1 g0285(.A(G264), .B(new_n275), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n474), .A2(new_n255), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n476), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n324), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n297), .A2(G33), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n296), .A2(KEYINPUT80), .A3(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n291), .A2(new_n293), .A3(new_n490), .A4(new_n295), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT80), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n224), .B1(KEYINPUT89), .B2(KEYINPUT25), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n293), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G87), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(KEYINPUT88), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n267), .A2(new_n215), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n267), .A2(KEYINPUT22), .A3(new_n215), .A4(new_n504), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G116), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G20), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n215), .B2(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n224), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n507), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT24), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n507), .A2(new_n517), .A3(new_n508), .A4(new_n514), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n349), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n477), .B(new_n489), .C1(new_n502), .C2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G257), .B(new_n275), .C1(new_n484), .C2(new_n485), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT4), .A2(G244), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n259), .B(new_n522), .C1(new_n256), .C2(new_n257), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n223), .B1(new_n265), .B2(new_n266), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(KEYINPUT4), .ZN(new_n526));
  OAI21_X1  g0326(.A(G250), .B1(new_n256), .B2(new_n257), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n259), .B1(new_n527), .B2(KEYINPUT4), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n255), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n521), .A2(new_n529), .A3(new_n476), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n374), .ZN(new_n531));
  INV_X1    g0331(.A(new_n494), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n492), .A2(new_n493), .ZN(new_n533));
  OAI21_X1  g0333(.A(G97), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n311), .A2(new_n229), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n304), .A2(G77), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n536), .B(KEYINPUT79), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n538), .A2(new_n229), .A3(G107), .ZN(new_n539));
  XNOR2_X1  g0339(.A(G97), .B(G107), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n537), .B1(new_n215), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n224), .B1(new_n343), .B2(new_n331), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n290), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n534), .A2(new_n535), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n521), .A2(new_n529), .A3(new_n476), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n324), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n531), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n516), .A2(new_n518), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n290), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n475), .A2(G190), .A3(new_n476), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n500), .B1(new_n495), .B2(G107), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n488), .A2(G200), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n550), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n544), .A2(new_n535), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n546), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n521), .A2(new_n529), .A3(G190), .A4(new_n476), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n534), .A4(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n520), .A2(new_n548), .A3(new_n554), .A4(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n401), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n495), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT83), .ZN(new_n563));
  AOI21_X1  g0363(.A(G20), .B1(new_n431), .B2(KEYINPUT19), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n267), .A2(new_n215), .A3(G68), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n302), .A2(new_n229), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(KEYINPUT19), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n290), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n311), .A2(new_n401), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n561), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n259), .C1(new_n256), .C2(new_n257), .ZN(new_n572));
  OAI211_X1 g0372(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(new_n509), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n277), .A2(G1), .A3(G274), .ZN(new_n575));
  AOI21_X1  g0375(.A(G250), .B1(new_n297), .B2(G45), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n574), .A2(new_n255), .B1(new_n275), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(new_n324), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n255), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n275), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n580), .A2(G179), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n571), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n578), .A2(new_n379), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(G190), .B2(new_n578), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n569), .A2(new_n570), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT84), .B1(new_n495), .B2(G87), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT84), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n589), .B(new_n503), .C1(new_n491), .C2(new_n494), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n585), .B(new_n587), .C1(new_n588), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n559), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G270), .B(new_n275), .C1(new_n484), .C2(new_n485), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n595));
  OAI211_X1 g0395(.A(G257), .B(new_n259), .C1(new_n256), .C2(new_n257), .ZN(new_n596));
  XNOR2_X1  g0396(.A(KEYINPUT85), .B(G303), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n595), .B(new_n596), .C1(new_n267), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n255), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(new_n476), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT86), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n524), .B(new_n215), .C1(G33), .C2(new_n229), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(new_n290), .C1(new_n215), .C2(G116), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G116), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n297), .B2(G33), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n215), .A2(G116), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n398), .A2(new_n607), .B1(new_n608), .B2(new_n292), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n324), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT86), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n594), .A2(new_n611), .A3(new_n476), .A4(new_n599), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n601), .A2(KEYINPUT21), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT87), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n605), .A2(new_n609), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n616), .A2(new_n374), .A3(new_n600), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n601), .A2(new_n612), .A3(new_n610), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n601), .A2(new_n612), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G190), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n622), .B(new_n616), .C1(new_n379), .C2(new_n621), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n593), .A2(new_n615), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n462), .A2(new_n624), .ZN(G372));
  AOI21_X1  g0425(.A(KEYINPUT17), .B1(new_n388), .B2(new_n381), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n382), .A2(new_n383), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n453), .A2(new_n455), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n426), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT91), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n410), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n408), .A2(KEYINPUT91), .A3(new_n409), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n459), .A3(new_n632), .ZN(new_n633));
  AOI211_X1 g0433(.A(new_n626), .B(new_n627), .C1(new_n629), .C2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n378), .A2(new_n389), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n323), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(new_n326), .ZN(new_n638));
  INV_X1    g0438(.A(new_n462), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT90), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n579), .B2(new_n582), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n578), .A2(G179), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n642), .B(KEYINPUT90), .C1(new_n324), .C2(new_n578), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n571), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n613), .A2(new_n614), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n613), .A2(new_n614), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n620), .B(new_n520), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n591), .A2(new_n548), .A3(new_n558), .A4(new_n554), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n531), .A2(new_n545), .A3(new_n547), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n645), .A3(new_n591), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n583), .A3(new_n591), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n639), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n638), .A2(new_n659), .ZN(G369));
  NAND2_X1  g0460(.A1(new_n292), .A2(new_n215), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(G213), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n616), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n615), .A2(new_n623), .A3(new_n620), .A4(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n615), .A2(new_n620), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n669), .ZN(new_n672));
  XOR2_X1   g0472(.A(KEYINPUT92), .B(G330), .Z(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n520), .A2(new_n666), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n550), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n667), .B1(new_n550), .B2(new_n552), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n520), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n666), .B1(new_n615), .B2(new_n620), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n683), .A2(new_n676), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(G399));
  NOR2_X1   g0485(.A1(new_n210), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G1), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n563), .A2(new_n606), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n688), .A2(new_n689), .B1(new_n217), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n374), .B1(new_n598), .B2(new_n255), .ZN(new_n692));
  AND4_X1   g0492(.A1(new_n578), .A2(new_n692), .A3(new_n486), .A4(new_n487), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n694), .A2(new_n469), .A3(new_n478), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n470), .A2(G270), .B1(new_n695), .B2(new_n284), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n693), .A2(KEYINPUT30), .A3(new_n696), .A4(new_n530), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT95), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n486), .A2(new_n692), .A3(new_n487), .A4(new_n578), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n594), .A2(new_n476), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n700), .A2(new_n546), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n692), .A2(new_n578), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n696), .A3(new_n475), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT93), .B1(new_n706), .B2(new_n546), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT93), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n693), .A2(new_n708), .A3(new_n696), .A4(new_n530), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n578), .A2(G179), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n546), .A2(new_n488), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n621), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n704), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n693), .A2(new_n696), .A3(new_n530), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT30), .B1(new_n720), .B2(KEYINPUT93), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n714), .B1(new_n721), .B2(new_n709), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT96), .A3(new_n704), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n719), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n666), .ZN(new_n725));
  INV_X1    g0525(.A(new_n624), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n719), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n667), .A2(new_n719), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n722), .A2(KEYINPUT94), .B1(new_n699), .B2(new_n703), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n673), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n658), .A2(new_n667), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n495), .A2(G87), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n589), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n495), .A2(KEYINPUT84), .A3(G87), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n586), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n740), .A2(new_n585), .B1(new_n644), .B2(new_n571), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n654), .B1(new_n741), .B2(new_n652), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n656), .A2(KEYINPUT26), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n666), .B1(new_n744), .B2(new_n651), .ZN(new_n745));
  MUX2_X1   g0545(.A(new_n736), .B(new_n745), .S(KEYINPUT29), .Z(new_n746));
  AND2_X1   g0546(.A1(new_n735), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n691), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n207), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n688), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n209), .A2(G355), .A3(new_n267), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n247), .A2(new_n277), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n209), .B(new_n258), .C1(G45), .C2(new_n217), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n754), .B1(G116), .B2(new_n209), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n214), .B1(G20), .B2(new_n324), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(G20), .A2(G179), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n316), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n215), .A2(G179), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(new_n316), .A3(G200), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n768), .A2(new_n312), .B1(new_n770), .B2(new_n224), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n771), .B1(G87), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n764), .A2(new_n316), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n267), .B1(new_n776), .B2(new_n227), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G190), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n765), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n777), .B1(G77), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n769), .A2(new_n778), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G159), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT32), .Z(new_n785));
  NOR2_X1   g0585(.A1(new_n766), .A2(G190), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n374), .A2(new_n379), .A3(G190), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n786), .A2(G68), .B1(G97), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n774), .A2(new_n781), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G329), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n782), .A2(new_n791), .B1(new_n779), .B2(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n267), .B(new_n793), .C1(G322), .C2(new_n775), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n772), .B(KEYINPUT98), .Z(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G303), .ZN(new_n796));
  INV_X1    g0596(.A(new_n770), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n797), .A2(G283), .B1(new_n788), .B2(G294), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G326), .A2(new_n767), .B1(new_n786), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n794), .A2(new_n796), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n790), .A2(KEYINPUT99), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT99), .B1(new_n790), .B2(new_n801), .ZN(new_n803));
  INV_X1    g0603(.A(new_n761), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n753), .B(new_n763), .C1(new_n802), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT100), .ZN(new_n807));
  INV_X1    g0607(.A(new_n760), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n672), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n672), .A2(new_n673), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT97), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n674), .A2(new_n753), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT101), .ZN(G396));
  NOR2_X1   g0614(.A1(new_n411), .A2(new_n666), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n658), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n736), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n631), .A2(new_n405), .A3(new_n632), .A4(new_n666), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n405), .A2(new_n666), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n407), .A2(new_n410), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n816), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n752), .B1(new_n735), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n735), .B2(new_n822), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n804), .A2(new_n759), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n752), .B1(G77), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n776), .A2(new_n827), .B1(new_n779), .B2(new_n606), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n267), .B(new_n828), .C1(G311), .C2(new_n783), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n795), .A2(G107), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n770), .A2(new_n503), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G97), .B2(new_n788), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G283), .A2(new_n786), .B1(new_n767), .B2(G303), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n829), .A2(new_n830), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n780), .A2(G159), .B1(G143), .B2(new_n775), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  INV_X1    g0636(.A(new_n786), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n768), .B2(new_n836), .C1(new_n303), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(KEYINPUT102), .B(KEYINPUT34), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n795), .A2(G50), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n267), .B1(new_n782), .B2(new_n842), .C1(new_n308), .C2(new_n770), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G58), .B2(new_n788), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n840), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n838), .A2(new_n839), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n834), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n826), .B1(new_n847), .B2(new_n761), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n821), .B2(new_n759), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n824), .A2(new_n849), .ZN(G384));
  INV_X1    g0650(.A(new_n541), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n851), .A2(KEYINPUT35), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(KEYINPUT35), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(G116), .A3(new_n216), .A4(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT36), .Z(new_n855));
  OAI211_X1 g0655(.A(new_n218), .B(G77), .C1(new_n227), .C2(new_n308), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n312), .A2(G68), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n297), .B(G13), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT108), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n382), .B1(new_n388), .B2(new_n376), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n388), .A2(new_n664), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n862), .A2(KEYINPUT37), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n352), .A2(KEYINPUT104), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n344), .B2(new_n338), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n333), .A2(new_n339), .A3(new_n865), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n300), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n329), .ZN(new_n870));
  AND4_X1   g0670(.A1(new_n374), .A2(new_n366), .A3(new_n367), .A4(new_n368), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n871), .A2(new_n373), .B1(new_n324), .B2(new_n369), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n872), .A3(new_n370), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n382), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n382), .A2(new_n873), .A3(KEYINPUT106), .ZN(new_n877));
  INV_X1    g0677(.A(new_n664), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT105), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n880), .B(new_n664), .C1(new_n869), .C2(new_n329), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n876), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n864), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n627), .A2(new_n626), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n635), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n861), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n300), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n333), .A2(new_n339), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n866), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n385), .B1(new_n890), .B2(new_n868), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n880), .B1(new_n891), .B2(new_n664), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n870), .A2(KEYINPUT105), .A3(new_n878), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n391), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT106), .B1(new_n382), .B2(new_n873), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n894), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n898), .B2(new_n877), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT38), .B(new_n895), .C1(new_n899), .C2(new_n864), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n887), .A2(new_n900), .A3(KEYINPUT39), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n629), .A2(new_n666), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n862), .B2(new_n863), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n355), .A2(new_n377), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n355), .A2(new_n878), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n896), .A4(new_n382), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n391), .A2(new_n863), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n886), .B1(new_n910), .B2(new_n906), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n909), .B1(new_n911), .B2(KEYINPUT38), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n901), .B(new_n902), .C1(new_n912), .C2(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n636), .A2(new_n664), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n427), .A2(new_n667), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n629), .A2(new_n459), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n916), .B1(new_n456), .B2(new_n460), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n815), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n651), .B2(new_n657), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n408), .A2(new_n409), .A3(new_n667), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT103), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n920), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n887), .A2(new_n900), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT107), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n887), .A2(new_n900), .A3(KEYINPUT107), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n860), .B1(new_n915), .B2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n816), .A2(new_n924), .B1(new_n918), .B2(new_n919), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n887), .A2(KEYINPUT107), .A3(new_n900), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT107), .B1(new_n887), .B2(new_n900), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n936), .A2(KEYINPUT108), .A3(new_n914), .A4(new_n913), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n638), .B1(new_n746), .B2(new_n462), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n938), .B(new_n939), .Z(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n934), .A2(new_n935), .ZN(new_n942));
  INV_X1    g0742(.A(new_n821), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n918), .B2(new_n919), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n718), .A2(new_n723), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT109), .B1(new_n945), .B2(new_n728), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT109), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n947), .B(new_n729), .C1(new_n718), .C2(new_n723), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n724), .A2(new_n666), .B1(new_n624), .B2(KEYINPUT31), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n941), .B1(new_n942), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n909), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n941), .B1(new_n953), .B2(new_n900), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n954), .B(new_n944), .C1(new_n949), .C2(new_n950), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n716), .A2(new_n717), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT96), .B1(new_n722), .B2(new_n704), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n728), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n947), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n945), .A2(KEYINPUT109), .A3(new_n728), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n950), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n462), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n956), .A2(new_n963), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n673), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n940), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n297), .B2(new_n749), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n940), .A2(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n859), .B1(new_n968), .B2(new_n969), .ZN(G367));
  NAND2_X1  g0770(.A1(new_n652), .A2(new_n666), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n545), .A2(new_n666), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n558), .A2(new_n548), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n680), .A2(new_n682), .A3(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n548), .B1(new_n973), .B2(new_n520), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n975), .A2(KEYINPUT42), .B1(new_n667), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n740), .A2(new_n667), .ZN(new_n979));
  MUX2_X1   g0779(.A(new_n741), .B(new_n646), .S(new_n979), .Z(new_n980));
  AOI22_X1  g0780(.A1(new_n976), .A2(new_n978), .B1(new_n980), .B2(KEYINPUT43), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n681), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n974), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n983), .B(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n751), .A2(new_n297), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n686), .B(KEYINPUT41), .Z(new_n988));
  NAND3_X1  g0788(.A1(new_n683), .A2(new_n676), .A3(new_n974), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n684), .B2(new_n974), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n683), .A2(new_n676), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n995), .A2(KEYINPUT44), .A3(new_n973), .A4(new_n971), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT45), .B1(new_n990), .B2(new_n991), .ZN(new_n999));
  OAI211_X1 g0799(.A(KEYINPUT111), .B(new_n984), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n999), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n984), .A2(KEYINPUT111), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n1001), .A2(new_n1002), .A3(new_n992), .A4(new_n997), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n680), .B(new_n682), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n675), .B(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1000), .A2(new_n1003), .A3(new_n747), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n988), .B1(new_n1006), .B2(new_n747), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT112), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n987), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(KEYINPUT112), .B(new_n988), .C1(new_n1006), .C2(new_n747), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n986), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT113), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(KEYINPUT113), .B(new_n986), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n242), .A2(new_n209), .A3(new_n258), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n762), .B1(new_n209), .B2(new_n401), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n752), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n606), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n795), .A2(G116), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(KEYINPUT46), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G294), .A2(new_n786), .B1(new_n797), .B2(G97), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n597), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n267), .B1(new_n1023), .B2(new_n775), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n767), .A2(G311), .B1(G107), .B2(new_n788), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G317), .A2(new_n783), .B1(new_n780), .B2(G283), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n776), .A2(new_n303), .B1(new_n782), .B2(new_n836), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G50), .B2(new_n780), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n773), .A2(G58), .B1(new_n788), .B2(G68), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G143), .A2(new_n767), .B1(new_n786), .B2(G159), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n267), .B1(new_n770), .B2(new_n222), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT114), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1021), .A2(new_n1027), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1018), .B1(new_n1036), .B2(new_n761), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n980), .B2(new_n808), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT115), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1015), .A2(new_n1040), .ZN(G387));
  INV_X1    g0841(.A(new_n987), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1005), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n680), .A2(new_n808), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n301), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n1045), .A2(KEYINPUT50), .A3(new_n312), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT50), .B1(new_n1045), .B2(new_n312), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n277), .B1(new_n308), .B2(new_n222), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n689), .B1(new_n1048), .B2(new_n258), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n267), .A2(new_n277), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1049), .B1(new_n238), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1051), .A2(new_n210), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n762), .B1(new_n224), .B2(new_n209), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n780), .A2(new_n1023), .B1(G317), .B2(new_n775), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n767), .A2(G322), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n792), .C2(new_n837), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT48), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n773), .A2(G294), .B1(new_n788), .B2(G283), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n770), .A2(new_n606), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n267), .B(new_n1065), .C1(G326), .C2(new_n783), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n776), .A2(new_n312), .B1(new_n779), .B2(new_n308), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n258), .B(new_n1068), .C1(G150), .C2(new_n783), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n786), .A2(new_n1045), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n767), .A2(G159), .B1(new_n560), .B2(new_n788), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n773), .A2(G77), .B1(new_n797), .B2(G97), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT116), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n752), .B1(new_n1052), .B2(new_n1053), .C1(new_n1075), .C2(new_n804), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n747), .A2(new_n1005), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n686), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n747), .A2(new_n1005), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1043), .B1(new_n1044), .B2(new_n1076), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT117), .ZN(G393));
  NOR2_X1   g0881(.A1(new_n681), .A2(KEYINPUT118), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n998), .A2(new_n999), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT118), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n984), .ZN(new_n1085));
  OAI211_X1 g0885(.A(KEYINPUT118), .B(new_n681), .C1(new_n998), .C2(new_n999), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1077), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n686), .A3(new_n1006), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n209), .A2(new_n258), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n762), .B1(new_n229), .B2(new_n209), .C1(new_n250), .C2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n752), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n974), .A2(new_n808), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n767), .A2(G317), .B1(G311), .B2(new_n775), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT52), .Z(new_n1094));
  OAI21_X1  g0894(.A(new_n258), .B1(new_n779), .B2(new_n827), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G322), .B2(new_n783), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n797), .A2(G107), .B1(new_n788), .B2(G116), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1023), .A2(new_n786), .B1(new_n773), .B2(G283), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n767), .A2(G150), .B1(G159), .B2(new_n775), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT51), .Z(new_n1101));
  AOI211_X1 g0901(.A(new_n258), .B(new_n831), .C1(G143), .C2(new_n783), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n308), .C2(new_n772), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n788), .A2(G77), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n301), .B2(new_n779), .C1(new_n837), .C2(new_n312), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT119), .Z(new_n1106));
  OAI21_X1  g0906(.A(new_n1099), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1091), .B(new_n1092), .C1(new_n761), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n1042), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1088), .A2(new_n1110), .ZN(G390));
  OAI21_X1  g0911(.A(new_n752), .B1(new_n1045), .B2(new_n825), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n782), .A2(new_n827), .B1(new_n779), .B2(new_n229), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n267), .B(new_n1113), .C1(G116), .C2(new_n775), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n795), .A2(G87), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n797), .A2(G68), .B1(new_n788), .B2(G77), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G107), .A2(new_n786), .B1(new_n767), .B2(G283), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G128), .A2(new_n767), .B1(new_n797), .B2(G50), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n786), .A2(G137), .B1(G159), .B2(new_n788), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1122));
  OR3_X1    g0922(.A1(new_n1122), .A2(new_n772), .A3(new_n303), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G125), .A2(new_n783), .B1(new_n780), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1122), .B1(new_n772), .B2(new_n303), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n258), .B1(G132), .B2(new_n775), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1123), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1118), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1130), .A2(KEYINPUT122), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n804), .B1(new_n1130), .B2(KEYINPUT122), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1112), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n901), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT39), .B1(new_n953), .B2(new_n900), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1133), .B1(new_n1136), .B2(new_n759), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT123), .ZN(new_n1138));
  OAI211_X1 g0938(.A(G330), .B(new_n944), .C1(new_n949), .C2(new_n950), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT39), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n884), .A2(new_n861), .A3(new_n886), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n909), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n902), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1143), .A2(new_n901), .B1(new_n926), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1142), .B2(new_n909), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT120), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n917), .B1(new_n629), .B2(new_n459), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n456), .A2(new_n460), .A3(new_n916), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n918), .A2(KEYINPUT120), .A3(new_n919), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n744), .A2(new_n651), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n667), .A3(new_n821), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n924), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1146), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1140), .B1(new_n1145), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1151), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT120), .B1(new_n918), .B2(new_n919), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1146), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1134), .A2(new_n1135), .B1(new_n933), .B2(new_n902), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n734), .A2(new_n673), .A3(new_n821), .A4(new_n920), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1157), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n1042), .ZN(new_n1168));
  OAI21_X1  g0968(.A(G330), .B1(new_n949), .B2(new_n950), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1151), .B(new_n1150), .C1(new_n1169), .C2(new_n943), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n673), .B(new_n821), .C1(new_n950), .C2(new_n732), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1155), .B1(new_n1172), .B2(new_n920), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n920), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n1139), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n816), .A2(new_n924), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1170), .A2(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(G330), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n962), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n639), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n638), .C1(new_n462), .C2(new_n746), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n686), .B1(new_n1183), .B2(new_n1167), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1169), .A2(new_n462), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n939), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(new_n1166), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1138), .B(new_n1168), .C1(new_n1184), .C2(new_n1191), .ZN(G378));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n1178), .B2(new_n1166), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n929), .A2(new_n930), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n821), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n960), .A2(new_n961), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n727), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT40), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n955), .A2(G330), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n314), .A2(new_n878), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n327), .B(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1201), .B(new_n1203), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1198), .A2(new_n1199), .A3(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1201), .B(new_n1202), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1179), .B1(new_n1197), .B2(new_n954), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1206), .B1(new_n952), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n938), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1204), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n952), .A2(new_n1207), .A3(new_n1206), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n932), .A4(new_n937), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1193), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1193), .A2(new_n1209), .A3(KEYINPUT57), .A4(new_n1212), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n686), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1209), .A2(new_n1042), .A3(new_n1212), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n752), .B1(G50), .B2(new_n825), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n837), .A2(new_n229), .B1(new_n770), .B2(new_n227), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G116), .B2(new_n767), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n258), .A2(new_n276), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G283), .B2(new_n783), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n780), .A2(new_n560), .B1(G107), .B2(new_n775), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n773), .A2(G77), .B1(new_n788), .B2(G68), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT58), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1223), .B(new_n312), .C1(G33), .C2(G41), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n767), .A2(G125), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n837), .B2(new_n842), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n780), .A2(G137), .B1(G128), .B2(new_n775), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n772), .B2(new_n1124), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(G150), .C2(new_n788), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n797), .A2(G159), .ZN(new_n1239));
  AOI211_X1 g1039(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1231), .B1(new_n1228), .B2(new_n1227), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1220), .B1(new_n1243), .B2(new_n761), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1206), .B2(new_n759), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1219), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1218), .A2(new_n1246), .ZN(G375));
  NOR2_X1   g1047(.A1(new_n1183), .A2(new_n988), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1189), .B2(new_n1187), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1152), .A2(new_n759), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT124), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n752), .B1(G68), .B2(new_n825), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n776), .A2(new_n836), .B1(new_n779), .B2(new_n303), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n258), .B(new_n1253), .C1(G128), .C2(new_n783), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n795), .A2(G159), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n797), .A2(G58), .B1(new_n788), .B2(G50), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G132), .A2(new_n767), .B1(new_n786), .B2(new_n1125), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n775), .A2(G283), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n224), .B2(new_n779), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n267), .B(new_n1260), .C1(G303), .C2(new_n783), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n795), .A2(G97), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n797), .A2(G77), .B1(new_n560), .B2(new_n788), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G116), .A2(new_n786), .B1(new_n767), .B2(G294), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1258), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1252), .B1(new_n1266), .B2(new_n761), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1187), .A2(new_n1042), .B1(new_n1251), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1249), .A2(new_n1268), .ZN(G381));
  AOI211_X1 g1069(.A(new_n1039), .B(G390), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1168), .A2(new_n1138), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1184), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1191), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(G375), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1270), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(G407));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n665), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G375), .C2(new_n1278), .ZN(G409));
  NAND2_X1  g1079(.A1(G387), .A2(G390), .ZN(new_n1280));
  INV_X1    g1080(.A(G390), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1015), .A2(new_n1040), .A3(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G393), .B(G396), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(new_n1282), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1281), .B1(new_n1015), .B2(new_n1040), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1283), .B1(new_n1286), .B2(new_n1270), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(G213), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(G343), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1209), .A2(KEYINPUT125), .A3(new_n1212), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1042), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT125), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1245), .B1(new_n1213), .B2(new_n988), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1274), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G378), .B(new_n1246), .C1(new_n1215), .C2(new_n1217), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1290), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n686), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT60), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT60), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1178), .A2(new_n1182), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1300), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(G384), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1268), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n687), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1303), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1302), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1311), .B2(new_n1268), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1299), .B1(new_n1307), .B2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1305), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1311), .A2(G384), .A3(new_n1268), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(KEYINPUT126), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT62), .B1(new_n1298), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1290), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  AOI211_X1 g1122(.A(KEYINPUT127), .B(new_n1290), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1318), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1290), .A2(G2897), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1317), .B2(new_n1327), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1288), .B1(new_n1326), .B2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1317), .A2(KEYINPUT63), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1324), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1298), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1329), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT63), .B1(new_n1298), .B2(new_n1317), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1339), .A2(KEYINPUT61), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1334), .A2(new_n1336), .A3(new_n1338), .A4(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1333), .A2(new_n1341), .ZN(G405));
  NAND2_X1  g1142(.A1(G375), .A2(new_n1274), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1297), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1317), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1307), .A2(new_n1312), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1334), .B(new_n1345), .C1(new_n1346), .C2(new_n1344), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1345), .B1(new_n1346), .B2(new_n1344), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1288), .A2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(G402));
endmodule


