//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(new_n456), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n465), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .A3(G137), .A4(new_n469), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n474), .A2(new_n478), .A3(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n468), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n469), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n472), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(new_n472), .B2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n493), .B2(G124), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT71), .ZN(G162));
  NAND2_X1  g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n469), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n505), .A2(new_n507), .A3(G2104), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(G138), .B(new_n469), .C1(new_n466), .C2(new_n467), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n472), .A2(new_n513), .A3(G138), .A4(new_n469), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n503), .A2(new_n510), .B1(new_n512), .B2(new_n514), .ZN(G164));
  OAI21_X1  g090(.A(KEYINPUT5), .B1(KEYINPUT74), .B2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT75), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(KEYINPUT74), .A2(KEYINPUT75), .A3(KEYINPUT5), .A4(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n525), .B1(new_n522), .B2(KEYINPUT73), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(KEYINPUT6), .A3(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(new_n528), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n523), .A2(new_n534), .ZN(G166));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n540), .A2(new_n542), .B1(G51), .B2(new_n529), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n518), .A2(new_n519), .B1(new_n526), .B2(new_n528), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT78), .B(G89), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT76), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT79), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n548), .B(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n552), .A2(new_n553), .A3(new_n546), .A4(new_n543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n550), .A2(new_n554), .ZN(G168));
  AOI22_X1  g130(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n522), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n529), .A2(G52), .ZN(new_n558));
  INV_X1    g133(.A(G90), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n532), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(G171));
  AOI22_X1  g136(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OR3_X1    g137(.A1(new_n562), .A2(KEYINPUT80), .A3(new_n522), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT80), .B1(new_n562), .B2(new_n522), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n544), .A2(G81), .B1(G43), .B2(new_n529), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n529), .A2(new_n573), .A3(G53), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n573), .B1(new_n529), .B2(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT81), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n576), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(new_n579), .A3(new_n574), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(new_n520), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G91), .B2(new_n544), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n581), .A2(new_n586), .ZN(G299));
  INV_X1    g162(.A(G171), .ZN(G301));
  INV_X1    g163(.A(G168), .ZN(G286));
  OR2_X1    g164(.A1(new_n523), .A2(new_n534), .ZN(G303));
  INV_X1    g165(.A(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n518), .A2(new_n591), .A3(new_n519), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n529), .A2(G49), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n596));
  INV_X1    g171(.A(G87), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n532), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n544), .A2(KEYINPUT82), .A3(G87), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G288));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n518), .B2(new_n519), .ZN(new_n603));
  AND2_X1   g178(.A1(G73), .A2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT83), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n607), .B(G651), .C1(new_n603), .C2(new_n604), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n544), .A2(G86), .B1(G48), .B2(new_n529), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(G305));
  AND2_X1   g185(.A1(new_n520), .A2(G60), .ZN(new_n611));
  AND2_X1   g186(.A1(G72), .A2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n544), .A2(G85), .B1(G47), .B2(new_n529), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n544), .A2(G92), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT10), .Z(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  INV_X1    g197(.A(G66), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n583), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n624), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n619), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n619), .B1(new_n627), .B2(G868), .ZN(G321));
  NOR2_X1   g204(.A1(G299), .A2(G868), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g206(.A(new_n630), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n627), .B1(new_n633), .B2(G860), .ZN(G148));
  OAI21_X1  g209(.A(G868), .B1(new_n626), .B2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n472), .A2(new_n480), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(G111), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(G2105), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n483), .B2(G135), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n493), .B2(G123), .ZN(new_n648));
  AOI22_X1  g223(.A1(new_n640), .A2(new_n641), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G2096), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n649), .B(new_n651), .C1(new_n641), .C2(new_n640), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(G156));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n657), .B(new_n663), .Z(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n667), .A3(G14), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT86), .Z(G401));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT17), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(new_n670), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT87), .Z(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(new_n672), .A3(new_n670), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT18), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n672), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n671), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT89), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(KEYINPUT89), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT20), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n687), .A3(new_n688), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n687), .B(new_n688), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n697), .B(new_n698), .C1(new_n694), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT91), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(G1981), .B(G1986), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT90), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n703), .B(new_n707), .ZN(G229));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G25), .ZN(new_n710));
  INV_X1    g285(.A(G119), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n492), .A2(KEYINPUT92), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT92), .B1(new_n492), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(G107), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G2105), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n483), .B2(G131), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n710), .B1(new_n719), .B2(new_n709), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n723), .A2(G24), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G290), .B2(G16), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n722), .B1(G1986), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n600), .A2(new_n723), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n723), .B2(G23), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT33), .B(G1976), .Z(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n723), .A2(G22), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G166), .B2(new_n723), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(G1971), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(G1971), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n732), .A2(new_n733), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G6), .B(G305), .S(G16), .Z(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT32), .B(G1981), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT34), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n738), .A2(KEYINPUT34), .A3(new_n741), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n726), .A2(G1986), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n727), .A2(new_n742), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT36), .Z(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G35), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G162), .B2(G29), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT29), .Z(new_n749));
  INV_X1    g324(.A(G2090), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n723), .A2(G19), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n567), .B2(new_n723), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1341), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n723), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n751), .A2(new_n752), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT31), .B(G11), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT100), .B(G28), .Z(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n762), .B2(KEYINPUT30), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(KEYINPUT101), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(KEYINPUT101), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(KEYINPUT30), .B2(new_n762), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n761), .B1(new_n764), .B2(new_n766), .C1(new_n650), .C2(new_n709), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT102), .Z(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT98), .B(KEYINPUT26), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G105), .B2(new_n480), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n483), .A2(G141), .ZN(new_n773));
  INV_X1    g348(.A(G129), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n772), .B(new_n773), .C1(new_n774), .C2(new_n492), .ZN(new_n775));
  MUX2_X1   g350(.A(G32), .B(new_n775), .S(G29), .Z(new_n776));
  XOR2_X1   g351(.A(KEYINPUT27), .B(G1996), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G164), .A2(new_n709), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G27), .B2(new_n709), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(G160), .A2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n785), .B2(KEYINPUT24), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT24), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2084), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n778), .A2(new_n782), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n709), .A2(G26), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT94), .ZN(new_n796));
  INV_X1    g371(.A(G116), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n479), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  AOI22_X1  g373(.A1(G140), .A2(new_n483), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G128), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n492), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n794), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  NOR2_X1   g378(.A1(G171), .A2(new_n723), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G5), .B2(new_n723), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n803), .B1(new_n806), .B2(G1961), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n768), .A2(new_n791), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G16), .A2(G21), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G168), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G1966), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n806), .A2(G1961), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT103), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n723), .A2(G4), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n627), .B2(new_n723), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT93), .B(G1348), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n808), .A2(new_n812), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n709), .A2(G33), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT25), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n483), .A2(G139), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n469), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n820), .B1(new_n827), .B2(new_n709), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT96), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G2072), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT97), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(G2072), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n776), .A2(new_n777), .B1(new_n789), .B2(new_n788), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT99), .Z(new_n836));
  NOR4_X1   g411(.A1(new_n746), .A2(new_n760), .A3(new_n819), .A4(new_n836), .ZN(G311));
  INV_X1    g412(.A(G311), .ZN(G150));
  NAND2_X1  g413(.A1(new_n627), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n522), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n529), .A2(G55), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n532), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n566), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n846), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n840), .B(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n853), .A2(new_n854), .A3(G860), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n847), .A2(G860), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT104), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  OR2_X1    g433(.A1(new_n855), .A2(new_n858), .ZN(G145));
  NAND2_X1  g434(.A1(new_n483), .A2(G142), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT106), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n493), .A2(G130), .ZN(new_n862));
  OR2_X1    g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n863), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT107), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n639), .ZN(new_n867));
  INV_X1    g442(.A(new_n719), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n512), .A2(new_n514), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n504), .A2(new_n508), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n870), .A2(KEYINPUT105), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT105), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n801), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n775), .ZN(new_n878));
  INV_X1    g453(.A(new_n827), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n869), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n867), .B(new_n719), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT108), .ZN(new_n886));
  XNOR2_X1  g461(.A(G162), .B(new_n650), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G160), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(new_n889), .A3(new_n884), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n883), .B2(new_n884), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n892), .B2(new_n882), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g470(.A(G290), .B(G305), .Z(new_n896));
  XNOR2_X1  g471(.A(G303), .B(new_n600), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n627), .A2(new_n633), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n850), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n621), .A2(new_n581), .A3(new_n586), .A4(new_n625), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n621), .A2(new_n625), .B1(new_n581), .B2(new_n586), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT41), .B1(new_n904), .B2(new_n905), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n626), .A2(G299), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n903), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n906), .A2(KEYINPUT109), .A3(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n907), .B1(new_n915), .B2(new_n902), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT111), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(KEYINPUT111), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n900), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n900), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(G868), .B2(new_n846), .ZN(G295));
  OAI21_X1  g497(.A(new_n921), .B1(G868), .B2(new_n846), .ZN(G331));
  INV_X1    g498(.A(new_n898), .ZN(new_n924));
  NAND2_X1  g499(.A1(G168), .A2(G171), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n550), .A2(new_n554), .A3(G301), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n851), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n550), .A2(new_n554), .A3(G301), .ZN(new_n928));
  AOI21_X1  g503(.A(G301), .B1(new_n550), .B2(new_n554), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n850), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n913), .A3(new_n914), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n932), .A2(KEYINPUT112), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n931), .A2(new_n913), .A3(new_n914), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n927), .A2(new_n930), .A3(new_n906), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n924), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(KEYINPUT112), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n941), .A2(new_n898), .A3(new_n936), .A4(new_n935), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n908), .A2(new_n912), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n931), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n936), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n924), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n947), .A2(new_n942), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n943), .B(KEYINPUT44), .C1(new_n948), .C2(new_n939), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n938), .A2(new_n940), .A3(new_n942), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n942), .A3(new_n939), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI211_X1 g531(.A(KEYINPUT113), .B(KEYINPUT44), .C1(new_n952), .C2(new_n953), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n949), .B1(new_n956), .B2(new_n957), .ZN(G397));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n875), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n474), .A2(new_n478), .A3(G40), .A4(new_n481), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n801), .B(G2067), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT114), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n775), .B(G1996), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n868), .A2(new_n721), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n868), .A2(new_n721), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(G290), .B(G1986), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n964), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n503), .A2(new_n510), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n870), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n961), .A2(G1384), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AND4_X1   g554(.A1(G40), .A2(new_n474), .A3(new_n478), .A4(new_n481), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n871), .B1(new_n512), .B2(new_n514), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n961), .B1(new_n981), .B2(G1384), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n811), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT120), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n976), .B2(new_n870), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n981), .A2(G1384), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n963), .B1(new_n990), .B2(new_n988), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT117), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n989), .A2(new_n991), .A3(new_n789), .A4(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT120), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n983), .A2(new_n994), .A3(new_n811), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n985), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G8), .ZN(new_n997));
  INV_X1    g572(.A(G8), .ZN(new_n998));
  NOR2_X1   g573(.A1(G168), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(KEYINPUT51), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(G8), .C1(new_n996), .C2(G286), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT123), .B1(new_n996), .B2(new_n999), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n996), .A2(KEYINPUT123), .A3(new_n999), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1001), .B(new_n1003), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n963), .B1(new_n875), .B2(new_n978), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT115), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(new_n961), .C1(G164), .C2(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1008), .A2(new_n1012), .A3(new_n781), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n1014));
  INV_X1    g589(.A(G1961), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1013), .A2(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OR3_X1    g592(.A1(new_n983), .A2(new_n1014), .A3(G2078), .ZN(new_n1018));
  AOI21_X1  g593(.A(G301), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(G166), .B2(new_n998), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(G166), .A2(new_n1020), .A3(new_n998), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1022), .A2(KEYINPUT118), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n1025));
  NAND3_X1  g600(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(new_n1021), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1971), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n1029), .A2(new_n1030), .B1(G2090), .B2(new_n1016), .ZN(new_n1031));
  AOI211_X1 g606(.A(KEYINPUT116), .B(G1971), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1032));
  OAI211_X1 g607(.A(G8), .B(new_n1028), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n592), .A2(G651), .B1(new_n529), .B2(G49), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n544), .A2(KEYINPUT82), .A3(G87), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT82), .B1(new_n544), .B2(G87), .ZN(new_n1036));
  OAI211_X1 g611(.A(G1976), .B(new_n1034), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n870), .A2(new_n872), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n959), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1037), .B(G8), .C1(new_n963), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n600), .B2(G1976), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n998), .B1(new_n980), .B2(new_n990), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1044), .B2(new_n1037), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n609), .A2(new_n608), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(new_n606), .ZN(new_n1050));
  AND4_X1   g625(.A1(new_n1048), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G305), .A2(G1981), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1048), .A3(new_n606), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(KEYINPUT49), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1044), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1046), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n987), .A2(new_n988), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1060));
  AND4_X1   g635(.A1(new_n750), .A2(new_n1059), .A3(new_n1060), .A4(new_n980), .ZN(new_n1061));
  OAI21_X1  g636(.A(G8), .B1(new_n1029), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1057), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1033), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1007), .A2(new_n1019), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n996), .A2(G8), .A3(G168), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT63), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1069));
  INV_X1    g644(.A(G1971), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1061), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1058), .B1(new_n1071), .B2(new_n998), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1067), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1033), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1057), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1058), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT116), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1016), .A2(G2090), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1077), .B1(new_n1082), .B2(G8), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1067), .A2(new_n1075), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT63), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(G288), .A2(G1976), .ZN(new_n1086));
  XOR2_X1   g661(.A(new_n1086), .B(KEYINPUT119), .Z(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1044), .B1(new_n1088), .B2(new_n1051), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1076), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1008), .A2(new_n1012), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1059), .A2(new_n1060), .A3(new_n980), .ZN(new_n1093));
  INV_X1    g668(.A(G1956), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n581), .B2(new_n586), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n578), .A2(new_n574), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n586), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT121), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1092), .A2(new_n1101), .A3(new_n1095), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1105), .A2(KEYINPUT61), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1096), .A2(new_n1107), .A3(new_n1102), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT122), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  INV_X1    g686(.A(G1996), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1008), .A2(new_n1012), .A3(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT58), .B(G1341), .Z(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1039), .B2(new_n963), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1116), .B2(new_n567), .ZN(new_n1117));
  AOI211_X1 g692(.A(KEYINPUT59), .B(new_n566), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT61), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1104), .A2(new_n1106), .A3(new_n1122), .A4(new_n1108), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1016), .A2(new_n817), .ZN(new_n1124));
  OR3_X1    g699(.A1(new_n1039), .A2(new_n963), .A3(G2067), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT60), .A3(new_n627), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n626), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1128), .B(new_n1130), .C1(KEYINPUT60), .C2(new_n1127), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1110), .A2(new_n1121), .A3(new_n1123), .A4(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1104), .B(new_n1108), .C1(new_n626), .C2(new_n1127), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1105), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1016), .A2(new_n1015), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n962), .A2(KEYINPUT53), .A3(new_n781), .A4(new_n1008), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G171), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1136), .A2(G301), .A3(new_n1137), .A4(new_n1018), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1142), .A2(KEYINPUT54), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1144), .A3(G171), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1147));
  NOR2_X1   g722(.A1(new_n1139), .A2(G171), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(new_n1019), .ZN(new_n1149));
  AND4_X1   g724(.A1(new_n1146), .A2(new_n1149), .A3(new_n1006), .A4(new_n1064), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1090), .B1(new_n1135), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1066), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(KEYINPUT126), .B(new_n1090), .C1(new_n1135), .C2(new_n1150), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n975), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n969), .A2(new_n971), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n801), .A2(G2067), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n964), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n964), .A2(new_n1112), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT46), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n964), .B1(new_n775), .B2(new_n965), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G290), .A2(G1986), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n964), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT48), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n969), .A2(new_n972), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1158), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1158), .A2(KEYINPUT127), .A3(new_n1163), .A4(new_n1167), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1155), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g748(.A(new_n668), .ZN(new_n1175));
  NOR4_X1   g749(.A1(G229), .A2(new_n463), .A3(new_n1175), .A4(G227), .ZN(new_n1176));
  NAND3_X1  g750(.A1(new_n894), .A2(new_n954), .A3(new_n1176), .ZN(G225));
  INV_X1    g751(.A(G225), .ZN(G308));
endmodule


