//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  XNOR2_X1  g000(.A(G116), .B(G119), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT2), .B(G113), .Z(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(new_n187), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT66), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT0), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n194), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT68), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n198), .A2(new_n206), .A3(new_n201), .A4(new_n203), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G137), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(G134), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI211_X1 g031(.A(KEYINPUT69), .B(KEYINPUT11), .C1(new_n209), .C2(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n213), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(new_n212), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n216), .B1(new_n211), .B2(G137), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT69), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(new_n214), .A3(new_n216), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NOR3_X1   g044(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n231));
  OAI22_X1  g045(.A1(new_n230), .A2(new_n231), .B1(new_n199), .B2(new_n200), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n196), .A2(G143), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n194), .A2(KEYINPUT66), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n235), .A2(G143), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n195), .A2(new_n197), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT67), .B1(new_n242), .B2(new_n235), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n233), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n208), .A2(new_n228), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n226), .B1(new_n215), .B2(new_n212), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n225), .B2(new_n226), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n200), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n248));
  AOI21_X1  g062(.A(G146), .B1(new_n195), .B2(new_n197), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT67), .B1(new_n249), .B2(new_n239), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n234), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  AND4_X1   g067(.A1(new_n253), .A2(new_n198), .A3(G128), .A4(new_n203), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n247), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n245), .A2(KEYINPUT30), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n205), .A2(new_n207), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n232), .B1(new_n250), .B2(new_n251), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n254), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT66), .B(G143), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n240), .B1(new_n261), .B2(G146), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n243), .B1(KEYINPUT67), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n263), .B2(new_n248), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n228), .A2(new_n259), .B1(new_n264), .B2(new_n247), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n193), .B(new_n256), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G237), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G210), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n270), .B(KEYINPUT27), .Z(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G101), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g087(.A(new_n193), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n245), .A2(new_n274), .A3(new_n255), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n267), .A2(KEYINPUT31), .A3(new_n273), .A4(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(G472), .A2(G902), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n267), .A2(new_n273), .A3(new_n275), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n245), .A2(new_n274), .A3(new_n255), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n274), .B1(new_n245), .B2(new_n255), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT28), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n275), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n273), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n276), .B(new_n277), .C1(new_n280), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT28), .B1(new_n265), .B2(new_n274), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n245), .A2(new_n255), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n193), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n275), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n279), .B(new_n278), .C1(new_n293), .C2(new_n273), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n276), .A4(new_n277), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n283), .A2(KEYINPUT29), .A3(new_n273), .A4(new_n285), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n283), .A2(new_n273), .A3(new_n285), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n273), .B1(new_n267), .B2(new_n275), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n298), .B(new_n299), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n304), .A2(KEYINPUT70), .A3(G472), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT70), .B1(new_n304), .B2(G472), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n297), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  OAI21_X1  g122(.A(G125), .B1(new_n257), .B2(new_n258), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n310), .B(new_n260), .C1(new_n263), .C2(new_n248), .ZN(new_n311));
  INV_X1    g125(.A(G224), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G953), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT7), .A4(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G104), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(new_n316), .B2(G107), .ZN(new_n317));
  AOI21_X1  g131(.A(G101), .B1(new_n316), .B2(G107), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n319));
  INV_X1    g133(.A(G107), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G104), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G101), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(G104), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n316), .A2(G107), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n187), .A2(KEYINPUT5), .ZN(new_n329));
  INV_X1    g143(.A(G116), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n330), .A2(KEYINPUT5), .A3(G119), .ZN(new_n331));
  INV_X1    g145(.A(G113), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n329), .A2(new_n333), .B1(new_n191), .B2(new_n187), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n328), .A2(new_n334), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G122), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT8), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n315), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n309), .A2(new_n311), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT7), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n313), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT85), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(KEYINPUT85), .A3(new_n344), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n340), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n322), .B2(new_n326), .ZN(new_n351));
  INV_X1    g165(.A(new_n326), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(KEYINPUT78), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n354), .A3(new_n334), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT82), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n317), .A2(new_n321), .A3(new_n325), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n353), .A2(KEYINPUT4), .B1(new_n357), .B2(G101), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n357), .A2(KEYINPUT4), .A3(G101), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n193), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n351), .A2(new_n334), .A3(new_n354), .A4(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n356), .A2(new_n337), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n362), .A2(new_n360), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n366), .A2(KEYINPUT83), .A3(new_n337), .A4(new_n356), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n349), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT6), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n356), .A2(new_n360), .A3(new_n362), .ZN(new_n371));
  INV_X1    g185(.A(new_n337), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n355), .A2(KEYINPUT82), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n362), .A2(new_n360), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n370), .B(new_n372), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n371), .A2(KEYINPUT84), .A3(new_n370), .A4(new_n372), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n341), .B(new_n313), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n374), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G210), .B1(G237), .B2(G902), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n369), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n384), .B(KEYINPUT86), .Z(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n369), .B2(new_n383), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n308), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n316), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT90), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n268), .A2(new_n269), .A3(G214), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n394), .A2(KEYINPUT87), .A3(new_n195), .A4(new_n197), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n268), .A2(new_n269), .A3(G143), .A4(G214), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT87), .B1(new_n261), .B2(new_n394), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n393), .B1(new_n399), .B2(new_n226), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n268), .A2(new_n269), .A3(G214), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n401), .B1(new_n242), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n396), .A3(new_n395), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT90), .A3(G131), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n226), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G140), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G125), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n310), .A2(G140), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT88), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(KEYINPUT19), .A3(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(new_n235), .C1(KEYINPUT19), .C2(new_n411), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n409), .A2(new_n410), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT16), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n418), .B(G146), .C1(KEYINPUT16), .C2(new_n409), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n407), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n403), .A2(new_n422), .A3(new_n396), .A4(new_n395), .ZN(new_n423));
  NAND2_X1  g237(.A1(KEYINPUT18), .A2(G131), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(G146), .A3(new_n414), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n417), .A2(new_n235), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n392), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n423), .A2(new_n424), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n423), .A2(new_n424), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n431), .A2(new_n432), .B1(new_n427), .B2(new_n426), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n418), .B1(KEYINPUT16), .B2(new_n409), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n235), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n419), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n400), .A2(new_n405), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(KEYINPUT17), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT17), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n400), .A2(new_n439), .A3(new_n405), .A4(new_n406), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n433), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n430), .B1(new_n441), .B2(new_n392), .ZN(new_n442));
  NOR2_X1   g256(.A1(G475), .A2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT20), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n405), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT90), .B1(new_n404), .B2(G131), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT17), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n436), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n440), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n392), .A3(new_n429), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n421), .A2(new_n429), .ZN(new_n452));
  INV_X1    g266(.A(new_n392), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n443), .ZN(new_n457));
  AOI211_X1 g271(.A(new_n453), .B(new_n433), .C1(new_n438), .C2(new_n440), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n392), .B1(new_n450), .B2(new_n429), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n298), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT91), .B(G475), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n445), .A2(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n269), .A2(G952), .ZN(new_n463));
  INV_X1    g277(.A(G234), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(new_n268), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n298), .B(new_n269), .C1(G234), .C2(G237), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(G898), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G478), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT9), .B(G234), .ZN(new_n474));
  INV_X1    g288(.A(G217), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n474), .A2(new_n475), .A3(G953), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n261), .A2(G128), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n200), .A2(G143), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n211), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G116), .B(G122), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G107), .ZN(new_n482));
  INV_X1    g296(.A(new_n481), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n320), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT13), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n479), .B1(new_n478), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(KEYINPUT92), .A3(new_n486), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT92), .B1(new_n478), .B2(new_n486), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n485), .B1(new_n492), .B2(G134), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n478), .A2(new_n479), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G134), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n480), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(G116), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n481), .B1(new_n499), .B2(new_n320), .ZN(new_n500));
  OR3_X1    g314(.A1(new_n481), .A2(new_n499), .A3(new_n320), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n477), .B1(new_n493), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n485), .ZN(new_n504));
  INV_X1    g318(.A(new_n491), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n487), .B1(new_n505), .B2(new_n489), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n506), .B2(new_n211), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n476), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n473), .B1(new_n510), .B2(new_n298), .ZN(new_n511));
  AOI211_X1 g325(.A(G902), .B(new_n472), .C1(new_n503), .C2(new_n509), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n462), .A2(new_n470), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n390), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n475), .B1(G234), .B2(new_n298), .ZN(new_n516));
  INV_X1    g330(.A(G119), .ZN(new_n517));
  OR3_X1    g331(.A1(new_n517), .A2(KEYINPUT71), .A3(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(G128), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT71), .B1(new_n517), .B2(G128), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT24), .B(G110), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT23), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n517), .B2(G128), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n525), .A2(new_n526), .A3(new_n519), .ZN(new_n527));
  INV_X1    g341(.A(G110), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n419), .A3(new_n427), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n530), .A2(new_n419), .A3(new_n533), .A4(new_n427), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n527), .A2(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n527), .A2(KEYINPUT72), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(G110), .A3(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n436), .B(new_n538), .C1(new_n522), .C2(new_n521), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT74), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT22), .B(G137), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n535), .A2(new_n539), .A3(new_n544), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n516), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n547), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n544), .B1(new_n535), .B2(new_n539), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n298), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(KEYINPUT25), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n516), .A2(G902), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n546), .B2(new_n547), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G221), .B1(new_n474), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G469), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT81), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n269), .A2(G227), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT76), .ZN(new_n566));
  XNOR2_X1  g380(.A(G110), .B(G140), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT1), .B1(new_n261), .B2(G146), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n570), .A2(G128), .B1(new_n203), .B2(new_n198), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT77), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n260), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n198), .A2(new_n203), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n253), .B1(new_n242), .B2(new_n235), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n572), .B(new_n574), .C1(new_n575), .C2(new_n200), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n327), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n358), .A2(new_n359), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n351), .A2(KEYINPUT10), .A3(new_n354), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n259), .A2(new_n581), .B1(new_n264), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n228), .B(KEYINPUT79), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n228), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n580), .B2(new_n583), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n564), .B(new_n569), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT80), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n574), .B1(new_n575), .B2(new_n200), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n254), .B1(new_n591), .B2(KEYINPUT77), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n328), .B1(new_n592), .B2(new_n576), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n252), .A2(new_n254), .A3(new_n327), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n228), .B(new_n590), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n586), .B1(new_n578), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n568), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n588), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n264), .A2(new_n582), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n581), .A2(new_n208), .A3(new_n244), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n591), .A2(KEYINPUT77), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n260), .A3(new_n576), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT10), .B1(new_n607), .B2(new_n327), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n228), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n600), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n564), .B1(new_n610), .B2(new_n569), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n563), .B(new_n298), .C1(new_n602), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n599), .A2(new_n600), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n605), .A2(new_n608), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n569), .B1(new_n614), .B2(new_n584), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n613), .A2(new_n569), .B1(new_n615), .B2(new_n609), .ZN(new_n616));
  OAI21_X1  g430(.A(G469), .B1(new_n616), .B2(G902), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n562), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n307), .A2(new_n515), .A3(new_n560), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT93), .B(G101), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G3));
  NAND4_X1  g435(.A1(new_n369), .A2(KEYINPUT94), .A3(new_n383), .A4(new_n384), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(new_n308), .ZN(new_n623));
  INV_X1    g437(.A(new_n384), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n374), .A2(new_n381), .A3(new_n382), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT85), .B1(new_n341), .B2(new_n344), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n346), .B(new_n343), .C1(new_n309), .C2(new_n311), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n339), .B(new_n315), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n368), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n298), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n624), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT94), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n385), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT95), .B(G478), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n510), .B2(new_n298), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n510), .A2(KEYINPUT33), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n503), .B2(new_n509), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n471), .A2(G902), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n636), .B1(new_n462), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n460), .A2(new_n461), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n456), .B1(new_n455), .B2(new_n443), .ZN(new_n647));
  AOI211_X1 g461(.A(KEYINPUT20), .B(new_n444), .C1(new_n451), .C2(new_n454), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n643), .B1(new_n639), .B2(new_n641), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n503), .A2(new_n509), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(G902), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n650), .B1(new_n652), .B2(new_n637), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n649), .A2(KEYINPUT96), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n635), .A2(new_n655), .A3(new_n470), .ZN(new_n656));
  INV_X1    g470(.A(new_n560), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n298), .B(new_n276), .C1(new_n280), .C2(new_n286), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(G472), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n287), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n618), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n445), .A2(new_n666), .A3(new_n457), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n647), .A2(KEYINPUT97), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n472), .B1(new_n651), .B2(G902), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n510), .A2(new_n298), .A3(new_n473), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n460), .A2(new_n461), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n667), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n470), .A2(new_n672), .A3(new_n633), .A4(new_n623), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n618), .A3(new_n661), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NOR2_X1   g490(.A1(new_n544), .A2(KEYINPUT36), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n540), .B(new_n677), .Z(new_n678));
  OAI22_X1  g492(.A1(new_n550), .A2(new_n554), .B1(new_n557), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n659), .A2(new_n287), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT98), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT98), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n659), .A2(new_n679), .A3(new_n682), .A4(new_n287), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n646), .B(new_n513), .C1(new_n647), .C2(new_n648), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n469), .ZN(new_n686));
  INV_X1    g500(.A(new_n308), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n387), .B1(new_n625), .B2(new_n630), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n687), .B1(new_n688), .B2(new_n385), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n618), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  INV_X1    g507(.A(new_n679), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT70), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n299), .A2(new_n298), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT29), .B1(new_n293), .B2(new_n273), .ZN(new_n697));
  INV_X1    g511(.A(new_n303), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(G472), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n304), .A2(KEYINPUT70), .A3(G472), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n694), .B1(new_n703), .B2(new_n297), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n466), .B1(new_n467), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n667), .A2(new_n671), .A3(new_n668), .A4(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT99), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n704), .A2(new_n710), .A3(new_n618), .A4(new_n635), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G128), .ZN(G30));
  NOR2_X1   g526(.A1(new_n386), .A2(new_n389), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT38), .ZN(new_n714));
  INV_X1    g528(.A(new_n513), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n649), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n714), .A2(new_n687), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n273), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n267), .B2(new_n275), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n298), .B1(new_n292), .B2(new_n273), .ZN(new_n720));
  OAI21_X1  g534(.A(G472), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n679), .B1(new_n297), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n706), .B(KEYINPUT39), .Z(new_n724));
  NAND2_X1  g538(.A1(new_n618), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT100), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT40), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n723), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n242), .ZN(G45));
  NOR3_X1   g545(.A1(new_n462), .A2(new_n644), .A3(new_n706), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n704), .A2(new_n618), .A3(new_n635), .A4(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT101), .B(G146), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G48));
  OAI21_X1  g549(.A(new_n298), .B1(new_n602), .B2(new_n611), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n563), .A2(KEYINPUT102), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI221_X1 g552(.A(new_n298), .B1(KEYINPUT102), .B2(new_n563), .C1(new_n602), .C2(new_n611), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n561), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n307), .A3(new_n560), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n656), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT41), .B(G113), .Z(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G15));
  NAND4_X1  g559(.A1(new_n673), .A2(new_n307), .A3(new_n560), .A4(new_n741), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G116), .ZN(G18));
  NOR2_X1   g561(.A1(new_n740), .A2(new_n634), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n307), .A3(new_n686), .A4(new_n679), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NAND3_X1  g564(.A1(new_n649), .A2(new_n470), .A3(new_n715), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n657), .A2(new_n660), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  INV_X1    g568(.A(KEYINPUT103), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n680), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n659), .A2(new_n679), .A3(KEYINPUT103), .A4(new_n287), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n748), .A2(new_n732), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT104), .B(G125), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G27));
  NAND3_X1  g574(.A1(new_n688), .A2(new_n308), .A3(new_n385), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n688), .A2(KEYINPUT105), .A3(new_n308), .A4(new_n385), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n618), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n763), .A2(new_n618), .A3(KEYINPUT106), .A4(new_n764), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n701), .A2(new_n702), .B1(new_n288), .B2(new_n296), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT107), .B1(new_n770), .B2(new_n657), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n307), .A2(new_n772), .A3(new_n560), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n769), .A2(new_n732), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n307), .A2(new_n560), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n767), .B2(new_n768), .ZN(new_n776));
  INV_X1    g590(.A(new_n732), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT42), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n774), .A2(KEYINPUT42), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n710), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  NAND2_X1  g596(.A1(new_n763), .A2(new_n764), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n660), .A2(new_n679), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT110), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n644), .B1(new_n649), .B2(KEYINPUT109), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(KEYINPUT43), .C1(KEYINPUT109), .C2(new_n649), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT43), .B1(new_n462), .B2(new_n653), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT108), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n783), .B1(new_n790), .B2(KEYINPUT44), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n616), .A2(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n616), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(G469), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(G469), .A2(G902), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT46), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n612), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n795), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n562), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n724), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n791), .B(new_n802), .C1(KEYINPUT44), .C2(new_n790), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  XNOR2_X1  g618(.A(new_n800), .B(KEYINPUT47), .ZN(new_n805));
  INV_X1    g619(.A(new_n783), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n307), .A2(new_n777), .A3(new_n560), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT111), .B(G140), .Z(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(G42));
  INV_X1    g624(.A(new_n714), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n297), .A2(new_n560), .A3(new_n721), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n811), .A2(new_n562), .A3(new_n687), .A4(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n786), .B1(KEYINPUT109), .B2(new_n649), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n738), .A2(new_n739), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n813), .B(new_n818), .C1(new_n817), .C2(new_n816), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n756), .A2(new_n732), .A3(new_n757), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n307), .A2(new_n618), .A3(new_n679), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n667), .A2(new_n668), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n646), .A2(new_n513), .A3(new_n707), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n783), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n769), .A2(new_n821), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(new_n781), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n746), .A2(new_n749), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n390), .A2(new_n469), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n462), .A2(new_n653), .ZN(new_n830));
  INV_X1    g644(.A(new_n685), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n661), .A2(new_n829), .A3(new_n832), .A4(new_n618), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n691), .A2(new_n833), .A3(new_n619), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n753), .B1(new_n742), .B2(new_n656), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n828), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n827), .A2(new_n779), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n634), .A2(new_n716), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n618), .A3(new_n707), .A4(new_n722), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n711), .A2(new_n733), .A3(new_n839), .A4(new_n758), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n822), .B(new_n635), .C1(new_n710), .C2(new_n732), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n758), .A4(new_n839), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n820), .B1(new_n837), .B2(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n837), .A2(new_n820), .A3(new_n845), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(KEYINPUT112), .ZN(new_n848));
  INV_X1    g662(.A(new_n769), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n771), .A2(new_n732), .A3(new_n773), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT42), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n776), .A2(new_n778), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n746), .A2(new_n749), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n691), .A2(new_n833), .A3(new_n619), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n635), .A2(new_n655), .A3(new_n470), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n770), .A2(new_n657), .A3(new_n740), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n856), .A2(new_n857), .B1(new_n748), .B2(new_n752), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n841), .A2(new_n844), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT53), .A4(new_n827), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT54), .B1(new_n848), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n854), .A2(new_n866), .A3(new_n858), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT113), .B1(new_n828), .B2(new_n835), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n834), .A2(new_n820), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n861), .A3(new_n779), .A4(new_n827), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n846), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n815), .A2(new_n561), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n805), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n789), .A2(new_n787), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n466), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n657), .A3(new_n660), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n877), .A2(new_n880), .A3(new_n806), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n811), .A2(new_n308), .A3(new_n740), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT50), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(KEYINPUT50), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n806), .A2(new_n741), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n756), .A3(new_n757), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n812), .A2(new_n465), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n806), .A3(KEYINPUT115), .A4(new_n741), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n462), .A3(new_n644), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n880), .A2(new_n882), .A3(new_n886), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n888), .A2(new_n891), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n875), .B1(new_n881), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n771), .A2(new_n773), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n890), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT48), .Z(new_n903));
  NAND3_X1  g717(.A1(new_n895), .A2(new_n655), .A3(new_n896), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n880), .A2(KEYINPUT116), .A3(new_n748), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT116), .B1(new_n880), .B2(new_n748), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n463), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n881), .A2(new_n899), .A3(new_n875), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n874), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(G952), .A2(G953), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n819), .B1(new_n911), .B2(new_n912), .ZN(G75));
  NOR2_X1   g727(.A1(new_n269), .A2(G952), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n374), .A2(new_n381), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n382), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT55), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n826), .A2(new_n781), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n853), .A2(new_n918), .A3(new_n859), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n919), .B2(new_n861), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n851), .A2(new_n826), .A3(new_n852), .A4(new_n781), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n845), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n298), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(G210), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n917), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n387), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n917), .A2(new_n927), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n914), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(G51));
  OAI21_X1  g745(.A(KEYINPUT54), .B1(new_n920), .B2(new_n923), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n873), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n795), .B(KEYINPUT57), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n934), .A2(new_n935), .B1(new_n611), .B2(new_n602), .ZN(new_n936));
  OR3_X1    g750(.A1(new_n924), .A2(new_n298), .A3(new_n794), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n914), .B1(new_n936), .B2(new_n937), .ZN(G54));
  NAND4_X1  g752(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .A4(new_n455), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT117), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(KEYINPUT117), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n925), .A2(KEYINPUT58), .A3(G475), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n914), .B1(new_n942), .B2(new_n442), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(G60));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n945));
  INV_X1    g759(.A(new_n914), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n642), .B(KEYINPUT118), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(G478), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT59), .Z(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT119), .B1(new_n933), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n953));
  INV_X1    g767(.A(new_n951), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n953), .B(new_n954), .C1(new_n932), .C2(new_n873), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n946), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n950), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n947), .B1(new_n874), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n945), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n873), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n872), .B1(new_n871), .B2(new_n846), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n951), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n953), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n933), .A2(KEYINPUT119), .A3(new_n951), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n847), .A2(KEYINPUT112), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n862), .A2(new_n863), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n967), .A3(new_n846), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n960), .B1(new_n968), .B2(KEYINPUT54), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n948), .B1(new_n969), .B2(new_n950), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n965), .A2(new_n970), .A3(KEYINPUT120), .A4(new_n946), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n959), .A2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT121), .Z(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n924), .A2(new_n678), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n546), .A2(new_n547), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n924), .A2(new_n975), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n976), .B(new_n946), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G66));
  OAI21_X1  g795(.A(G953), .B1(new_n468), .B2(new_n312), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n836), .B2(G953), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n915), .B1(G898), .B2(new_n269), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G69));
  NAND2_X1  g799(.A1(new_n779), .A2(new_n781), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT124), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n803), .A2(new_n808), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n901), .A2(new_n838), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n758), .B(new_n842), .C1(new_n989), .C2(new_n801), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n269), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n256), .B1(new_n265), .B2(new_n266), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n415), .B1(KEYINPUT19), .B2(new_n411), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n993), .B(new_n994), .Z(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(G900), .B2(G953), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n988), .ZN(new_n998));
  INV_X1    g812(.A(new_n730), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n842), .A2(new_n758), .ZN(new_n1000));
  OR3_X1    g814(.A1(new_n999), .A2(KEYINPUT62), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT62), .B1(new_n999), .B2(new_n1000), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n832), .B(KEYINPUT122), .ZN(new_n1003));
  INV_X1    g817(.A(new_n775), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n726), .A2(new_n1003), .A3(new_n1004), .A4(new_n806), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n269), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n995), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT123), .Z(new_n1010));
  NAND3_X1  g824(.A1(new_n997), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n997), .A2(KEYINPUT125), .A3(new_n1008), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1009), .B1(new_n997), .B2(KEYINPUT125), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(G72));
  XNOR2_X1  g828(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n700), .A2(new_n298), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1015), .B(new_n1016), .Z(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(new_n1006), .B2(new_n859), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n914), .B1(new_n1019), .B2(new_n719), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1017), .B1(new_n991), .B2(new_n836), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n267), .A2(new_n718), .A3(new_n275), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1017), .B1(new_n698), .B2(new_n278), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT127), .Z(new_n1025));
  AOI21_X1  g839(.A(new_n1023), .B1(new_n968), .B2(new_n1025), .ZN(G57));
endmodule


