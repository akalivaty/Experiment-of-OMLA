//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT68), .A3(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT2), .B(G113), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n189), .A2(new_n191), .B1(G116), .B2(new_n188), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n193), .B2(KEYINPUT5), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT5), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n202), .A2(new_n188), .A3(KEYINPUT87), .A4(G116), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(G113), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n197), .B1(new_n199), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT82), .B(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n207), .A2(KEYINPUT3), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g028(.A(KEYINPUT81), .B(KEYINPUT3), .C1(new_n207), .C2(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n211), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n209), .A2(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(G107), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n206), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(KEYINPUT4), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n211), .A2(new_n216), .A3(KEYINPUT83), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT83), .B1(new_n211), .B2(new_n216), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n224), .B1(new_n227), .B2(G101), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n211), .A2(new_n216), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n211), .A2(new_n216), .A3(KEYINPUT83), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n196), .B1(new_n194), .B2(new_n235), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n198), .A2(KEYINPUT67), .A3(new_n195), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n223), .B1(new_n228), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n223), .B(new_n241), .C1(new_n228), .C2(new_n239), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(KEYINPUT6), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT64), .A2(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT64), .A2(G143), .ZN(new_n250));
  AOI21_X1  g064(.A(G146), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  INV_X1    g066(.A(G146), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT65), .A3(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n248), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n249), .A2(G146), .A3(new_n250), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n253), .A2(G143), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n246), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT88), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n255), .A2(G146), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n266));
  OAI21_X1  g080(.A(G128), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n251), .B2(new_n257), .ZN(new_n268));
  INV_X1    g082(.A(G125), .ZN(new_n269));
  INV_X1    g083(.A(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n259), .A2(new_n260), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT88), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n262), .A2(new_n274), .A3(G125), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n264), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT89), .B(G224), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n240), .A2(new_n280), .A3(new_n242), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n245), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n218), .A2(new_n221), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n206), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n241), .B(KEYINPUT8), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n199), .A2(KEYINPUT90), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n204), .B1(new_n199), .B2(KEYINPUT90), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n197), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n284), .B(new_n285), .C1(new_n288), .C2(new_n283), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n278), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n264), .A2(new_n273), .A3(new_n275), .A4(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n263), .B2(new_n273), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(KEYINPUT91), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT91), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n295), .B(new_n291), .C1(new_n263), .C2(new_n273), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n289), .B(new_n292), .C1(new_n294), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n298), .B2(new_n244), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n282), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT92), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n282), .A2(new_n299), .A3(KEYINPUT92), .ZN(new_n303));
  OAI21_X1  g117(.A(G210), .B1(G237), .B2(G902), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT93), .Z(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n282), .A2(new_n299), .A3(new_n304), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT94), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n305), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n300), .B2(new_n301), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n307), .B1(new_n314), .B2(new_n303), .ZN(new_n315));
  INV_X1    g129(.A(new_n311), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT94), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G221), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT9), .B(G234), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n268), .A2(new_n272), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT10), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n325), .A2(new_n283), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n259), .A2(new_n260), .A3(new_n271), .ZN(new_n329));
  AND2_X1   g143(.A1(KEYINPUT64), .A2(G143), .ZN(new_n330));
  NOR2_X1   g144(.A1(KEYINPUT64), .A2(G143), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n265), .B1(new_n332), .B2(G146), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G128), .B1(new_n251), .B2(new_n266), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n328), .B1(new_n336), .B2(new_n283), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n253), .B1(new_n330), .B2(new_n331), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n270), .B1(new_n338), .B2(KEYINPUT1), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n272), .B1(new_n339), .B2(new_n333), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n340), .A2(KEYINPUT85), .A3(new_n218), .A4(new_n221), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n327), .B1(new_n342), .B2(new_n326), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT11), .ZN(new_n344));
  INV_X1    g158(.A(G134), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(G137), .ZN(new_n346));
  INV_X1    g160(.A(G137), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT11), .A3(G134), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(G137), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G131), .ZN(new_n351));
  INV_X1    g165(.A(G131), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n346), .A2(new_n348), .A3(new_n352), .A4(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n338), .A2(new_n254), .A3(new_n256), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n356), .A2(new_n248), .B1(new_n333), .B2(new_n246), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n234), .A2(new_n357), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n228), .A2(new_n358), .A3(KEYINPUT84), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n262), .B1(new_n227), .B2(new_n233), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n231), .A2(G101), .A3(new_n232), .ZN(new_n362));
  INV_X1    g176(.A(new_n224), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n343), .B(new_n355), .C1(new_n359), .C2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G110), .B(G140), .ZN(new_n367));
  INV_X1    g181(.A(G953), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n368), .A2(G227), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n367), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n343), .B1(new_n359), .B2(new_n365), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n354), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n324), .B1(new_n218), .B2(new_n221), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT85), .B1(new_n222), .B2(new_n340), .ZN(new_n377));
  INV_X1    g191(.A(new_n341), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT12), .A3(new_n354), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT12), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n375), .B1(new_n337), .B2(new_n341), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(new_n355), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n366), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n372), .A2(new_n374), .B1(new_n385), .B2(new_n370), .ZN(new_n386));
  OAI21_X1  g200(.A(G469), .B1(new_n386), .B2(G902), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT84), .B1(new_n228), .B2(new_n358), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n361), .A2(new_n360), .A3(new_n364), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n390), .A2(new_n355), .A3(new_n343), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n355), .B1(new_n390), .B2(new_n343), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n370), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n366), .A2(new_n384), .A3(new_n371), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XOR2_X1   g209(.A(KEYINPUT86), .B(G469), .Z(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n322), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n323), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n368), .A3(G214), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n249), .A3(new_n250), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n400), .A2(new_n368), .A3(G143), .A4(G214), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n352), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G125), .B(G140), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(new_n253), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n402), .A2(new_n403), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n406), .A2(new_n352), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n207), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT96), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n269), .A2(KEYINPUT16), .A3(G140), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G140), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G125), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n269), .A2(G140), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT16), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n419), .A2(KEYINPUT75), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT76), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(G146), .ZN(new_n429));
  INV_X1    g243(.A(new_n426), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n419), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n430), .B(G146), .C1(new_n431), .C2(new_n418), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT76), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n253), .B1(new_n425), .B2(new_n426), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n402), .A2(new_n352), .A3(new_n403), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n436), .B1(new_n438), .B2(new_n404), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n405), .A2(KEYINPUT17), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n414), .B(new_n417), .C1(new_n435), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n440), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n444), .A2(new_n433), .A3(new_n434), .A4(new_n429), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n416), .B1(new_n445), .B2(new_n414), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n322), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT97), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n449), .B(new_n322), .C1(new_n443), .C2(new_n446), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(G475), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n321), .A2(G217), .A3(new_n368), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n190), .A2(G122), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n190), .A2(G122), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(new_n209), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n249), .A2(G128), .A3(new_n250), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n270), .A2(G143), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(KEYINPUT13), .A3(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n462), .B(G134), .C1(KEYINPUT13), .C2(new_n460), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n345), .A3(new_n461), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n458), .A2(new_n209), .ZN(new_n467));
  INV_X1    g281(.A(new_n464), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n345), .B1(new_n460), .B2(new_n461), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT99), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT98), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n457), .A2(new_n472), .A3(KEYINPUT14), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n456), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n457), .B2(KEYINPUT14), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n457), .A2(KEYINPUT14), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n457), .A2(KEYINPUT14), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT98), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(KEYINPUT99), .A3(new_n456), .A4(new_n473), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n470), .B1(G107), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n455), .B1(new_n466), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n455), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n481), .A2(G107), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n465), .B(new_n484), .C1(new_n485), .C2(new_n470), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n454), .B1(new_n487), .B2(new_n322), .ZN(new_n488));
  AOI211_X1 g302(.A(G902), .B(new_n453), .C1(new_n483), .C2(new_n486), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n413), .B1(new_n491), .B2(new_n444), .ZN(new_n492));
  INV_X1    g306(.A(new_n416), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n408), .A2(KEYINPUT95), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT19), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n408), .A2(KEYINPUT95), .A3(KEYINPUT19), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n253), .A2(new_n498), .B1(new_n405), .B2(new_n437), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n432), .A2(KEYINPUT77), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT77), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n427), .A2(new_n501), .A3(G146), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n414), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n492), .A2(new_n417), .B1(new_n493), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(G475), .A2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT20), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n493), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n442), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT20), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n506), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(G234), .A2(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(G952), .A3(new_n368), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT21), .B(G898), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(G902), .A3(G953), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT100), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n451), .A2(new_n490), .A3(new_n513), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT101), .ZN(new_n522));
  INV_X1    g336(.A(G475), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n447), .B2(KEYINPUT97), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n524), .A2(new_n450), .B1(new_n508), .B2(new_n512), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT101), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n490), .A4(new_n520), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n399), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(G472), .A2(G902), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n354), .A2(new_n258), .A3(new_n261), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n345), .A2(G137), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n347), .A2(G134), .ZN(new_n535));
  OAI21_X1  g349(.A(G131), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n353), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n268), .B2(new_n272), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT66), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n353), .A2(new_n536), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n270), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n254), .A2(new_n256), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n338), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n539), .B(new_n541), .C1(new_n544), .C2(new_n329), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n532), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n357), .A2(new_n354), .B1(new_n324), .B2(new_n541), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT69), .B1(new_n548), .B2(KEYINPUT30), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n541), .B1(new_n544), .B2(new_n329), .ZN(new_n550));
  AND4_X1   g364(.A1(KEYINPUT69), .A2(new_n550), .A3(new_n533), .A4(KEYINPUT30), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n547), .B(new_n238), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n236), .A2(new_n237), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n550), .A3(new_n533), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n400), .A2(new_n368), .A3(G210), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT27), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT26), .B(G101), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n552), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT31), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n552), .A2(KEYINPUT31), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n238), .B1(new_n540), .B2(new_n546), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n548), .A2(KEYINPUT28), .A3(new_n553), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n554), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n560), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n531), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n567), .A2(new_n570), .A3(new_n568), .A4(new_n559), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT69), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n550), .A2(new_n533), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n578), .B2(new_n532), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n548), .A2(KEYINPUT69), .A3(KEYINPUT30), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n550), .A2(KEYINPUT66), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n545), .A3(new_n533), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n579), .A2(new_n580), .B1(new_n582), .B2(new_n532), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n555), .B1(new_n583), .B2(new_n238), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n576), .B1(new_n584), .B2(new_n559), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT71), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n548), .A2(new_n553), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n586), .B(KEYINPUT28), .C1(new_n587), .C2(new_n555), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n578), .A2(new_n238), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n569), .B1(new_n589), .B2(new_n554), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n570), .A2(KEYINPUT71), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n560), .A2(new_n575), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n573), .A2(KEYINPUT32), .B1(G472), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT70), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n573), .B2(KEYINPUT32), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n552), .A2(KEYINPUT31), .A3(new_n561), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT31), .B1(new_n552), .B2(new_n561), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n572), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n530), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT32), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(KEYINPUT70), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n596), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT80), .ZN(new_n606));
  OR3_X1    g420(.A1(new_n188), .A2(KEYINPUT73), .A3(G128), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT73), .B1(new_n188), .B2(G128), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n188), .A2(G128), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT24), .B(G110), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT74), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n188), .B2(G128), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n614), .A2(KEYINPUT23), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(KEYINPUT23), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n615), .A2(new_n609), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G110), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n435), .A2(new_n612), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n618), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n610), .A2(new_n611), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n621), .A2(new_n622), .B1(new_n253), .B2(new_n408), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n500), .A3(new_n502), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT22), .B(G137), .ZN(new_n626));
  INV_X1    g440(.A(G234), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n319), .A2(new_n627), .A3(G953), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n626), .B(new_n628), .Z(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n620), .A2(new_n624), .A3(new_n629), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n322), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n634), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n631), .A2(new_n322), .A3(new_n632), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G217), .B1(new_n627), .B2(G902), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT72), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(G902), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n631), .A2(new_n632), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT79), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n605), .A2(new_n606), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n606), .B1(new_n605), .B2(new_n647), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n318), .B(new_n529), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G101), .ZN(G3));
  NAND2_X1  g465(.A1(new_n601), .A2(new_n322), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G472), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n602), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n646), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n399), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n452), .A2(new_n322), .ZN(new_n658));
  INV_X1    g472(.A(new_n487), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(G902), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n658), .B1(new_n660), .B2(new_n452), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n487), .A2(KEYINPUT33), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n487), .A2(KEYINPUT33), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(G478), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n525), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n520), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n304), .B1(new_n282), .B2(new_n299), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n311), .B1(new_n307), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n657), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT102), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n511), .B1(new_n510), .B2(new_n506), .ZN(new_n676));
  AOI211_X1 g490(.A(KEYINPUT20), .B(new_n507), .C1(new_n509), .C2(new_n442), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n508), .A2(KEYINPUT103), .A3(new_n512), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n490), .B1(new_n524), .B2(new_n450), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n520), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n683));
  INV_X1    g497(.A(new_n669), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n680), .A2(new_n681), .A3(new_n685), .A4(new_n520), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n657), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT35), .B(G107), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G9));
  NOR2_X1   g504(.A1(new_n630), .A2(KEYINPUT36), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT105), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n625), .B(new_n692), .Z(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n639), .A2(new_n641), .B1(new_n694), .B2(new_n643), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n654), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n318), .A2(new_n529), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT37), .B(G110), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  OR2_X1    g513(.A1(new_n518), .A2(G900), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n515), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n680), .A2(new_n681), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT106), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n669), .A2(new_n695), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n703), .A2(new_n399), .A3(new_n704), .A4(new_n605), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  XNOR2_X1  g520(.A(new_n701), .B(KEYINPUT39), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n399), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT40), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n573), .A2(KEYINPUT32), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n587), .A2(new_n555), .A3(new_n559), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n711), .B(new_n713), .C1(new_n584), .C2(new_n560), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n560), .B1(new_n552), .B2(new_n554), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT108), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n716), .A3(new_n322), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G472), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n598), .A2(new_n710), .A3(new_n604), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n695), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n451), .A2(new_n513), .ZN(new_n721));
  INV_X1    g535(.A(new_n490), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n720), .A2(new_n316), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n315), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n709), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(new_n332), .Z(G45));
  NAND4_X1  g542(.A1(new_n721), .A2(new_n664), .A3(new_n661), .A4(new_n701), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n399), .A2(new_n605), .A3(new_n704), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  INV_X1    g546(.A(new_n323), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n371), .B1(new_n374), .B2(new_n366), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n366), .A2(new_n384), .A3(new_n371), .ZN(new_n735));
  OAI211_X1 g549(.A(KEYINPUT109), .B(new_n322), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT109), .B1(new_n395), .B2(new_n322), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n733), .B(new_n398), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT110), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n322), .B1(new_n734), .B2(new_n735), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(G469), .A3(new_n736), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n745), .A3(new_n733), .A4(new_n398), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT70), .B1(new_n602), .B2(new_n603), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n597), .B(KEYINPUT32), .C1(new_n601), .C2(new_n530), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n646), .B1(new_n749), .B2(new_n596), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n740), .A2(new_n746), .A3(new_n750), .A4(new_n670), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT41), .B(G113), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT111), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n751), .B(new_n753), .ZN(G15));
  NAND4_X1  g568(.A1(new_n740), .A2(new_n687), .A3(new_n746), .A4(new_n750), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G116), .ZN(G18));
  INV_X1    g570(.A(new_n695), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n605), .A2(new_n528), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n740), .A3(new_n684), .A4(new_n746), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NOR2_X1   g574(.A1(new_n669), .A2(new_n723), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(new_n520), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n566), .B1(new_n559), .B2(new_n592), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n530), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n653), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n646), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n740), .A2(new_n762), .A3(new_n746), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  NOR3_X1   g582(.A1(new_n765), .A2(new_n729), .A3(new_n695), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n740), .A2(new_n746), .A3(new_n684), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  OAI21_X1  g585(.A(new_n596), .B1(KEYINPUT32), .B2(new_n573), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n647), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(G469), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n385), .A2(new_n370), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n374), .A2(new_n366), .A3(new_n371), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n775), .B1(new_n778), .B2(new_n322), .ZN(new_n779));
  AOI211_X1 g593(.A(G902), .B(new_n396), .C1(new_n393), .C2(new_n394), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n733), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n306), .A2(new_n311), .A3(new_n308), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n774), .A2(KEYINPUT42), .A3(new_n730), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n316), .B(new_n307), .C1(new_n314), .C2(new_n303), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n399), .A3(new_n605), .A4(new_n647), .ZN(new_n787));
  OAI211_X1 g601(.A(KEYINPUT112), .B(new_n785), .C1(new_n787), .C2(new_n729), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n783), .A2(new_n750), .A3(new_n730), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT112), .B1(new_n790), .B2(new_n785), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n784), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  INV_X1    g607(.A(new_n703), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n787), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n345), .ZN(G36));
  NOR2_X1   g610(.A1(new_n775), .A2(new_n322), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n778), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT113), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n775), .B1(new_n778), .B2(new_n798), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n398), .B1(new_n802), .B2(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n733), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n721), .A2(new_n665), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT43), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n654), .A3(new_n757), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n782), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  INV_X1    g625(.A(new_n707), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n805), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n347), .ZN(G39));
  XNOR2_X1  g628(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n805), .B(new_n816), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n605), .A2(new_n782), .A3(new_n647), .A4(new_n729), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  AND2_X1   g634(.A1(new_n744), .A2(new_n398), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT49), .Z(new_n822));
  NAND4_X1  g636(.A1(new_n647), .A2(new_n311), .A3(new_n733), .A4(new_n806), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT115), .Z(new_n824));
  OR4_X1    g638(.A1(new_n719), .A2(new_n822), .A3(new_n726), .A4(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n767), .A2(new_n751), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n755), .A4(new_n759), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n759), .A2(new_n755), .A3(new_n767), .A4(new_n751), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT119), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n765), .A2(new_n695), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n605), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n490), .A2(new_n701), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n757), .A2(new_n451), .A3(new_n680), .A4(new_n836), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n834), .A2(new_n729), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n795), .B1(new_n783), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n792), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n701), .B(KEYINPUT117), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n399), .A2(new_n761), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT118), .B1(new_n843), .B2(new_n720), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n710), .A2(new_n718), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n757), .B1(new_n749), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n847));
  INV_X1    g661(.A(new_n842), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n323), .B(new_n848), .C1(new_n387), .C2(new_n398), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n847), .A3(new_n849), .A4(new_n761), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n844), .A2(new_n850), .A3(new_n731), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n770), .A2(new_n705), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT52), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n844), .A2(new_n850), .A3(new_n731), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n770), .A2(new_n705), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n667), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n860));
  AOI211_X1 g674(.A(KEYINPUT94), .B(new_n316), .C1(new_n306), .C2(new_n308), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT116), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n318), .A2(new_n864), .A3(new_n859), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n656), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n525), .A2(new_n722), .A3(new_n520), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n657), .A2(new_n318), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n650), .A2(new_n697), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n866), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n832), .A2(new_n841), .A3(new_n858), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n866), .A2(new_n869), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n751), .A2(new_n759), .A3(new_n755), .A4(new_n767), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n792), .A3(new_n839), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT52), .B1(new_n851), .B2(new_n852), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n855), .A2(new_n856), .A3(new_n854), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n870), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n872), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n650), .A2(new_n697), .A3(new_n868), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n864), .B1(new_n318), .B2(new_n859), .ZN(new_n883));
  AOI211_X1 g697(.A(KEYINPUT116), .B(new_n667), .C1(new_n312), .C2(new_n317), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n657), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n874), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n840), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT53), .B1(new_n887), .B2(new_n858), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n875), .A2(new_n878), .A3(new_n870), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n881), .B1(new_n890), .B2(new_n880), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n740), .A2(new_n746), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n786), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT43), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n806), .B(new_n894), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n895), .A2(KEYINPUT120), .A3(new_n515), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT120), .B1(new_n895), .B2(new_n515), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n719), .A2(new_n515), .A3(new_n646), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n525), .A2(new_n665), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n899), .A2(new_n834), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n646), .B(new_n765), .C1(new_n896), .C2(new_n897), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n726), .A2(new_n311), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n892), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT50), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n821), .A2(new_n323), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n786), .B(new_n904), .C1(new_n817), .C2(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n910), .A2(new_n913), .A3(KEYINPUT51), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT51), .B1(new_n910), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n899), .A2(new_n773), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT48), .Z(new_n917));
  NAND3_X1  g731(.A1(new_n904), .A2(new_n684), .A3(new_n892), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT121), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n901), .A2(new_n525), .A3(new_n665), .ZN(new_n920));
  INV_X1    g734(.A(G952), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(G953), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  NOR4_X1   g737(.A1(new_n891), .A2(new_n914), .A3(new_n915), .A4(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(G952), .A2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n825), .B1(new_n924), .B2(new_n925), .ZN(G75));
  NAND2_X1  g740(.A1(new_n921), .A2(G953), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT123), .Z(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT124), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n872), .A2(new_n879), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(G902), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n313), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n245), .A2(new_n281), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n279), .ZN(new_n934));
  XOR2_X1   g748(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n929), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n930), .A2(G210), .A3(G902), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n940), .B2(new_n937), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(G51));
  INV_X1    g756(.A(new_n928), .ZN(new_n943));
  AND4_X1   g757(.A1(G902), .A2(new_n930), .A3(new_n800), .A4(new_n801), .ZN(new_n944));
  INV_X1    g758(.A(new_n395), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n792), .A4(new_n839), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n946), .A2(new_n878), .A3(new_n831), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT54), .B1(new_n888), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n881), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n797), .B(KEYINPUT57), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n944), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n950), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n948), .B2(new_n881), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT125), .B1(new_n955), .B2(new_n945), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n943), .B1(new_n953), .B2(new_n956), .ZN(G54));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n931), .A2(new_n510), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n510), .B1(new_n931), .B2(new_n958), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n943), .B1(new_n959), .B2(new_n960), .ZN(G60));
  NAND2_X1  g775(.A1(new_n662), .A2(new_n663), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n658), .B(KEYINPUT59), .Z(new_n963));
  NAND3_X1  g777(.A1(new_n949), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n929), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n891), .B2(new_n963), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(G63));
  XNOR2_X1  g781(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n631), .A2(new_n632), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n888), .A2(new_n947), .ZN(new_n972));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n929), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n972), .A2(new_n693), .A3(new_n974), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n977), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n979), .A2(new_n929), .A3(new_n975), .A4(new_n968), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n978), .A2(new_n980), .ZN(G66));
  OAI21_X1  g795(.A(G953), .B1(new_n277), .B2(new_n516), .ZN(new_n982));
  INV_X1    g796(.A(new_n886), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n933), .B1(G898), .B2(new_n368), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(G69));
  AND2_X1   g800(.A1(new_n852), .A2(new_n731), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(new_n727), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n648), .A2(new_n649), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n666), .B1(new_n722), .B2(new_n525), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n708), .A2(new_n782), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n813), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n988), .A2(new_n989), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n990), .A2(new_n994), .A3(new_n819), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n368), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n583), .B(new_n498), .Z(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n774), .A2(new_n761), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n805), .A2(new_n812), .A3(new_n1002), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n813), .A2(new_n1003), .A3(new_n795), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1004), .A2(new_n819), .A3(new_n792), .A4(new_n987), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1001), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n999), .A2(new_n1000), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n368), .B1(G227), .B2(G900), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1008), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n999), .A2(new_n1000), .A3(new_n1010), .A4(new_n1006), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(G72));
  OAI21_X1  g826(.A(new_n562), .B1(new_n584), .B2(new_n559), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n928), .B1(new_n890), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n584), .A2(new_n560), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n819), .A2(new_n792), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1019), .A2(new_n983), .A3(new_n987), .A4(new_n1004), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1018), .B1(new_n1020), .B2(new_n1015), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n996), .B2(new_n886), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n1017), .B(new_n1021), .C1(new_n715), .C2(new_n1022), .ZN(G57));
endmodule


