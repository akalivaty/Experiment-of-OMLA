//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G234), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  XNOR2_X1  g013(.A(G119), .B(G128), .ZN(new_n200));
  OAI22_X1  g014(.A1(new_n198), .A2(G110), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT16), .ZN(new_n206));
  OR3_X1    g020(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G146), .ZN(new_n208));
  XNOR2_X1  g022(.A(G125), .B(G140), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n201), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n199), .A2(new_n200), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n206), .A2(G146), .A3(new_n207), .ZN(new_n214));
  AOI21_X1  g028(.A(G146), .B1(new_n206), .B2(new_n207), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT70), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n198), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n194), .A2(new_n197), .A3(KEYINPUT70), .A4(new_n195), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n212), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT71), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(G953), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n224), .B(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT71), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(new_n212), .C1(new_n216), .C2(new_n221), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n227), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n222), .A2(KEYINPUT71), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n189), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(G902), .B1(new_n230), .B2(new_n232), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT25), .B1(new_n238), .B2(KEYINPUT72), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n191), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n190), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n187), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n236), .B1(new_n234), .B2(new_n235), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n238), .A2(KEYINPUT72), .A3(KEYINPUT25), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n190), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT73), .A3(new_n242), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT11), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G137), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n252), .A2(new_n254), .A3(new_n258), .A4(new_n255), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT65), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n210), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT0), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n196), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n263), .A2(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n263), .A2(new_n265), .A3(new_n268), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n262), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n263), .A2(new_n265), .A3(new_n268), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n267), .A2(new_n268), .ZN(new_n273));
  XNOR2_X1  g087(.A(G143), .B(G146), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n272), .B(KEYINPUT64), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n257), .A2(new_n277), .A3(new_n259), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n261), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n264), .A2(KEYINPUT1), .A3(G146), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n274), .B2(G128), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n282), .A2(new_n263), .A3(new_n265), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n251), .A2(G137), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n253), .A2(G134), .ZN(new_n286));
  OAI21_X1  g100(.A(G131), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n259), .A2(new_n287), .A3(KEYINPUT66), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT66), .B1(new_n259), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n284), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(KEYINPUT30), .A3(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT2), .B(G113), .Z(new_n292));
  XNOR2_X1  g106(.A(G116), .B(G119), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n193), .A2(G116), .ZN(new_n295));
  INV_X1    g109(.A(G116), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G119), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT2), .B(G113), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n260), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n269), .A2(new_n270), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n281), .A2(new_n283), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n259), .A2(new_n287), .ZN(new_n305));
  OAI22_X1  g119(.A1(new_n302), .A2(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT30), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n291), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  NOR2_X1   g124(.A1(G237), .A2(G953), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G210), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n310), .B(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n314));
  XOR2_X1   g128(.A(new_n313), .B(new_n314), .Z(new_n315));
  NOR2_X1   g129(.A1(new_n301), .A2(KEYINPUT67), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n294), .B2(new_n300), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n279), .A2(new_n319), .A3(new_n290), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n309), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT31), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n309), .A2(KEYINPUT31), .A3(new_n315), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n306), .A2(new_n301), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n329), .B2(new_n326), .ZN(new_n330));
  INV_X1    g144(.A(new_n315), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G472), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(new_n189), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT32), .ZN(new_n336));
  AOI21_X1  g150(.A(G902), .B1(new_n325), .B2(new_n332), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n334), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n309), .A2(new_n320), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n331), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n342), .B(new_n343), .C1(new_n330), .C2(new_n331), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n320), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n279), .A2(new_n319), .A3(KEYINPUT69), .A4(new_n290), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n279), .A2(new_n290), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n319), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT28), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n327), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n315), .A2(KEYINPUT29), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n344), .B(new_n189), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G472), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n249), .B1(new_n340), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n357));
  INV_X1    g171(.A(G107), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(G104), .ZN(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n358), .A3(G104), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(KEYINPUT75), .A3(G107), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n359), .A2(new_n361), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n356), .B1(new_n365), .B2(G101), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n359), .A2(new_n364), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n361), .A2(new_n363), .ZN(new_n368));
  INV_X1    g182(.A(G101), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n356), .A3(G101), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n371), .A2(new_n301), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n374), .B(G113), .C1(KEYINPUT5), .C2(new_n295), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n294), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n365), .A2(G101), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n358), .B2(G104), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n360), .A2(KEYINPUT76), .A3(G107), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n358), .A2(G104), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n369), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n377), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n360), .A2(KEYINPUT76), .A3(G107), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT76), .B1(new_n360), .B2(G107), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G101), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n370), .A2(new_n389), .A3(KEYINPUT78), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n376), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n373), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G110), .B(G122), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n304), .A2(new_n204), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n303), .A2(G125), .ZN(new_n395));
  INV_X1    g209(.A(G224), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT7), .B1(new_n396), .B2(G953), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n395), .ZN(new_n399));
  INV_X1    g213(.A(new_n397), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n392), .A2(new_n393), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n393), .B(KEYINPUT80), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT8), .ZN(new_n404));
  INV_X1    g218(.A(new_n376), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n370), .B2(new_n389), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n406), .B2(new_n391), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n393), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n373), .B2(new_n391), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n385), .A2(new_n390), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n405), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n365), .A2(new_n356), .A3(G101), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n370), .B2(new_n366), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n301), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n415), .A3(new_n393), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n416), .A3(KEYINPUT6), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n418), .B(new_n409), .C1(new_n373), .C2(new_n391), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n396), .A2(G953), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n399), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n408), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n408), .B2(new_n422), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT79), .Z(new_n429));
  NOR2_X1   g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G237), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n225), .A3(G214), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G143), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT82), .ZN(new_n435));
  AOI211_X1 g249(.A(G143), .B(new_n435), .C1(new_n311), .C2(G214), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT82), .B1(new_n432), .B2(new_n264), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G131), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT17), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n258), .B(new_n434), .C1(new_n436), .C2(new_n437), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n214), .A2(new_n215), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n439), .A2(KEYINPUT87), .A3(new_n440), .A4(new_n441), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n438), .A2(KEYINPUT17), .A3(G131), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n444), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n209), .B(G146), .ZN(new_n449));
  INV_X1    g263(.A(new_n437), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n432), .A2(KEYINPUT82), .A3(new_n264), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n450), .A2(new_n451), .B1(G143), .B2(new_n433), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(KEYINPUT18), .A3(G131), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n449), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n438), .A2(new_n453), .A3(KEYINPUT18), .A4(G131), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G113), .B(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(new_n360), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT86), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n448), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n448), .B2(new_n457), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n189), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT88), .B(G475), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n264), .A2(G128), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT13), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n264), .A2(G128), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n251), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n196), .A2(G143), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n467), .A2(new_n474), .A3(new_n251), .ZN(new_n475));
  INV_X1    g289(.A(G122), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G116), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n296), .A2(G122), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n358), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n358), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n475), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n251), .B1(new_n467), .B2(new_n474), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n478), .A2(KEYINPUT14), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n296), .A2(G122), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n478), .B1(new_n487), .B2(KEYINPUT14), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n358), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI22_X1  g303(.A1(new_n473), .A2(new_n482), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT9), .B(G234), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n491), .A2(new_n188), .A3(G953), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI221_X1 g308(.A(new_n492), .B1(new_n482), .B2(new_n473), .C1(new_n485), .C2(new_n489), .ZN(new_n495));
  AOI21_X1  g309(.A(G902), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G478), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(G234), .A2(G237), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(G952), .A3(new_n225), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT21), .B(G898), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(G902), .A3(G953), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n439), .A2(new_n441), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n209), .A2(new_n511), .A3(KEYINPUT19), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n209), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n214), .B1(new_n514), .B2(new_n210), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n456), .A2(new_n455), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n509), .B1(new_n516), .B2(new_n459), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n510), .A2(new_n515), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n457), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n459), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(KEYINPUT85), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n461), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT20), .ZN(new_n523));
  NOR2_X1   g337(.A1(G475), .A2(G902), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n522), .B2(new_n524), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n466), .B(new_n508), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G221), .ZN(new_n530));
  INV_X1    g344(.A(new_n491), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(new_n189), .ZN(new_n532));
  INV_X1    g346(.A(G469), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n189), .ZN(new_n534));
  XOR2_X1   g348(.A(G110), .B(G140), .Z(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT74), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n225), .A2(G227), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT10), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n304), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n411), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n261), .A2(new_n278), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n371), .A2(new_n276), .A3(new_n372), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n282), .A2(new_n263), .A3(new_n265), .A4(KEYINPUT77), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n545), .B(new_n280), .C1(G128), .C2(new_n274), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n283), .A2(KEYINPUT77), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n370), .B(new_n389), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n540), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n385), .A2(new_n390), .A3(new_n304), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n548), .ZN(new_n552));
  INV_X1    g366(.A(new_n543), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT12), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n302), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n551), .B2(new_n548), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n550), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n550), .A2(new_n538), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n549), .A2(new_n544), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n284), .A2(KEYINPUT10), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n385), .B2(new_n390), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n553), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n539), .A2(new_n559), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n534), .B1(new_n565), .B2(G469), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n561), .A2(new_n563), .A3(new_n553), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n414), .A2(new_n276), .B1(new_n548), .B2(new_n540), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n543), .B1(new_n568), .B2(new_n542), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n539), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n538), .B(new_n550), .C1(new_n554), .C2(new_n558), .ZN(new_n571));
  AOI21_X1  g385(.A(G902), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n533), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n532), .B1(new_n566), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n430), .A2(new_n529), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n355), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  AOI22_X1  g391(.A1(new_n323), .A2(new_n324), .B1(new_n330), .B2(new_n331), .ZN(new_n578));
  OAI21_X1  g392(.A(G472), .B1(new_n578), .B2(G902), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n335), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n559), .A2(new_n539), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n560), .A2(new_n564), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(G469), .ZN(new_n584));
  INV_X1    g398(.A(new_n534), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n573), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n532), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n581), .A2(new_n249), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n466), .B1(new_n525), .B2(new_n527), .ZN(new_n590));
  INV_X1    g404(.A(new_n496), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT91), .A3(new_n497), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT91), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n496), .B2(G478), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n490), .B2(KEYINPUT89), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n494), .A2(new_n495), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n495), .A3(new_n494), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n497), .A2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(KEYINPUT90), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT90), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n595), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n590), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n408), .A2(new_n422), .ZN(new_n611));
  INV_X1    g425(.A(new_n423), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n424), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n428), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n610), .A2(new_n615), .A3(new_n507), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n589), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT92), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n428), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n613), .B2(new_n424), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n507), .B(KEYINPUT93), .Z(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n625), .A2(new_n527), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n499), .B1(new_n464), .B2(new_n465), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n589), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT94), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n227), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n222), .B(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(new_n241), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n247), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n575), .A2(new_n580), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT95), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(G12));
  XNOR2_X1  g456(.A(new_n502), .B(KEYINPUT96), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(G900), .B2(new_n505), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n627), .B(new_n644), .C1(new_n625), .C2(new_n527), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n588), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n338), .B1(new_n337), .B2(new_n334), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n578), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n354), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n622), .A2(new_n638), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XNOR2_X1  g467(.A(new_n644), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n574), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT40), .Z(new_n656));
  AOI21_X1  g470(.A(new_n319), .B1(new_n279), .B2(new_n290), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n345), .B2(new_n320), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n315), .B1(new_n658), .B2(new_n347), .ZN(new_n659));
  INV_X1    g473(.A(new_n321), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT97), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n349), .A2(new_n331), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n321), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n661), .A2(new_n664), .A3(new_n189), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT98), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n668), .A3(G472), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n340), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n614), .B(KEYINPUT38), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n590), .A2(new_n500), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n674), .A2(new_n621), .A3(new_n638), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n656), .A2(new_n672), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NAND3_X1  g491(.A1(new_n590), .A2(new_n609), .A3(new_n644), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n588), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n649), .A3(new_n651), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n570), .A2(new_n571), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT99), .B1(new_n683), .B2(new_n189), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  AOI211_X1 g499(.A(new_n685), .B(G902), .C1(new_n570), .C2(new_n571), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n682), .B(G469), .C1(new_n684), .C2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n552), .A2(new_n553), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n555), .ZN(new_n689));
  INV_X1    g503(.A(new_n558), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n564), .A2(new_n550), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n691), .A2(new_n560), .B1(new_n692), .B2(new_n539), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n685), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n572), .A2(KEYINPUT99), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n533), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT100), .B1(new_n572), .B2(new_n533), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n687), .B(new_n587), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n355), .A2(new_n699), .A3(new_n616), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND3_X1  g516(.A1(new_n355), .A2(new_n699), .A3(new_n629), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NAND2_X1  g518(.A1(new_n649), .A2(new_n651), .ZN(new_n705));
  OAI21_X1  g519(.A(G469), .B1(new_n684), .B2(new_n686), .ZN(new_n706));
  INV_X1    g520(.A(new_n697), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n587), .A3(new_n529), .A4(new_n687), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n193), .ZN(G21));
  NOR2_X1   g525(.A1(new_n240), .A2(new_n243), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n334), .A2(new_n189), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT101), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n315), .B1(new_n350), .B2(new_n327), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n323), .A2(new_n324), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n712), .A2(new_n579), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n622), .A2(new_n590), .A3(new_n500), .A4(new_n623), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n698), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT102), .B(G122), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G24));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n579), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n240), .A2(new_n636), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n678), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n699), .A2(new_n622), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND2_X1  g541(.A1(new_n427), .A2(new_n428), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n588), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n244), .A2(new_n248), .ZN(new_n730));
  INV_X1    g544(.A(new_n678), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n729), .A2(new_n649), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n734));
  INV_X1    g548(.A(new_n524), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n517), .A2(new_n521), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(new_n736), .B2(new_n461), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n734), .B1(new_n737), .B2(new_n526), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n608), .B1(new_n738), .B2(new_n466), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n425), .A2(new_n426), .A3(new_n621), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n574), .A3(new_n644), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n733), .ZN(new_n742));
  INV_X1    g556(.A(new_n712), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n340), .B2(new_n354), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n732), .A2(new_n733), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n258), .ZN(G33));
  NAND2_X1  g560(.A1(new_n645), .A2(KEYINPUT103), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n626), .A2(new_n748), .A3(new_n627), .A4(new_n644), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n649), .A3(new_n730), .A4(new_n729), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  XNOR2_X1  g566(.A(new_n565), .B(KEYINPUT45), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n533), .B1(new_n753), .B2(new_n189), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n755), .A2(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(KEYINPUT46), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n573), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n587), .A3(new_n654), .ZN(new_n759));
  INV_X1    g573(.A(new_n590), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n609), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT104), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT104), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n761), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n581), .A2(new_n638), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n740), .B1(new_n768), .B2(new_n769), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n759), .B(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  NAND2_X1  g589(.A1(new_n758), .A2(new_n587), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n649), .A2(new_n730), .A3(new_n678), .A4(new_n728), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  INV_X1    g595(.A(new_n672), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n698), .A2(new_n728), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n730), .A2(new_n782), .A3(new_n503), .A4(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n760), .A3(new_n608), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n766), .A2(new_n643), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT110), .Z(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n783), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n723), .A2(new_n724), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n792));
  INV_X1    g606(.A(new_n718), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n673), .A2(new_n428), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n698), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n792), .B(KEYINPUT50), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n792), .A2(KEYINPUT50), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n794), .A2(new_n698), .A3(new_n799), .A4(new_n796), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n791), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n803), .B(new_n791), .C1(new_n798), .C2(new_n800), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n708), .A2(new_n532), .A3(new_n687), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n795), .B(new_n740), .C1(new_n778), .C2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n802), .A2(KEYINPUT51), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n724), .A2(new_n586), .A3(new_n587), .A4(new_n644), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n622), .A2(new_n590), .A3(new_n500), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n340), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n670), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n726), .A2(new_n814), .A3(new_n652), .A4(new_n680), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT52), .Z(new_n816));
  AND2_X1   g630(.A1(new_n499), .A2(new_n644), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n466), .A2(new_n638), .A3(new_n626), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n729), .A3(new_n649), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n679), .A2(new_n790), .A3(new_n740), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n751), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n745), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n650), .B1(new_n340), .B2(new_n354), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n699), .A3(new_n529), .ZN(new_n824));
  INV_X1    g638(.A(new_n719), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n699), .A2(new_n793), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n700), .A2(new_n703), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n610), .B1(new_n590), .B2(new_n499), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n430), .A2(new_n623), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n589), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n576), .A3(new_n639), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n827), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n816), .A2(new_n822), .A3(new_n833), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n700), .A2(new_n703), .A3(new_n824), .A4(new_n826), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT106), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT107), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n827), .A2(KEYINPUT106), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n822), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n710), .A2(new_n720), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n836), .A3(new_n700), .A4(new_n703), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n830), .A2(new_n576), .A3(new_n639), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n839), .A2(new_n842), .A3(new_n843), .A4(new_n822), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT107), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n840), .A2(new_n845), .A3(new_n816), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n834), .B1(new_n846), .B2(new_n832), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n832), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n815), .B(KEYINPUT52), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n844), .B2(KEYINPUT107), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(KEYINPUT53), .A3(new_n840), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n809), .B(new_n849), .C1(new_n854), .C2(new_n848), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n848), .B1(new_n850), .B2(new_n853), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT53), .B1(new_n852), .B2(new_n840), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(KEYINPUT54), .A3(new_n834), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT108), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n795), .A2(new_n622), .A3(new_n699), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n225), .A2(G952), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n784), .B2(new_n739), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT48), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n789), .B2(new_n744), .ZN(new_n864));
  INV_X1    g678(.A(new_n744), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n788), .A2(KEYINPUT48), .A3(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n860), .B(new_n862), .C1(new_n864), .C2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n791), .B(new_n807), .C1(new_n798), .C2(new_n800), .ZN(new_n868));
  XNOR2_X1  g682(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n808), .A2(new_n855), .A3(new_n859), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n708), .A2(new_n687), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT49), .Z(new_n874));
  OR2_X1    g688(.A1(new_n532), .A2(new_n429), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n673), .A2(new_n761), .A3(new_n743), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n782), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n877), .ZN(G75));
  NOR2_X1   g692(.A1(new_n225), .A2(G952), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n417), .A2(new_n419), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n421), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n847), .A2(new_n189), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n612), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT114), .B1(new_n847), .B2(new_n189), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n612), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n883), .A2(new_n886), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n879), .B(new_n887), .C1(new_n891), .C2(new_n892), .ZN(G51));
  XNOR2_X1  g707(.A(new_n847), .B(new_n848), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n534), .B(KEYINPUT57), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n693), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n753), .A2(new_n533), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n889), .A2(new_n898), .A3(new_n890), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n899), .A2(new_n897), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n879), .B1(new_n900), .B2(new_n901), .ZN(G54));
  AND2_X1   g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n889), .A2(new_n890), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n461), .A3(new_n736), .ZN(new_n905));
  INV_X1    g719(.A(new_n879), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n889), .A2(new_n522), .A3(new_n890), .A4(new_n903), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT116), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n905), .A2(new_n910), .A3(new_n906), .A4(new_n907), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(G60));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT59), .Z(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n602), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n879), .B1(new_n894), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n855), .B2(new_n859), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n602), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT117), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n921), .B(new_n917), .C1(new_n918), .C2(new_n602), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(G63));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n188), .A2(new_n189), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n857), .B2(new_n834), .ZN(new_n928));
  INV_X1    g742(.A(new_n233), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n879), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n635), .B(new_n927), .C1(new_n857), .C2(new_n834), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n924), .B(KEYINPUT61), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n927), .ZN(new_n933));
  INV_X1    g747(.A(new_n834), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n850), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n906), .B(new_n931), .C1(new_n935), .C2(new_n233), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT119), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n929), .B1(new_n847), .B2(new_n933), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n940), .A2(KEYINPUT61), .A3(new_n906), .A4(new_n931), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT120), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n930), .A2(new_n943), .A3(KEYINPUT61), .A4(new_n931), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT121), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n936), .A2(new_n937), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n924), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n936), .A2(KEYINPUT119), .A3(new_n937), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n942), .A2(new_n944), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT121), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n946), .A2(new_n953), .ZN(G66));
  NOR3_X1   g768(.A1(new_n504), .A2(new_n396), .A3(new_n225), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n837), .A2(new_n839), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n957), .B2(new_n225), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n880), .B1(G898), .B2(new_n225), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G69));
  AOI21_X1  g774(.A(new_n225), .B1(G227), .B2(G900), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT123), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n726), .A2(new_n652), .A3(new_n680), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n676), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  NOR2_X1   g780(.A1(new_n655), .A2(new_n728), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n355), .A2(new_n828), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n774), .A2(new_n780), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n291), .A2(new_n308), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n514), .B(KEYINPUT122), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n969), .A2(new_n225), .A3(new_n973), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n865), .A2(new_n811), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n751), .B1(new_n759), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g790(.A(new_n963), .B(new_n976), .C1(new_n778), .C2(new_n779), .ZN(new_n977));
  INV_X1    g791(.A(new_n745), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n774), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n973), .B1(new_n979), .B2(new_n225), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n962), .B1(new_n974), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(G900), .B1(new_n972), .B2(G227), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(G953), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(G72));
  NOR2_X1   g798(.A1(new_n341), .A2(new_n315), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n979), .A2(new_n956), .ZN(new_n986));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(KEYINPUT125), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT125), .B1(new_n986), .B2(new_n988), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n342), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n988), .B1(new_n993), .B2(new_n660), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT126), .Z(new_n995));
  NOR2_X1   g809(.A1(new_n854), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT127), .Z(new_n997));
  OAI21_X1  g811(.A(new_n988), .B1(new_n969), .B2(new_n956), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1000), .A2(new_n315), .A3(new_n341), .A4(new_n1001), .ZN(new_n1002));
  AND4_X1   g816(.A1(new_n906), .A2(new_n992), .A3(new_n997), .A4(new_n1002), .ZN(G57));
endmodule


