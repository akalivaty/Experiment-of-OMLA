//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n208), .A2(new_n209), .B1(new_n202), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n211), .B(new_n217), .C1(G116), .C2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT68), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n222), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n219), .A2(new_n213), .ZN(new_n234));
  OR2_X1    g0034(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n235), .A2(G50), .A3(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT67), .Z(new_n238));
  AOI21_X1  g0038(.A(new_n230), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g0039(.A1(new_n225), .A2(new_n229), .A3(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n220), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n209), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  INV_X1    g0047(.A(G264), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G270), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G358));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(new_n202), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(G107), .ZN(new_n256));
  INV_X1    g0056(.A(G116), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n254), .B(new_n258), .ZN(G351));
  INV_X1    g0059(.A(KEYINPUT12), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n260), .B1(new_n262), .B2(G68), .ZN(new_n263));
  INV_X1    g0063(.A(new_n262), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(KEYINPUT12), .A3(new_n213), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n231), .B1(new_n222), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n261), .A2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n263), .B(new_n265), .C1(new_n272), .C2(new_n213), .ZN(new_n273));
  XOR2_X1   g0073(.A(new_n273), .B(KEYINPUT78), .Z(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n232), .A2(G33), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n276), .A2(new_n208), .B1(new_n277), .B2(new_n202), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n232), .A2(G68), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n267), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n280), .B(KEYINPUT11), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G226), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(G232), .A3(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G97), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n231), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT71), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT77), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n291), .B2(new_n231), .ZN(new_n299));
  AND2_X1   g0099(.A1(G1), .A2(G13), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(KEYINPUT70), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  AOI21_X1  g0105(.A(G1), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(G274), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT77), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n306), .B1(new_n299), .B2(new_n302), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G238), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n297), .A2(new_n307), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT13), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n295), .A2(new_n296), .B1(G238), .B2(new_n309), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n307), .A4(new_n308), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n284), .B1(new_n316), .B2(G169), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI211_X1 g0118(.A(KEYINPUT14), .B(new_n318), .C1(new_n312), .C2(new_n315), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n312), .A2(G179), .A3(new_n315), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n283), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n316), .A2(G200), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n312), .A2(G190), .A3(new_n315), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n283), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n328));
  INV_X1    g0128(.A(G107), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n285), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n334), .A2(new_n220), .A3(G1698), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n294), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n309), .A2(G244), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n307), .A3(new_n337), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(G179), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n318), .ZN(new_n340));
  INV_X1    g0140(.A(new_n272), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G77), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT8), .B(G58), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n343), .A2(new_n276), .B1(new_n232), .B2(new_n202), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT15), .B(G87), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n277), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n267), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n264), .A2(new_n202), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT73), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n342), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n339), .A2(new_n340), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n338), .A2(G200), .ZN(new_n352));
  INV_X1    g0152(.A(new_n350), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n352), .B(new_n353), .C1(new_n354), .C2(new_n338), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT74), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n275), .A2(G150), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n359), .B1(new_n201), .B2(new_n232), .C1(new_n343), .C2(new_n277), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n267), .B1(new_n208), .B2(new_n264), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n208), .B2(new_n272), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT9), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT75), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n285), .A2(G223), .A3(G1698), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(new_n202), .C2(new_n285), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n294), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n309), .A2(G226), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n307), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(new_n354), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n367), .A2(new_n374), .A3(KEYINPUT76), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(G200), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n366), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT10), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT10), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n366), .A2(new_n375), .A3(new_n379), .A4(new_n376), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT79), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n332), .A2(new_n333), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n331), .A2(KEYINPUT79), .A3(G33), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n232), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT7), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT80), .B(KEYINPUT7), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n388), .A2(new_n383), .A3(new_n232), .A4(new_n384), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(G68), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(G58), .B(G68), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(G20), .B1(G159), .B2(new_n275), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n387), .B1(new_n285), .B2(G20), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n334), .A2(new_n395), .A3(new_n232), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n396), .A3(G68), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n392), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n393), .A2(new_n267), .A3(new_n400), .ZN(new_n401));
  XOR2_X1   g0201(.A(KEYINPUT8), .B(G58), .Z(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n262), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n341), .B2(new_n402), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n309), .A2(G232), .ZN(new_n405));
  INV_X1    g0205(.A(G87), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n266), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n383), .B2(new_n384), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n286), .A2(G226), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n292), .B(KEYINPUT71), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n307), .B(new_n405), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G200), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n410), .B(new_n408), .C1(new_n383), .C2(new_n384), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n294), .B1(new_n416), .B2(new_n407), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n417), .A2(G190), .A3(new_n307), .A4(new_n405), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n401), .A2(new_n404), .A3(new_n415), .A4(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n401), .A2(new_n404), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(G169), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n417), .A2(G179), .A3(new_n307), .A4(new_n405), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n422), .A2(KEYINPUT18), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT18), .B1(new_n422), .B2(new_n425), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n420), .A2(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n373), .A2(new_n318), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n362), .B1(new_n373), .B2(G179), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n356), .A2(new_n357), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n381), .A2(new_n429), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n327), .A2(new_n358), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n383), .A2(new_n384), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n216), .A2(G1698), .ZN(new_n439));
  OR2_X1    g0239(.A1(G250), .A2(G1698), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G294), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n266), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n261), .B(G45), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n291), .A2(new_n298), .A3(new_n231), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT70), .B1(new_n300), .B2(new_n301), .ZN(new_n450));
  OAI211_X1 g0250(.A(G264), .B(new_n448), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT87), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT87), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n303), .A2(new_n453), .A3(G264), .A4(new_n448), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n445), .A2(new_n294), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n448), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n303), .A3(G274), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G169), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(G179), .A3(new_n457), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT85), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n438), .A2(new_n232), .A3(G87), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n406), .A2(G20), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(new_n332), .A3(new_n333), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n285), .A2(KEYINPUT84), .A3(new_n466), .A4(new_n465), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n464), .A2(KEYINPUT22), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n232), .B2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n329), .A2(KEYINPUT23), .A3(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G116), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n473), .A2(new_n474), .B1(new_n476), .B2(new_n232), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n463), .B1(new_n471), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(G20), .B1(new_n383), .B2(new_n384), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n466), .B1(new_n480), .B2(G87), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n469), .A2(new_n470), .ZN(new_n482));
  OAI211_X1 g0282(.A(KEYINPUT85), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(KEYINPUT24), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n463), .B(new_n485), .C1(new_n471), .C2(new_n478), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n267), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n264), .A2(new_n329), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT25), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n261), .A2(G33), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n268), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT81), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n491), .B(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n489), .B1(new_n493), .B2(G107), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n487), .A2(KEYINPUT86), .A3(new_n494), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n462), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n248), .A2(G1698), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n438), .B(new_n500), .C1(G257), .C2(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n334), .A2(G303), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n413), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G179), .ZN(new_n504));
  INV_X1    g0304(.A(new_n457), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n303), .A2(G270), .A3(new_n448), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR4_X1   g0307(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n268), .A2(G116), .A3(new_n490), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n510), .B(new_n232), .C1(G33), .C2(new_n215), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n511), .B(new_n267), .C1(new_n232), .C2(G116), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT20), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n512), .A2(new_n513), .ZN(new_n515));
  OAI221_X1 g0315(.A(new_n509), .B1(G116), .B2(new_n262), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n501), .A2(new_n502), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n505), .B1(new_n518), .B2(new_n294), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n506), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(new_n516), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n354), .C2(new_n520), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n516), .A3(G169), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n520), .A2(new_n516), .A3(KEYINPUT21), .A4(G169), .ZN(new_n527));
  AND4_X1   g0327(.A1(new_n517), .A2(new_n523), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n261), .A2(G45), .ZN(new_n530));
  OAI211_X1 g0330(.A(G250), .B(new_n530), .C1(new_n449), .C2(new_n450), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n298), .A2(new_n261), .A3(G45), .A4(G274), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G238), .A2(G1698), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n286), .A2(G244), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n438), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n475), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n533), .B1(new_n539), .B2(new_n294), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n318), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT83), .ZN(new_n543));
  AOI211_X1 g0343(.A(G20), .B(new_n213), .C1(new_n383), .C2(new_n384), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n289), .A2(KEYINPUT19), .A3(G20), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n205), .A2(new_n406), .B1(new_n289), .B2(new_n232), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n547), .B2(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n480), .A2(G68), .ZN(new_n550));
  INV_X1    g0350(.A(new_n545), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(KEYINPUT83), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n554), .A3(new_n267), .ZN(new_n555));
  INV_X1    g0355(.A(new_n345), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n491), .A2(new_n492), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT81), .B1(new_n268), .B2(new_n490), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n345), .A2(new_n264), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n540), .A2(new_n504), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n542), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n540), .A2(G190), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n413), .B1(new_n475), .B2(new_n538), .ZN(new_n565));
  OAI21_X1  g0365(.A(G200), .B1(new_n565), .B2(new_n533), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n493), .A2(G87), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n560), .A3(new_n555), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n455), .A2(G190), .A3(new_n457), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n458), .A2(G200), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n487), .A2(new_n494), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(G1698), .B1(new_n383), .B2(new_n384), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT4), .B1(new_n575), .B2(G244), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n332), .A2(new_n333), .A3(G250), .A4(G1698), .ZN(new_n577));
  AND2_X1   g0377(.A1(KEYINPUT4), .A2(G244), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n332), .A2(new_n333), .A3(new_n578), .A4(new_n286), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n579), .A3(new_n510), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n294), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n303), .A2(G257), .A3(new_n448), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n457), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT82), .ZN(new_n584));
  INV_X1    g0384(.A(new_n580), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n210), .B(G1698), .C1(new_n383), .C2(new_n384), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(KEYINPUT4), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n505), .B1(new_n587), .B2(new_n294), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT82), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n582), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n584), .A2(new_n590), .A3(G200), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n493), .A2(G97), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT6), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n215), .A2(new_n329), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(new_n205), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n329), .A2(KEYINPUT6), .A3(G97), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G20), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n394), .A2(new_n396), .A3(G107), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(new_n202), .C2(new_n276), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n267), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n592), .B(new_n601), .C1(G97), .C2(new_n262), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n583), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G190), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n591), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n504), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n583), .A2(new_n318), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n602), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n571), .A2(new_n574), .A3(new_n606), .A4(new_n609), .ZN(new_n610));
  NOR4_X1   g0410(.A1(new_n437), .A2(new_n499), .A3(new_n529), .A4(new_n610), .ZN(G372));
  INV_X1    g0411(.A(KEYINPUT89), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n419), .B(KEYINPUT17), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n326), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n351), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n615), .B1(new_n322), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n401), .A2(new_n404), .B1(new_n423), .B2(new_n424), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n618), .B(KEYINPUT18), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n617), .A2(new_n619), .B1(new_n378), .B2(new_n380), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n612), .B1(new_n620), .B2(new_n432), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n316), .A2(G169), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT14), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n316), .A2(new_n284), .A3(G169), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n321), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n616), .B1(new_n625), .B2(new_n282), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n619), .B1(new_n626), .B2(new_n614), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n381), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(KEYINPUT89), .A3(new_n433), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  AOI221_X4 g0430(.A(KEYINPUT88), .B1(new_n459), .B2(new_n460), .C1(new_n487), .C2(new_n494), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT88), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n495), .B2(new_n461), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n526), .A2(new_n517), .A3(new_n527), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n610), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n609), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n571), .A2(new_n638), .A3(KEYINPUT26), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n542), .A2(new_n561), .A3(new_n562), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n569), .B2(new_n567), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n642), .B2(new_n609), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n641), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n630), .B1(new_n437), .B2(new_n646), .ZN(G369));
  INV_X1    g0447(.A(new_n498), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT86), .B1(new_n487), .B2(new_n494), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n461), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n261), .A2(new_n232), .A3(G13), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT27), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(new_n261), .A3(new_n232), .A4(G13), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n652), .A2(G213), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G343), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT90), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n648), .B2(new_n649), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n650), .A2(new_n658), .A3(new_n574), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n499), .A2(new_n657), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n657), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n522), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n635), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n529), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT91), .Z(new_n669));
  NAND2_X1  g0469(.A1(new_n635), .A2(new_n663), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT92), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n661), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n634), .A2(new_n657), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n669), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n226), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n237), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n663), .B1(new_n637), .B2(new_n645), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(KEYINPUT93), .A2(KEYINPUT31), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n588), .A2(new_n455), .A3(new_n540), .A4(new_n582), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n519), .A2(G179), .A3(new_n506), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(G179), .B1(new_n519), .B2(new_n506), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n458), .A3(new_n541), .A4(new_n583), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n445), .A2(new_n294), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n452), .A2(new_n454), .ZN(new_n695));
  AOI211_X1 g0495(.A(new_n534), .B(new_n536), .C1(new_n383), .C2(new_n384), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n294), .B1(new_n696), .B2(new_n476), .ZN(new_n697));
  INV_X1    g0497(.A(new_n533), .ZN(new_n698));
  AND4_X1   g0498(.A1(new_n694), .A2(new_n695), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n604), .A2(new_n699), .A3(new_n508), .A4(KEYINPUT30), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n691), .A2(new_n693), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n657), .ZN(new_n702));
  NAND2_X1  g0502(.A1(KEYINPUT93), .A2(KEYINPUT31), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n687), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI211_X1 g0504(.A(KEYINPUT93), .B(KEYINPUT31), .C1(new_n701), .C2(new_n657), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AND4_X1   g0507(.A1(new_n571), .A2(new_n574), .A3(new_n606), .A4(new_n609), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n650), .A3(new_n528), .A4(new_n663), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(G330), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n708), .B1(new_n499), .B2(new_n635), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n563), .B1(new_n639), .B2(new_n643), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n657), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n686), .A2(new_n711), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n683), .B1(new_n719), .B2(G1), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT94), .ZN(G364));
  AOI21_X1  g0521(.A(new_n231), .B1(G20), .B2(new_n318), .ZN(new_n722));
  INV_X1    g0522(.A(G303), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n232), .A2(new_n354), .ZN(new_n724));
  INV_X1    g0524(.A(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G179), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n354), .A2(G20), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n728), .A2(new_n504), .A3(G200), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n334), .B1(new_n723), .B2(new_n727), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n728), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n504), .A2(new_n725), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G317), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT33), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n737), .A2(KEYINPUT33), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n733), .A2(new_n726), .ZN(new_n742));
  INV_X1    g0542(.A(G322), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n504), .A2(G200), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n724), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n740), .B1(new_n741), .B2(new_n742), .C1(new_n743), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT95), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n728), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n732), .B(new_n747), .C1(G329), .C2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(G20), .B1(new_n749), .B2(new_n354), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n751), .B1(new_n442), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n734), .A2(new_n724), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n754), .B1(G326), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT96), .ZN(new_n758));
  INV_X1    g0558(.A(new_n742), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G107), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n219), .B2(new_n746), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n285), .B1(new_n208), .B2(new_n755), .C1(new_n730), .C2(new_n202), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n727), .A2(new_n406), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT32), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n750), .B2(G159), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G97), .B2(new_n752), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n750), .A2(new_n765), .A3(G159), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n764), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G68), .B2(new_n736), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n722), .B1(new_n758), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n238), .A2(new_n305), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n438), .A2(new_n677), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(new_n305), .C2(new_n254), .ZN(new_n774));
  NAND3_X1  g0574(.A1(G355), .A2(new_n285), .A3(new_n226), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n774), .B(new_n775), .C1(G116), .C2(new_n226), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n722), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G13), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G45), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n679), .A2(G1), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n771), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n789));
  INV_X1    g0589(.A(new_n779), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n788), .B(new_n789), .C1(new_n666), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n786), .B1(new_n666), .B2(G330), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G330), .B2(new_n666), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(G396));
  INV_X1    g0594(.A(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n657), .A2(new_n350), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT98), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n356), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT98), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n796), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n800), .A2(KEYINPUT99), .A3(new_n351), .A4(new_n355), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n663), .B(new_n802), .C1(new_n637), .C2(new_n645), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n646), .A2(new_n657), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n616), .A2(new_n657), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n798), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(new_n711), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n711), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(new_n785), .A3(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n736), .A2(G150), .B1(new_n756), .B2(G137), .ZN(new_n811));
  INV_X1    g0611(.A(G143), .ZN(new_n812));
  INV_X1    g0612(.A(G159), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n812), .B2(new_n746), .C1(new_n813), .C2(new_n730), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT34), .Z(new_n815));
  NOR2_X1   g0615(.A1(new_n742), .A2(new_n213), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n750), .B2(G132), .ZN(new_n817));
  INV_X1    g0617(.A(new_n438), .ZN(new_n818));
  INV_X1    g0618(.A(new_n727), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(G50), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(new_n219), .C2(new_n753), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n742), .A2(new_n406), .B1(new_n727), .B2(new_n329), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n334), .B1(new_n755), .B2(new_n723), .C1(new_n741), .C2(new_n735), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(G116), .C2(new_n729), .ZN(new_n824));
  INV_X1    g0624(.A(new_n750), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n215), .B2(new_n753), .C1(new_n731), .C2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n746), .A2(new_n442), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n815), .A2(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n722), .A2(new_n777), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n828), .A2(new_n722), .B1(new_n202), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n786), .B(new_n830), .C1(new_n806), .C2(new_n778), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT100), .Z(new_n832));
  NAND2_X1  g0632(.A1(new_n810), .A2(new_n832), .ZN(G384));
  OAI21_X1  g0633(.A(G77), .B1(new_n219), .B2(new_n213), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n237), .A2(new_n834), .B1(G50), .B2(new_n213), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(G1), .A3(new_n782), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT101), .Z(new_n837));
  AOI21_X1  g0637(.A(new_n257), .B1(new_n597), .B2(KEYINPUT35), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n838), .B(new_n233), .C1(KEYINPUT35), .C2(new_n597), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT36), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT102), .Z(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT103), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n618), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n422), .A2(new_n655), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n419), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n618), .A2(new_n845), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n393), .A2(new_n267), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT16), .B1(new_n390), .B2(new_n392), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n404), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n425), .B2(new_n655), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n419), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n849), .A2(new_n850), .B1(KEYINPUT37), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n655), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n619), .B2(new_n613), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n843), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n422), .A2(new_n425), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT37), .B1(new_n860), .B2(KEYINPUT103), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n861), .A2(new_n419), .A3(new_n850), .A4(new_n847), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n857), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n428), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n806), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n282), .A2(new_n657), .ZN(new_n870));
  INV_X1    g0670(.A(new_n321), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n317), .A2(new_n319), .A3(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n326), .B(new_n870), .C1(new_n872), .C2(new_n283), .ZN(new_n873));
  INV_X1    g0673(.A(new_n326), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n282), .B(new_n657), .C1(new_n625), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n869), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT104), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(KEYINPUT31), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n702), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n702), .A2(new_n878), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n709), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g0681(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n876), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n876), .A2(new_n881), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n868), .B(new_n883), .C1(new_n884), .C2(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n876), .A2(new_n881), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n860), .A2(new_n847), .A3(new_n419), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n849), .A2(new_n850), .B1(KEYINPUT37), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n847), .B1(new_n619), .B2(new_n613), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n843), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(new_n867), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT40), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n436), .A2(new_n881), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(G330), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n436), .B1(new_n685), .B2(new_n716), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n630), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n351), .A2(new_n657), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n803), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n873), .A2(new_n875), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n868), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n619), .A2(new_n655), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n323), .A2(new_n657), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n890), .A2(new_n906), .A3(new_n867), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n859), .B2(new_n867), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n898), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n896), .B(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n783), .A2(new_n261), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n842), .B1(new_n912), .B2(new_n913), .ZN(G367));
  OAI22_X1  g0714(.A1(new_n735), .A2(new_n813), .B1(new_n755), .B2(new_n812), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n730), .A2(new_n208), .B1(new_n219), .B2(new_n727), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(G137), .C2(new_n750), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n752), .A2(G68), .ZN(new_n918));
  INV_X1    g0718(.A(G150), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n746), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n285), .B1(new_n742), .B2(new_n202), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT108), .Z(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT107), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n727), .B2(new_n257), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(KEYINPUT46), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(KEYINPUT46), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n737), .C2(new_n825), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n735), .A2(new_n442), .B1(new_n755), .B2(new_n731), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(G97), .B2(new_n759), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n438), .B1(G303), .B2(new_n745), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n930), .B(new_n931), .C1(new_n329), .C2(new_n753), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n928), .B(new_n932), .C1(G283), .C2(new_n729), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n923), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT47), .Z(new_n935));
  AOI21_X1  g0735(.A(new_n785), .B1(new_n935), .B2(new_n722), .ZN(new_n936));
  INV_X1    g0736(.A(new_n773), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n780), .B1(new_n226), .B2(new_n345), .C1(new_n250), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n569), .A2(new_n657), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n642), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n779), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n936), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n784), .A2(G1), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n606), .B(new_n609), .C1(new_n603), .C2(new_n663), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n638), .A2(new_n657), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n675), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT44), .Z(new_n949));
  NAND3_X1  g0749(.A1(new_n672), .A2(new_n674), .A3(new_n946), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n669), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n662), .A2(new_n667), .ZN(new_n955));
  INV_X1    g0755(.A(new_n668), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n671), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n671), .ZN(new_n958));
  INV_X1    g0758(.A(new_n955), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n668), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n718), .ZN(new_n962));
  INV_X1    g0762(.A(new_n669), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n949), .A2(new_n952), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n954), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n719), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n678), .B(KEYINPUT41), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n943), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n672), .A2(KEYINPUT42), .A3(new_n947), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT42), .B1(new_n672), .B2(new_n947), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n638), .B1(new_n499), .B2(new_n606), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n970), .C1(new_n657), .C2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT106), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n940), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(KEYINPUT106), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n940), .B(KEYINPUT43), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n973), .B2(new_n976), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n963), .A2(new_n947), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n977), .B2(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n942), .B1(new_n968), .B2(new_n983), .ZN(G387));
  AND2_X1   g0784(.A1(new_n750), .A2(G326), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n745), .A2(G317), .B1(new_n729), .B2(G303), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n731), .B2(new_n735), .C1(new_n743), .C2(new_n755), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT111), .Z(new_n988));
  AOI22_X1  g0788(.A1(new_n988), .A2(KEYINPUT48), .B1(G283), .B2(new_n752), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(KEYINPUT48), .B2(new_n988), .C1(new_n442), .C2(new_n727), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT49), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n438), .B(new_n985), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n991), .B2(new_n990), .C1(new_n257), .C2(new_n742), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n753), .A2(new_n345), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n746), .A2(new_n208), .B1(new_n813), .B2(new_n755), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n402), .B2(new_n736), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n213), .B2(new_n730), .C1(new_n202), .C2(new_n727), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n994), .B(new_n997), .C1(G150), .C2(new_n750), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n998), .B(new_n438), .C1(new_n215), .C2(new_n742), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT110), .Z(new_n1000));
  NAND2_X1  g0800(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n785), .B1(new_n1001), .B2(new_n722), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n662), .A2(new_n779), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n343), .A2(G50), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n680), .B1(new_n213), .B2(new_n202), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  AOI211_X1 g0807(.A(G45), .B(new_n1007), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n773), .B1(new_n245), .B2(new_n305), .ZN(new_n1009));
  OR3_X1    g0809(.A1(new_n680), .A2(new_n677), .A3(new_n334), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n226), .A2(G107), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n780), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n961), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1004), .A2(new_n1013), .B1(new_n1014), .B2(new_n943), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n962), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n678), .B(KEYINPUT112), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1014), .A2(new_n719), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(G393));
  INV_X1    g0821(.A(KEYINPUT113), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n954), .A2(new_n1022), .A3(new_n964), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n964), .A2(new_n1022), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n1016), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(new_n965), .A3(new_n1018), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n947), .A2(new_n779), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n780), .B1(new_n215), .B2(new_n226), .C1(new_n258), .C2(new_n937), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n753), .A2(new_n257), .B1(new_n723), .B2(new_n735), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT116), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n756), .A2(G317), .B1(new_n745), .B2(G311), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT52), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n825), .A2(new_n743), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n760), .B(new_n334), .C1(new_n442), .C2(new_n730), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n1030), .B2(new_n1029), .C1(new_n741), .C2(new_n727), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n756), .A2(G150), .B1(new_n745), .B2(G159), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT115), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT114), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n753), .A2(new_n202), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n759), .A2(G87), .B1(new_n402), .B2(new_n729), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n438), .C1(new_n213), .C2(new_n727), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(G143), .C2(new_n750), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n208), .B2(new_n735), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1037), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n785), .B1(new_n1047), .B2(new_n722), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1027), .A2(new_n1028), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n943), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1026), .A2(new_n1051), .ZN(G390));
  NOR2_X1   g0852(.A1(new_n907), .A2(new_n908), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n873), .A2(new_n875), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n803), .B2(new_n900), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1055), .B2(new_n905), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n891), .A2(new_n905), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n899), .B1(new_n714), .B2(new_n802), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n1054), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n806), .A2(G330), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n706), .B2(new_n709), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n1054), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1056), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1060), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n881), .A2(new_n902), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT117), .B1(new_n1061), .B2(new_n902), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n1066), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1061), .A2(KEYINPUT117), .A3(new_n902), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n901), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n881), .A2(new_n1065), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n1054), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n1058), .C1(new_n1054), .C2(new_n1062), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n436), .A2(G330), .A3(new_n881), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n630), .A2(new_n897), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1069), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1079), .B(new_n1077), .C1(new_n1064), .C2(new_n1068), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n1018), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1053), .A2(new_n777), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT54), .B(G143), .Z(new_n1085));
  AOI22_X1  g0885(.A1(new_n759), .A2(G50), .B1(new_n729), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(G128), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n755), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G125), .B2(new_n750), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n745), .A2(G132), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n752), .A2(G159), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n727), .A2(KEYINPUT53), .A3(new_n919), .ZN(new_n1092));
  OAI21_X1  g0892(.A(KEYINPUT53), .B1(new_n727), .B2(new_n919), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n285), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(G137), .C2(new_n736), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n736), .A2(G107), .B1(new_n745), .B2(G116), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n215), .B2(new_n730), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1098), .A2(new_n285), .A3(new_n763), .A4(new_n816), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n202), .B2(new_n753), .C1(new_n442), .C2(new_n825), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n755), .A2(new_n741), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(new_n722), .B1(new_n343), .B2(new_n829), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1084), .A2(new_n786), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1069), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n943), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1083), .A2(new_n1106), .ZN(G378));
  OAI21_X1  g0907(.A(new_n1079), .B1(new_n1069), .B2(new_n1080), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n893), .A2(G330), .A3(new_n910), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n910), .B1(new_n893), .B2(G330), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n362), .A2(new_n655), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n381), .A2(new_n433), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n381), .B2(new_n433), .ZN(new_n1113));
  OR3_X1    g0913(.A1(new_n1112), .A2(new_n1113), .A3(KEYINPUT55), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT55), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1114), .A2(KEYINPUT56), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT56), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1109), .A2(new_n1110), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n876), .A2(new_n881), .A3(new_n882), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT105), .B1(new_n876), .B2(new_n881), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n868), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n892), .ZN(new_n1125));
  OAI21_X1  g0925(.A(G330), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n910), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n893), .A2(G330), .A3(new_n910), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1118), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1108), .B(KEYINPUT57), .C1(new_n1120), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1018), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT122), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT122), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1134), .A3(new_n1018), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT123), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1119), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1128), .A2(new_n1118), .A3(new_n1129), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1137), .A2(new_n1138), .B1(new_n1082), .B2(new_n1079), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1136), .B1(new_n1139), .B2(KEYINPUT57), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1108), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(KEYINPUT123), .A3(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1133), .A2(new_n1135), .A3(new_n1140), .A4(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n736), .A2(G97), .B1(new_n745), .B2(G107), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n825), .B2(new_n741), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n304), .B1(new_n727), .B2(new_n202), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n818), .B1(new_n345), .B2(new_n730), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n742), .A2(new_n219), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n918), .C1(new_n257), .C2(new_n755), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT118), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(KEYINPUT58), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n752), .A2(G150), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G125), .A2(new_n756), .B1(new_n819), .B2(new_n1085), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n736), .A2(G132), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n745), .A2(G128), .B1(new_n729), .B2(G137), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G33), .B1(new_n759), .B2(G159), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT119), .B(G124), .Z(new_n1162));
  OAI211_X1 g0962(.A(new_n304), .B(new_n1161), .C1(new_n825), .C2(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT120), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(KEYINPUT120), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1160), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1153), .A2(KEYINPUT58), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n304), .B1(new_n818), .B2(new_n266), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n208), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1154), .A2(new_n1167), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1171), .A2(new_n722), .B1(new_n208), .B2(new_n829), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n786), .B(new_n1172), .C1(new_n1119), .C2(new_n778), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT121), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1141), .B2(new_n943), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1145), .A2(new_n1179), .ZN(G375));
  NAND3_X1  g0980(.A1(new_n630), .A2(new_n897), .A3(new_n1078), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT124), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n1073), .A3(KEYINPUT124), .A4(new_n1076), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n967), .A3(new_n1080), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT125), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n1054), .A2(new_n777), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n730), .A2(new_n329), .B1(new_n257), .B2(new_n735), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n334), .B1(new_n202), .B2(new_n742), .C1(new_n746), .C2(new_n741), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(G97), .C2(new_n819), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n994), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n756), .A2(G294), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n750), .A2(G303), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n756), .A2(G132), .B1(new_n729), .B2(G150), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n745), .A2(G137), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n813), .C2(new_n727), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n736), .B2(new_n1085), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n752), .A2(G50), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n750), .A2(G128), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1200), .A2(new_n438), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1196), .B1(new_n1203), .B2(new_n1150), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1204), .A2(new_n722), .B1(new_n213), .B2(new_n829), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1189), .A2(new_n786), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1077), .B2(new_n943), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1188), .A2(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(G378), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1145), .A2(new_n1210), .A3(new_n1179), .ZN(new_n1211));
  INV_X1    g1011(.A(G396), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(new_n1015), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(G387), .A2(G390), .A3(G384), .A4(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1214), .A3(new_n1208), .A4(new_n1188), .ZN(G407));
  INV_X1    g1015(.A(G343), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(G407), .A2(G213), .A3(new_n1217), .ZN(G409));
  INV_X1    g1018(.A(KEYINPUT127), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1213), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1026), .A2(new_n1051), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1026), .B2(new_n1051), .ZN(new_n1223));
  OAI21_X1  g1023(.A(G387), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1221), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G390), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n942), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n966), .A2(new_n967), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n943), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n981), .A2(new_n982), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1227), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1026), .A2(new_n1051), .A3(new_n1221), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1226), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1224), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT62), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1139), .A2(new_n967), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1210), .A2(new_n1176), .A3(new_n1237), .A4(new_n1177), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1216), .A2(G213), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G375), .B2(G378), .ZN(new_n1241));
  INV_X1    g1041(.A(G384), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1018), .B1(new_n1182), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1080), .A2(KEYINPUT60), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1186), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1208), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1242), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1184), .A2(new_n1185), .B1(new_n1080), .B2(KEYINPUT60), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G384), .B(new_n1208), .C1(new_n1249), .C2(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1236), .B1(new_n1241), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1210), .B1(new_n1145), .B2(new_n1179), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1254), .A2(KEYINPUT62), .A3(new_n1240), .A4(new_n1251), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1216), .A2(G213), .A3(G2897), .ZN(new_n1257));
  AOI211_X1 g1057(.A(KEYINPUT126), .B(new_n1257), .C1(new_n1248), .C2(new_n1250), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1257), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1259), .B1(new_n1251), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1251), .A2(new_n1260), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1258), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1254), .B2(new_n1240), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1235), .B1(new_n1256), .B2(new_n1266), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1264), .A2(KEYINPUT63), .B1(new_n1241), .B2(new_n1252), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1240), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1131), .A2(new_n1134), .A3(new_n1018), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1134), .B1(new_n1131), .B2(new_n1018), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1144), .A2(new_n1140), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1178), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1269), .B(new_n1252), .C1(new_n1274), .C2(new_n1210), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1235), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1268), .A2(new_n1277), .A3(KEYINPUT61), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1219), .B1(new_n1267), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(KEYINPUT62), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1241), .A2(new_n1236), .A3(new_n1252), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1265), .A4(new_n1264), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1235), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1277), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1264), .A2(KEYINPUT63), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1275), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1287), .A3(new_n1265), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1284), .A2(new_n1288), .A3(KEYINPUT127), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1279), .A2(new_n1289), .ZN(G405));
  NOR2_X1   g1090(.A1(new_n1211), .A2(new_n1254), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1252), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1283), .ZN(G402));
endmodule


