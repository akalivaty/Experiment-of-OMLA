

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(n730), .ZN(n705) );
  OR2_X1 U555 ( .A1(n709), .A2(n708), .ZN(n712) );
  OR2_X1 U556 ( .A1(n759), .A2(n758), .ZN(n765) );
  NOR2_X1 U557 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U558 ( .A1(n805), .A2(n814), .ZN(n806) );
  AND2_X1 U559 ( .A1(n605), .A2(G2105), .ZN(n882) );
  NOR2_X1 U560 ( .A1(G651), .A2(n653), .ZN(n648) );
  NAND2_X1 U561 ( .A1(G2104), .A2(G101), .ZN(n522) );
  NOR2_X1 U562 ( .A1(G2105), .A2(n522), .ZN(n523) );
  XNOR2_X1 U563 ( .A(KEYINPUT23), .B(n523), .ZN(n525) );
  INV_X1 U564 ( .A(G2104), .ZN(n605) );
  NAND2_X1 U565 ( .A1(n882), .A2(G125), .ZN(n524) );
  NAND2_X1 U566 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U567 ( .A(KEYINPUT64), .B(n526), .ZN(n532) );
  XNOR2_X1 U568 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n528) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X2 U570 ( .A(n528), .B(n527), .ZN(n876) );
  NAND2_X1 U571 ( .A1(n876), .A2(G137), .ZN(n530) );
  AND2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U573 ( .A1(n880), .A2(G113), .ZN(n529) );
  NAND2_X1 U574 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U575 ( .A1(n532), .A2(n531), .ZN(G160) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n639) );
  NAND2_X1 U577 ( .A1(G90), .A2(n639), .ZN(n534) );
  XOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  INV_X1 U579 ( .A(G651), .ZN(n536) );
  NOR2_X1 U580 ( .A1(n653), .A2(n536), .ZN(n642) );
  NAND2_X1 U581 ( .A1(G77), .A2(n642), .ZN(n533) );
  NAND2_X1 U582 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U583 ( .A(n535), .B(KEYINPUT9), .ZN(n539) );
  NOR2_X1 U584 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n537), .Z(n652) );
  NAND2_X1 U586 ( .A1(G64), .A2(n652), .ZN(n538) );
  NAND2_X1 U587 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U588 ( .A1(G52), .A2(n648), .ZN(n540) );
  XNOR2_X1 U589 ( .A(KEYINPUT67), .B(n540), .ZN(n541) );
  NOR2_X1 U590 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U591 ( .A(KEYINPUT68), .B(n543), .ZN(G171) );
  INV_X1 U592 ( .A(G171), .ZN(G301) );
  XOR2_X1 U593 ( .A(G2446), .B(G2430), .Z(n545) );
  XNOR2_X1 U594 ( .A(G2451), .B(KEYINPUT96), .ZN(n544) );
  XNOR2_X1 U595 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U596 ( .A(n546), .B(G2427), .Z(n548) );
  XNOR2_X1 U597 ( .A(G1341), .B(G1348), .ZN(n547) );
  XNOR2_X1 U598 ( .A(n548), .B(n547), .ZN(n552) );
  XOR2_X1 U599 ( .A(G2443), .B(G2435), .Z(n550) );
  XNOR2_X1 U600 ( .A(G2438), .B(G2454), .ZN(n549) );
  XNOR2_X1 U601 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U602 ( .A(n552), .B(n551), .Z(n553) );
  AND2_X1 U603 ( .A1(G14), .A2(n553), .ZN(G401) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U605 ( .A(G132), .ZN(G219) );
  INV_X1 U606 ( .A(G82), .ZN(G220) );
  INV_X1 U607 ( .A(G57), .ZN(G237) );
  NAND2_X1 U608 ( .A1(n648), .A2(G51), .ZN(n554) );
  XOR2_X1 U609 ( .A(KEYINPUT71), .B(n554), .Z(n556) );
  NAND2_X1 U610 ( .A1(n652), .A2(G63), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U612 ( .A(KEYINPUT6), .B(n557), .ZN(n564) );
  NAND2_X1 U613 ( .A1(n639), .A2(G89), .ZN(n558) );
  XNOR2_X1 U614 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G76), .A2(n642), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U617 ( .A(KEYINPUT5), .B(n561), .Z(n562) );
  XNOR2_X1 U618 ( .A(KEYINPUT70), .B(n562), .ZN(n563) );
  NOR2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(n565), .Z(G168) );
  XOR2_X1 U621 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U623 ( .A(n566), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U624 ( .A(G223), .ZN(n824) );
  NAND2_X1 U625 ( .A1(n824), .A2(G567), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U627 ( .A1(G56), .A2(n652), .ZN(n568) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n568), .Z(n574) );
  NAND2_X1 U629 ( .A1(n639), .A2(G81), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G68), .A2(n642), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT13), .B(n572), .Z(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n648), .A2(G43), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n968) );
  INV_X1 U637 ( .A(G860), .ZN(n595) );
  OR2_X1 U638 ( .A1(n968), .A2(n595), .ZN(G153) );
  NAND2_X1 U639 ( .A1(G301), .A2(G868), .ZN(n585) );
  NAND2_X1 U640 ( .A1(G79), .A2(n642), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G54), .A2(n648), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G92), .A2(n639), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G66), .A2(n652), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT15), .ZN(n969) );
  INV_X1 U648 ( .A(G868), .ZN(n666) );
  NAND2_X1 U649 ( .A1(n969), .A2(n666), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G78), .A2(n642), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G53), .A2(n648), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G91), .A2(n639), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G65), .A2(n652), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n592), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U659 ( .A1(G286), .A2(G868), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G299), .A2(n666), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U662 ( .A1(G559), .A2(n595), .ZN(n596) );
  XNOR2_X1 U663 ( .A(KEYINPUT72), .B(n596), .ZN(n597) );
  INV_X1 U664 ( .A(n969), .ZN(n612) );
  NAND2_X1 U665 ( .A1(n597), .A2(n612), .ZN(n598) );
  XNOR2_X1 U666 ( .A(KEYINPUT16), .B(n598), .ZN(G148) );
  NOR2_X1 U667 ( .A1(G868), .A2(n968), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G868), .A2(n612), .ZN(n599) );
  NOR2_X1 U669 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U671 ( .A1(G123), .A2(n882), .ZN(n602) );
  XNOR2_X1 U672 ( .A(n602), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n880), .A2(G111), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G135), .A2(n876), .ZN(n607) );
  NOR2_X1 U676 ( .A1(G2105), .A2(n605), .ZN(n877) );
  NAND2_X1 U677 ( .A1(G99), .A2(n877), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n911) );
  XNOR2_X1 U680 ( .A(G2096), .B(n911), .ZN(n611) );
  INV_X1 U681 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U683 ( .A1(G559), .A2(n612), .ZN(n613) );
  XOR2_X1 U684 ( .A(n968), .B(n613), .Z(n664) );
  XNOR2_X1 U685 ( .A(KEYINPUT73), .B(n664), .ZN(n614) );
  NOR2_X1 U686 ( .A1(G860), .A2(n614), .ZN(n615) );
  XNOR2_X1 U687 ( .A(n615), .B(KEYINPUT75), .ZN(n623) );
  NAND2_X1 U688 ( .A1(G93), .A2(n639), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G67), .A2(n652), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n642), .A2(G80), .ZN(n618) );
  XOR2_X1 U692 ( .A(KEYINPUT74), .B(n618), .Z(n619) );
  NOR2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n648), .A2(G55), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n667) );
  XNOR2_X1 U696 ( .A(n623), .B(n667), .ZN(G145) );
  NAND2_X1 U697 ( .A1(G50), .A2(n648), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G62), .A2(n652), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U700 ( .A(KEYINPUT77), .B(n626), .ZN(n630) );
  NAND2_X1 U701 ( .A1(G88), .A2(n639), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G75), .A2(n642), .ZN(n627) );
  AND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(G303) );
  INV_X1 U705 ( .A(G303), .ZN(G166) );
  NAND2_X1 U706 ( .A1(G86), .A2(n639), .ZN(n632) );
  NAND2_X1 U707 ( .A1(G61), .A2(n652), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n642), .A2(G73), .ZN(n633) );
  XOR2_X1 U710 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(KEYINPUT76), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G48), .A2(n648), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U715 ( .A1(G85), .A2(n639), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G60), .A2(n652), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G72), .A2(n642), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G47), .A2(n648), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U722 ( .A(KEYINPUT66), .B(n647), .Z(G290) );
  NAND2_X1 U723 ( .A1(G49), .A2(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(G288) );
  XNOR2_X1 U729 ( .A(G166), .B(G305), .ZN(n663) );
  XOR2_X1 U730 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n656) );
  XNOR2_X1 U731 ( .A(G288), .B(n656), .ZN(n657) );
  XOR2_X1 U732 ( .A(n657), .B(KEYINPUT19), .Z(n659) );
  INV_X1 U733 ( .A(G299), .ZN(n972) );
  XNOR2_X1 U734 ( .A(n972), .B(KEYINPUT79), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U736 ( .A(G290), .B(n660), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n661), .B(n667), .ZN(n662) );
  XNOR2_X1 U738 ( .A(n663), .B(n662), .ZN(n898) );
  XOR2_X1 U739 ( .A(n898), .B(n664), .Z(n665) );
  NOR2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n669) );
  NOR2_X1 U741 ( .A1(G868), .A2(n667), .ZN(n668) );
  NOR2_X1 U742 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n671), .ZN(n673) );
  XOR2_X1 U746 ( .A(KEYINPUT21), .B(KEYINPUT81), .Z(n672) );
  XNOR2_X1 U747 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U748 ( .A1(G2072), .A2(n674), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U750 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U751 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U752 ( .A1(G108), .A2(n676), .ZN(n833) );
  NAND2_X1 U753 ( .A1(n833), .A2(G567), .ZN(n682) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U756 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U757 ( .A1(G96), .A2(n679), .ZN(n832) );
  NAND2_X1 U758 ( .A1(G2106), .A2(n832), .ZN(n680) );
  XNOR2_X1 U759 ( .A(KEYINPUT82), .B(n680), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n834) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U762 ( .A1(n834), .A2(n683), .ZN(n831) );
  NAND2_X1 U763 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U764 ( .A1(n876), .A2(G138), .ZN(n686) );
  NAND2_X1 U765 ( .A1(G114), .A2(n880), .ZN(n684) );
  XOR2_X1 U766 ( .A(KEYINPUT83), .B(n684), .Z(n685) );
  NAND2_X1 U767 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U768 ( .A1(G126), .A2(n882), .ZN(n688) );
  NAND2_X1 U769 ( .A1(G102), .A2(n877), .ZN(n687) );
  NAND2_X1 U770 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U771 ( .A1(n690), .A2(n689), .ZN(G164) );
  NAND2_X1 U772 ( .A1(G40), .A2(G160), .ZN(n691) );
  XNOR2_X1 U773 ( .A(n691), .B(KEYINPUT84), .ZN(n773) );
  INV_X1 U774 ( .A(KEYINPUT90), .ZN(n692) );
  XNOR2_X1 U775 ( .A(n773), .B(n692), .ZN(n693) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n772) );
  NAND2_X2 U777 ( .A1(n693), .A2(n772), .ZN(n730) );
  OR2_X1 U778 ( .A1(n705), .A2(G1961), .ZN(n695) );
  XNOR2_X1 U779 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NAND2_X1 U780 ( .A1(n705), .A2(n943), .ZN(n694) );
  NAND2_X1 U781 ( .A1(n695), .A2(n694), .ZN(n723) );
  NAND2_X1 U782 ( .A1(n723), .A2(G171), .ZN(n722) );
  NAND2_X1 U783 ( .A1(G1956), .A2(n730), .ZN(n696) );
  XNOR2_X1 U784 ( .A(KEYINPUT91), .B(n696), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n705), .A2(G2072), .ZN(n697) );
  XNOR2_X1 U786 ( .A(KEYINPUT27), .B(n697), .ZN(n698) );
  NOR2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n715) );
  NAND2_X1 U788 ( .A1(n972), .A2(n715), .ZN(n714) );
  AND2_X1 U789 ( .A1(n705), .A2(G1996), .ZN(n700) );
  XNOR2_X1 U790 ( .A(n700), .B(KEYINPUT26), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n730), .A2(G1341), .ZN(n702) );
  INV_X1 U792 ( .A(n968), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n709) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n730), .ZN(n707) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n705), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n969), .A2(n710), .ZN(n708) );
  NAND2_X1 U799 ( .A1(n969), .A2(n710), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n719) );
  NOR2_X1 U802 ( .A1(n972), .A2(n715), .ZN(n717) );
  INV_X1 U803 ( .A(KEYINPUT28), .ZN(n716) );
  XNOR2_X1 U804 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U806 ( .A(KEYINPUT29), .B(n720), .Z(n721) );
  NAND2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n743) );
  NOR2_X1 U808 ( .A1(G171), .A2(n723), .ZN(n728) );
  NAND2_X2 U809 ( .A1(G8), .A2(n730), .ZN(n768) );
  NOR2_X1 U810 ( .A1(G1966), .A2(n768), .ZN(n745) );
  NOR2_X1 U811 ( .A1(G2084), .A2(n730), .ZN(n741) );
  NOR2_X1 U812 ( .A1(n745), .A2(n741), .ZN(n724) );
  NAND2_X1 U813 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U814 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U815 ( .A1(G168), .A2(n726), .ZN(n727) );
  XOR2_X1 U816 ( .A(KEYINPUT31), .B(n729), .Z(n742) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n768), .ZN(n732) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U820 ( .A1(n733), .A2(G303), .ZN(n735) );
  AND2_X1 U821 ( .A1(n742), .A2(n735), .ZN(n734) );
  NAND2_X1 U822 ( .A1(n743), .A2(n734), .ZN(n738) );
  INV_X1 U823 ( .A(n735), .ZN(n736) );
  OR2_X1 U824 ( .A1(n736), .A2(G286), .ZN(n737) );
  AND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n739), .A2(G8), .ZN(n740) );
  XNOR2_X1 U827 ( .A(n740), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U828 ( .A1(G8), .A2(n741), .ZN(n747) );
  AND2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U831 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U832 ( .A1(n749), .A2(n748), .ZN(n762) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n755) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U835 ( .A1(n755), .A2(n750), .ZN(n976) );
  NAND2_X1 U836 ( .A1(n762), .A2(n976), .ZN(n753) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n975) );
  INV_X1 U838 ( .A(n975), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n751), .A2(n768), .ZN(n752) );
  AND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U841 ( .A1(n754), .A2(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U842 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  OR2_X1 U843 ( .A1(n756), .A2(n768), .ZN(n757) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n965) );
  NAND2_X1 U845 ( .A1(n757), .A2(n965), .ZN(n758) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U849 ( .A1(n763), .A2(n768), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n765), .A2(n764), .ZN(n770) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XOR2_X1 U852 ( .A(n766), .B(KEYINPUT24), .Z(n767) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U854 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U855 ( .A(KEYINPUT92), .B(n771), .Z(n807) );
  NOR2_X1 U856 ( .A1(n773), .A2(n772), .ZN(n819) );
  XNOR2_X1 U857 ( .A(G290), .B(G1986), .ZN(n981) );
  NAND2_X1 U858 ( .A1(n819), .A2(n981), .ZN(n774) );
  XNOR2_X1 U859 ( .A(KEYINPUT85), .B(n774), .ZN(n792) );
  NAND2_X1 U860 ( .A1(G117), .A2(n880), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G141), .A2(n876), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U863 ( .A1(n877), .A2(G105), .ZN(n777) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(n777), .Z(n778) );
  NOR2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U866 ( .A1(n882), .A2(G129), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n871) );
  NAND2_X1 U868 ( .A1(G1996), .A2(n871), .ZN(n790) );
  NAND2_X1 U869 ( .A1(G119), .A2(n882), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G95), .A2(n877), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G107), .A2(n880), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G131), .A2(n876), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U876 ( .A(n788), .B(KEYINPUT89), .ZN(n892) );
  NAND2_X1 U877 ( .A1(G1991), .A2(n892), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n912) );
  AND2_X1 U879 ( .A1(n912), .A2(n819), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n805) );
  XNOR2_X1 U881 ( .A(KEYINPUT37), .B(G2067), .ZN(n816) );
  NAND2_X1 U882 ( .A1(n880), .A2(G116), .ZN(n793) );
  XOR2_X1 U883 ( .A(KEYINPUT87), .B(n793), .Z(n795) );
  NAND2_X1 U884 ( .A1(n882), .A2(G128), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U886 ( .A(KEYINPUT35), .B(n796), .Z(n802) );
  NAND2_X1 U887 ( .A1(G140), .A2(n876), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G104), .A2(n877), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U890 ( .A(KEYINPUT34), .B(n799), .ZN(n800) );
  XNOR2_X1 U891 ( .A(KEYINPUT86), .B(n800), .ZN(n801) );
  NOR2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n803), .ZN(n895) );
  NOR2_X1 U894 ( .A1(n816), .A2(n895), .ZN(n921) );
  NAND2_X1 U895 ( .A1(n819), .A2(n921), .ZN(n804) );
  XNOR2_X1 U896 ( .A(n804), .B(KEYINPUT88), .ZN(n814) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n822) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n871), .ZN(n808) );
  XOR2_X1 U899 ( .A(KEYINPUT93), .B(n808), .Z(n925) );
  NOR2_X1 U900 ( .A1(G1991), .A2(n892), .ZN(n913) );
  NOR2_X1 U901 ( .A1(G290), .A2(G1986), .ZN(n809) );
  XNOR2_X1 U902 ( .A(KEYINPUT94), .B(n809), .ZN(n810) );
  NOR2_X1 U903 ( .A1(n913), .A2(n810), .ZN(n811) );
  NOR2_X1 U904 ( .A1(n912), .A2(n811), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n925), .A2(n812), .ZN(n813) );
  XNOR2_X1 U906 ( .A(n813), .B(KEYINPUT39), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n816), .A2(n895), .ZN(n922) );
  NAND2_X1 U909 ( .A1(n817), .A2(n922), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U911 ( .A(KEYINPUT95), .B(n820), .Z(n821) );
  NAND2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U913 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U914 ( .A1(n824), .A2(G2106), .ZN(n825) );
  XOR2_X1 U915 ( .A(KEYINPUT97), .B(n825), .Z(G217) );
  INV_X1 U916 ( .A(G661), .ZN(n827) );
  NAND2_X1 U917 ( .A1(G2), .A2(G15), .ZN(n826) );
  NOR2_X1 U918 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT98), .B(n828), .Z(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n829) );
  XOR2_X1 U921 ( .A(KEYINPUT99), .B(n829), .Z(n830) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  NOR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  INV_X1 U929 ( .A(n834), .ZN(G319) );
  XOR2_X1 U930 ( .A(G2096), .B(KEYINPUT43), .Z(n836) );
  XNOR2_X1 U931 ( .A(G2072), .B(G2678), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U933 ( .A(n837), .B(KEYINPUT42), .Z(n839) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2090), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U936 ( .A(KEYINPUT100), .B(G2100), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2084), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U940 ( .A(G1986), .B(G1976), .Z(n845) );
  XNOR2_X1 U941 ( .A(G1961), .B(G1971), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U943 ( .A(G1991), .B(G1981), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1996), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U946 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U947 ( .A(KEYINPUT101), .B(G2474), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U949 ( .A(G1956), .B(KEYINPUT41), .Z(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U951 ( .A1(G124), .A2(n882), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n854), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U953 ( .A1(G112), .A2(n880), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n855), .B(KEYINPUT102), .ZN(n856) );
  NAND2_X1 U955 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U956 ( .A1(G136), .A2(n876), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G100), .A2(n877), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U959 ( .A1(n861), .A2(n860), .ZN(G162) );
  NAND2_X1 U960 ( .A1(G118), .A2(n880), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G130), .A2(n882), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U963 ( .A1(G142), .A2(n876), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G106), .A2(n877), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(KEYINPUT45), .B(n866), .ZN(n867) );
  XNOR2_X1 U967 ( .A(KEYINPUT103), .B(n867), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n891) );
  XOR2_X1 U969 ( .A(G164), .B(n911), .Z(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U971 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n873) );
  XNOR2_X1 U972 ( .A(KEYINPUT106), .B(KEYINPUT105), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U974 ( .A(n875), .B(n874), .Z(n889) );
  NAND2_X1 U975 ( .A1(G139), .A2(n876), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G103), .A2(n877), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n887) );
  NAND2_X1 U978 ( .A1(n880), .A2(G115), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n881), .B(KEYINPUT104), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n916) );
  XNOR2_X1 U984 ( .A(G160), .B(n916), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n892), .B(G162), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G286), .B(n898), .ZN(n901) );
  XNOR2_X1 U992 ( .A(KEYINPUT107), .B(n968), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n899), .B(n969), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U995 ( .A(n902), .B(G301), .ZN(n903) );
  NOR2_X1 U996 ( .A1(G37), .A2(n903), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n904) );
  XOR2_X1 U998 ( .A(KEYINPUT49), .B(n904), .Z(n905) );
  NAND2_X1 U999 ( .A1(G319), .A2(n905), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G401), .A2(n906), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(KEYINPUT108), .B(n907), .ZN(n909) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1006 ( .A(G160), .B(G2084), .Z(n910) );
  NOR2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(n934) );
  XOR2_X1 U1010 ( .A(n916), .B(KEYINPUT111), .Z(n917) );
  XOR2_X1 U1011 ( .A(G2072), .B(n917), .Z(n919) );
  XOR2_X1 U1012 ( .A(G164), .B(G2078), .Z(n918) );
  NOR2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(KEYINPUT50), .B(n920), .ZN(n932) );
  INV_X1 U1015 ( .A(n921), .ZN(n923) );
  NAND2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(n930) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n926), .Z(n928) );
  XNOR2_X1 U1020 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(n928), .B(n927), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1024 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1025 ( .A(KEYINPUT52), .B(n935), .Z(n936) );
  NOR2_X1 U1026 ( .A1(KEYINPUT55), .A2(n936), .ZN(n937) );
  XOR2_X1 U1027 ( .A(KEYINPUT112), .B(n937), .Z(n938) );
  NAND2_X1 U1028 ( .A1(n938), .A2(G29), .ZN(n939) );
  XOR2_X1 U1029 ( .A(KEYINPUT113), .B(n939), .Z(n1025) );
  XNOR2_X1 U1030 ( .A(G2084), .B(G34), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(n940), .B(KEYINPUT54), .ZN(n960) );
  XNOR2_X1 U1032 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1033 ( .A(KEYINPUT115), .B(G2067), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(G26), .ZN(n950) );
  XNOR2_X1 U1035 ( .A(G2072), .B(G33), .ZN(n948) );
  XNOR2_X1 U1036 ( .A(G1996), .B(G32), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n942), .B(KEYINPUT116), .ZN(n945) );
  XOR2_X1 U1038 ( .A(G27), .B(n943), .Z(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(n946), .B(KEYINPUT117), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1043 ( .A(G1991), .B(G25), .Z(n951) );
  NAND2_X1 U1044 ( .A1(n951), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(KEYINPUT114), .B(n952), .ZN(n953) );
  NOR2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1049 ( .A(KEYINPUT118), .B(n958), .Z(n959) );
  NOR2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(KEYINPUT55), .B(n961), .ZN(n963) );
  INV_X1 U1052 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1054 ( .A1(n964), .A2(G11), .ZN(n1023) );
  XNOR2_X1 U1055 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G168), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(KEYINPUT57), .B(n967), .ZN(n989) );
  XNOR2_X1 U1059 ( .A(n968), .B(G1341), .ZN(n971) );
  XNOR2_X1 U1060 ( .A(n969), .B(G1348), .ZN(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n986) );
  XNOR2_X1 U1062 ( .A(n972), .B(G1956), .ZN(n974) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n978) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(n979), .B(KEYINPUT119), .ZN(n980) );
  NOR2_X1 U1068 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1069 ( .A(KEYINPUT120), .B(n982), .Z(n984) );
  XNOR2_X1 U1070 ( .A(G301), .B(G1961), .ZN(n983) );
  NOR2_X1 U1071 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1072 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1073 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1075 ( .A1(n991), .A2(n990), .ZN(n1021) );
  INV_X1 U1076 ( .A(G16), .ZN(n1019) );
  XNOR2_X1 U1077 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n1017) );
  XOR2_X1 U1078 ( .A(G1956), .B(G20), .Z(n996) );
  XNOR2_X1 U1079 ( .A(G1341), .B(G19), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1981), .B(G6), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n994), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1084 ( .A(KEYINPUT59), .B(G1348), .Z(n997) );
  XNOR2_X1 U1085 ( .A(G4), .B(n997), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(n1000), .B(KEYINPUT123), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1001), .B(KEYINPUT60), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(G21), .B(G1966), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(KEYINPUT124), .B(n1004), .Z(n1006) );
  XNOR2_X1 U1092 ( .A(G1961), .B(G5), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT125), .B(n1007), .Z(n1015) );
  XOR2_X1 U1095 ( .A(G1971), .B(G22), .Z(n1010) );
  XOR2_X1 U1096 ( .A(G24), .B(KEYINPUT126), .Z(n1008) );
  XNOR2_X1 U1097 ( .A(n1008), .B(G1986), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

