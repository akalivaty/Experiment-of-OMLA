//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1301, new_n1302, new_n1303,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT64), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g0020(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n206), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n217), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n216), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n246), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G274), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n256), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n259), .A2(G226), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G222), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n263), .B1(new_n208), .B2(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n222), .A2(new_n252), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI211_X1 g0068(.A(new_n257), .B(new_n260), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G179), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT68), .ZN(new_n272));
  OAI21_X1  g0072(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G150), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n224), .A2(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n273), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n220), .A2(new_n221), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n278), .A2(new_n280), .B1(new_n201), .B2(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n220), .A2(new_n281), .A3(new_n221), .A4(new_n279), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n224), .A2(G1), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(G50), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n269), .B2(G169), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n272), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n269), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G190), .B2(new_n269), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n283), .A2(KEYINPUT69), .A3(new_n288), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n294), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n294), .B(new_n303), .C1(new_n300), .C2(new_n299), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n291), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n254), .ZN(new_n306));
  INV_X1    g0106(.A(new_n256), .ZN(new_n307));
  AOI22_X1  g0107(.A1(G232), .A2(new_n259), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  MUX2_X1   g0108(.A(G223), .B(G226), .S(G1698), .Z(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(G33), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT3), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n309), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G87), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n308), .B(G179), .C1(new_n319), .C2(new_n267), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n259), .A2(G232), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n306), .A2(new_n307), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n267), .B1(new_n317), .B2(new_n318), .ZN(new_n324));
  OAI21_X1  g0124(.A(G169), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G68), .ZN(new_n327));
  AOI21_X1  g0127(.A(G20), .B1(new_n314), .B2(new_n316), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n329), .ZN(new_n332));
  INV_X1    g0132(.A(new_n316), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n336), .B2(G33), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n332), .B1(new_n337), .B2(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n202), .A2(new_n327), .ZN(new_n340));
  NOR2_X1   g0140(.A1(G58), .A2(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(G20), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n274), .A2(G159), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n339), .A2(KEYINPUT16), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT16), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n315), .B1(new_n334), .B2(new_n335), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n311), .A2(G33), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(G20), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n261), .B2(G20), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n327), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n347), .B1(new_n355), .B2(new_n344), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n346), .A2(new_n280), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n277), .A2(new_n286), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n277), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n359), .A2(new_n284), .B1(new_n281), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n326), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n280), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n344), .B1(new_n330), .B2(new_n338), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(KEYINPUT16), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n361), .B1(new_n368), .B2(new_n356), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT18), .B1(new_n369), .B2(new_n326), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n308), .B(G190), .C1(new_n319), .C2(new_n267), .ZN(new_n372));
  OAI21_X1  g0172(.A(G200), .B1(new_n323), .B2(new_n324), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n357), .A2(new_n374), .A3(new_n362), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n369), .A2(KEYINPUT17), .A3(new_n374), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n261), .A2(G232), .A3(new_n262), .ZN(new_n381));
  INV_X1    g0181(.A(G238), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n381), .B1(new_n210), .B2(new_n261), .C1(new_n264), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n268), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n322), .B1(new_n209), .B2(new_n258), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G200), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n385), .B1(new_n268), .B2(new_n383), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G190), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n284), .A2(new_n208), .A3(new_n286), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n281), .A2(G77), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n360), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n276), .B2(new_n394), .ZN(new_n395));
  AOI211_X1 g0195(.A(new_n391), .B(new_n392), .C1(new_n395), .C2(new_n280), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n389), .A2(new_n270), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n392), .B1(new_n395), .B2(new_n280), .ZN(new_n399));
  INV_X1    g0199(.A(new_n391), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n398), .B(new_n401), .C1(G169), .C2(new_n389), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n305), .A2(new_n380), .A3(new_n397), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n316), .A2(new_n349), .A3(G226), .A4(new_n262), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT70), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT70), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n261), .A2(new_n407), .A3(G226), .A4(new_n262), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n316), .A2(new_n349), .A3(G232), .A4(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n267), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n322), .B1(new_n382), .B2(new_n258), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT13), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n257), .B1(G238), .B2(new_n259), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n412), .B1(new_n408), .B2(new_n406), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n417), .B(new_n418), .C1(new_n419), .C2(new_n267), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n404), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT14), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n416), .A2(new_n420), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n421), .A2(new_n422), .B1(new_n423), .B2(new_n270), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n422), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT71), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(KEYINPUT71), .A3(new_n422), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n327), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n208), .B2(new_n276), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n280), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT11), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n284), .A2(new_n327), .A3(new_n286), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n281), .A2(G68), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT12), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n433), .B2(new_n432), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n429), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G190), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n423), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n292), .B1(new_n416), .B2(new_n420), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OR3_X1    g0247(.A1(new_n403), .A2(new_n447), .A3(KEYINPUT74), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT74), .B1(new_n403), .B2(new_n447), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(G238), .A2(G1698), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n209), .B2(G1698), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n314), .A3(new_n316), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n315), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n267), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n253), .B(G250), .C1(G1), .C2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(G1), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n253), .A2(G274), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G190), .ZN(new_n464));
  OAI21_X1  g0264(.A(G200), .B1(new_n457), .B2(new_n462), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  INV_X1    g0266(.A(G87), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n466), .A2(new_n467), .B1(new_n411), .B2(new_n224), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT19), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G97), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n468), .A2(new_n469), .B1(new_n276), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n314), .A2(new_n224), .A3(G68), .A4(new_n316), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n366), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n394), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n281), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n315), .A2(G1), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n284), .A2(new_n467), .A3(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n464), .A2(new_n465), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n462), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n455), .B1(new_n337), .B2(new_n452), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n270), .B(new_n480), .C1(new_n481), .C2(new_n267), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n404), .B1(new_n457), .B2(new_n462), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n284), .A2(new_n394), .A3(new_n476), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n473), .A2(new_n475), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT78), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n482), .B(new_n483), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n475), .ZN(new_n488));
  INV_X1    g0288(.A(new_n484), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n471), .A2(new_n472), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n488), .B(new_n489), .C1(new_n490), .C2(new_n366), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(KEYINPUT78), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n479), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(KEYINPUT79), .B(new_n479), .C1(new_n487), .C2(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n284), .A2(new_n476), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT25), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n281), .B2(G107), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n282), .A2(KEYINPUT25), .A3(new_n210), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n498), .A2(G107), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT22), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n467), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n314), .A2(new_n224), .A3(new_n316), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n316), .A2(new_n349), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n224), .A2(G87), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT23), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n224), .B2(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n210), .A2(KEYINPUT23), .A3(G20), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n510), .A2(new_n511), .B1(new_n455), .B2(new_n224), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n505), .A2(new_n508), .A3(new_n515), .A4(new_n512), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n514), .A2(KEYINPUT24), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n280), .B1(new_n514), .B2(KEYINPUT24), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n502), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  NOR2_X1   g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n460), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n522), .A2(G264), .A3(new_n253), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G250), .A2(G1698), .ZN(new_n524));
  INV_X1    g0324(.A(G257), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G1698), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(new_n314), .A3(new_n316), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G294), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n523), .B1(new_n529), .B2(new_n268), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT5), .B(G41), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(new_n253), .A3(G274), .A4(new_n460), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n404), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n267), .B1(new_n527), .B2(new_n528), .ZN(new_n534));
  INV_X1    g0334(.A(new_n532), .ZN(new_n535));
  NOR4_X1   g0335(.A1(new_n534), .A2(new_n270), .A3(new_n523), .A4(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT86), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n530), .A2(G179), .A3(new_n532), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT86), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n534), .A2(new_n535), .A3(new_n523), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n538), .B(new_n539), .C1(new_n404), .C2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n519), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n514), .A2(KEYINPUT24), .A3(new_n516), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n543), .B(new_n280), .C1(KEYINPUT24), .C2(new_n514), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(G190), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n530), .A2(new_n532), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n544), .A2(new_n502), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n209), .A2(G1698), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT4), .B1(new_n337), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT76), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(G33), .A3(G283), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n268), .B1(new_n550), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n522), .A2(new_n253), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n532), .B1(new_n561), .B2(new_n525), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT77), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT77), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n532), .B(new_n564), .C1(new_n561), .C2(new_n525), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n498), .A2(G97), .ZN(new_n568));
  INV_X1    g0368(.A(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n282), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n352), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n348), .B2(new_n349), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT7), .B1(new_n506), .B2(new_n224), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g0375(.A(G97), .B(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(KEYINPUT75), .B2(KEYINPUT6), .ZN(new_n577));
  NOR2_X1   g0377(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(KEYINPUT6), .B2(new_n569), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n577), .B(G20), .C1(new_n576), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n274), .A2(G77), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n571), .B1(new_n582), .B2(new_n280), .ZN(new_n583));
  INV_X1    g0383(.A(new_n562), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n559), .A2(G190), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n567), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n583), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n563), .A2(new_n565), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n588), .A2(new_n270), .A3(new_n559), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n404), .B1(new_n560), .B2(new_n562), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n542), .A2(new_n548), .A3(new_n586), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(KEYINPUT84), .A2(KEYINPUT21), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT81), .B1(new_n498), .B2(G116), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT81), .ZN(new_n595));
  NOR4_X1   g0395(.A1(new_n284), .A2(new_n595), .A3(new_n454), .A4(new_n476), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n594), .A2(new_n596), .B1(G116), .B2(new_n281), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n454), .A2(G20), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n280), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n224), .B1(new_n569), .B2(G33), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n556), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n600), .A2(KEYINPUT82), .A3(KEYINPUT20), .A4(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT20), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n601), .B1(new_n553), .B2(new_n555), .ZN(new_n606));
  OAI211_X1 g0406(.A(KEYINPUT83), .B(new_n605), .C1(new_n599), .C2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n605), .B1(new_n599), .B2(new_n606), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT83), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n603), .A2(KEYINPUT20), .A3(new_n280), .A4(new_n598), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT82), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n609), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n597), .B1(new_n608), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n314), .A2(new_n316), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n211), .A2(G1698), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(G257), .B2(G1698), .ZN(new_n617));
  INV_X1    g0417(.A(G303), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n615), .A2(new_n617), .B1(new_n618), .B2(new_n261), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n268), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n522), .A2(G270), .A3(new_n253), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(KEYINPUT80), .A3(new_n532), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT80), .B1(new_n621), .B2(new_n532), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G169), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n593), .B1(new_n614), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n284), .A2(new_n476), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n595), .B1(new_n628), .B2(new_n454), .ZN(new_n629));
  INV_X1    g0429(.A(new_n596), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n629), .A2(new_n630), .B1(new_n454), .B2(new_n282), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n609), .A2(new_n610), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n611), .A2(new_n612), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n604), .A4(new_n607), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n620), .B(G179), .C1(new_n623), .C2(new_n624), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n624), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n622), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n404), .B1(new_n640), .B2(new_n620), .ZN(new_n641));
  INV_X1    g0441(.A(new_n593), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n635), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n625), .A2(G200), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n640), .A2(G190), .A3(new_n620), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n634), .A4(new_n631), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n627), .A2(new_n638), .A3(new_n643), .A4(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n497), .A2(new_n592), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n450), .A2(new_n648), .ZN(G372));
  AND3_X1   g0449(.A1(new_n459), .A2(KEYINPUT87), .A3(new_n461), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT87), .B1(new_n459), .B2(new_n461), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n650), .A2(new_n651), .B1(new_n481), .B2(new_n267), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n404), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n491), .A3(new_n482), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(G200), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n464), .A3(new_n478), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n654), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n591), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n519), .B1(new_n533), .B2(new_n536), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n627), .A2(new_n662), .A3(new_n638), .A4(new_n643), .ZN(new_n663));
  INV_X1    g0463(.A(new_n658), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n664), .A2(new_n548), .A3(new_n591), .A4(new_n586), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n661), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n496), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n482), .A2(new_n483), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n491), .A2(KEYINPUT78), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n485), .A2(new_n486), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT79), .B1(new_n672), .B2(new_n479), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n591), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n660), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n450), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n365), .A2(new_n370), .A3(KEYINPUT88), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT88), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n369), .A2(KEYINPUT18), .A3(new_n326), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n357), .A2(new_n362), .ZN(new_n683));
  INV_X1    g0483(.A(new_n326), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n364), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n681), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n445), .ZN(new_n687));
  INV_X1    g0487(.A(new_n402), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n441), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n680), .B(new_n686), .C1(new_n689), .C2(new_n379), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n302), .A2(new_n304), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n291), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n679), .A2(new_n692), .ZN(G369));
  NAND3_X1  g0493(.A1(new_n627), .A2(new_n638), .A3(new_n643), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n255), .A2(new_n224), .A3(G13), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G213), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n614), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n647), .B2(new_n702), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n542), .A2(new_n548), .ZN(new_n707));
  INV_X1    g0507(.A(new_n519), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n701), .ZN(new_n709));
  OAI22_X1  g0509(.A1(new_n707), .A2(new_n709), .B1(new_n542), .B2(new_n701), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n694), .A2(new_n701), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n707), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n662), .A2(new_n700), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n229), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n466), .A2(new_n467), .A3(new_n454), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n226), .B2(new_n719), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT89), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n559), .A2(new_n463), .A3(new_n530), .A4(new_n584), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  OR3_X1    g0527(.A1(new_n726), .A2(new_n727), .A3(new_n636), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n726), .B2(new_n636), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n546), .A2(new_n270), .A3(new_n652), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n625), .B1(new_n560), .B2(new_n566), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n733));
  NOR2_X1   g0533(.A1(new_n701), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT91), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n588), .A2(new_n559), .B1(new_n640), .B2(new_n620), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n546), .A2(new_n270), .A3(new_n652), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n731), .A2(new_n730), .A3(KEYINPUT91), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n728), .A2(new_n729), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n701), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n735), .B1(new_n743), .B2(KEYINPUT31), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT92), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n648), .B2(new_n701), .ZN(new_n747));
  AND4_X1   g0547(.A1(new_n542), .A2(new_n548), .A3(new_n591), .A4(new_n586), .ZN(new_n748));
  AND4_X1   g0548(.A1(new_n627), .A2(new_n638), .A3(new_n643), .A4(new_n646), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n674), .A3(new_n749), .A4(new_n701), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(KEYINPUT92), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n745), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT93), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n750), .A2(KEYINPUT92), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n497), .A2(new_n592), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n756), .A2(new_n746), .A3(new_n749), .A4(new_n701), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n744), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G330), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT93), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(KEYINPUT29), .B(new_n700), .C1(new_n667), .C2(new_n677), .ZN(new_n763));
  INV_X1    g0563(.A(new_n542), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n694), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n654), .B1(new_n765), .B2(new_n665), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n658), .A2(new_n591), .A3(new_n660), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n495), .A2(new_n496), .A3(new_n675), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(new_n768), .B2(new_n660), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n701), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(KEYINPUT29), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n763), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n725), .B1(new_n774), .B2(G1), .ZN(G364));
  XNOR2_X1  g0575(.A(new_n705), .B(KEYINPUT94), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n224), .A2(G13), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n255), .B1(new_n777), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OR3_X1    g0579(.A1(new_n779), .A2(new_n718), .A3(KEYINPUT95), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT95), .B1(new_n779), .B2(new_n718), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n776), .B(new_n782), .C1(G330), .C2(new_n704), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n223), .B1(G20), .B2(new_n404), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n246), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT97), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n337), .A2(new_n717), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n458), .B2(new_n227), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n790), .A2(G45), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n791), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n261), .A2(new_n229), .ZN(new_n797));
  INV_X1    g0597(.A(G355), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(KEYINPUT96), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(new_n800), .B1(new_n454), .B2(new_n717), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n789), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n784), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n224), .A2(G179), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(new_n442), .A3(G200), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n261), .B1(new_n805), .B2(new_n210), .C1(new_n467), .C2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT99), .Z(new_n808));
  NOR2_X1   g0608(.A1(G190), .A2(G200), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G159), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT32), .ZN(new_n813));
  NAND2_X1  g0613(.A1(G20), .A2(G179), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G190), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n813), .B1(G68), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n814), .A2(new_n442), .A3(G200), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n815), .A2(new_n809), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n820), .A2(new_n202), .B1(new_n821), .B2(new_n208), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT98), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n816), .A2(new_n442), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n442), .A2(G179), .A3(G200), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n224), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n826), .A2(new_n201), .B1(new_n569), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n823), .B2(new_n822), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n808), .A2(new_n818), .A3(new_n824), .A4(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n810), .A2(KEYINPUT100), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n810), .A2(KEYINPUT100), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G329), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n828), .A2(new_n837), .B1(new_n805), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT33), .B(G317), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n817), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G322), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n506), .B1(new_n820), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n821), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(G311), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n806), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G326), .A2(new_n825), .B1(new_n846), .B2(G303), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n836), .A2(new_n841), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n803), .B1(new_n831), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n802), .A2(new_n849), .A3(new_n782), .ZN(new_n850));
  INV_X1    g0650(.A(new_n787), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n704), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n783), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT101), .ZN(G396));
  NOR2_X1   g0654(.A1(new_n784), .A2(new_n785), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n782), .B1(new_n855), .B2(new_n208), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n844), .A2(G159), .B1(G143), .B2(new_n819), .ZN(new_n857));
  INV_X1    g0657(.A(new_n817), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n857), .B1(new_n858), .B2(new_n859), .C1(new_n860), .C2(new_n826), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT34), .ZN(new_n862));
  INV_X1    g0662(.A(new_n805), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n846), .A2(G50), .B1(new_n863), .B2(G68), .ZN(new_n864));
  INV_X1    g0664(.A(new_n828), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n615), .B1(new_n865), .B2(G58), .ZN(new_n866));
  INV_X1    g0666(.A(G132), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n864), .B(new_n866), .C1(new_n834), .C2(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n862), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n835), .A2(G311), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n467), .A2(new_n805), .B1(new_n806), .B2(new_n210), .ZN(new_n873));
  XOR2_X1   g0673(.A(KEYINPUT102), .B(G283), .Z(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n817), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n506), .B1(new_n821), .B2(new_n454), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G294), .B2(new_n819), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n865), .A2(G97), .B1(new_n825), .B2(G303), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n872), .A2(new_n876), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n387), .A2(new_n404), .B1(new_n399), .B2(new_n400), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n398), .A3(new_n701), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n401), .A2(new_n700), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n397), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n882), .B(new_n884), .C1(new_n886), .C2(new_n688), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n397), .A2(new_n885), .B1(new_n883), .B2(new_n398), .ZN(new_n888));
  INV_X1    g0688(.A(new_n884), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT104), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n856), .B1(new_n803), .B2(new_n881), .C1(new_n891), .C2(new_n786), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n678), .B2(new_n701), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n891), .B(new_n701), .C1(new_n666), .C2(new_n676), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n761), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n782), .B1(new_n761), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(G384));
  OAI21_X1  g0699(.A(new_n577), .B1(new_n576), .B2(new_n579), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT105), .Z(new_n901));
  OR2_X1    g0701(.A1(new_n901), .A2(KEYINPUT35), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(KEYINPUT35), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(G116), .A4(new_n225), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT36), .Z(new_n905));
  OAI211_X1 g0705(.A(new_n227), .B(G77), .C1(new_n202), .C2(new_n327), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n201), .A2(G68), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n255), .B(G13), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n894), .A2(new_n884), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n367), .A2(KEYINPUT16), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n361), .B1(new_n911), .B2(new_n368), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n375), .B1(new_n912), .B2(new_n698), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n326), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n363), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n698), .B1(new_n357), .B2(new_n362), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT37), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n375), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n912), .A2(new_n698), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n371), .B2(new_n379), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n921), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n440), .ZN(new_n929));
  INV_X1    g0729(.A(new_n424), .ZN(new_n930));
  INV_X1    g0730(.A(new_n428), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT71), .B1(new_n421), .B2(new_n422), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n929), .B(new_n700), .C1(new_n933), .C2(new_n445), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n929), .A2(new_n700), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n687), .B(new_n935), .C1(new_n429), .C2(new_n440), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n910), .A2(new_n928), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n686), .A2(new_n680), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n698), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(KEYINPUT106), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n441), .A2(new_n701), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n944));
  INV_X1    g0744(.A(new_n927), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n686), .A2(new_n377), .A3(new_n680), .A4(new_n378), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n917), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n916), .A2(new_n918), .A3(new_n375), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n357), .A2(new_n362), .A3(new_n374), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n949), .A2(new_n917), .A3(new_n681), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n948), .B1(new_n950), .B2(new_n919), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n949), .A2(new_n917), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n952), .A2(new_n681), .A3(KEYINPUT37), .A4(new_n916), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n945), .B1(new_n955), .B2(new_n925), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n943), .B(new_n944), .C1(new_n956), .C2(KEYINPUT39), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n941), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT106), .B1(new_n938), .B2(new_n940), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n450), .B1(new_n771), .B2(new_n763), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n692), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n960), .B(new_n962), .Z(new_n963));
  INV_X1    g0763(.A(KEYINPUT40), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n937), .A2(new_n891), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n755), .A2(new_n757), .ZN(new_n966));
  INV_X1    g0766(.A(new_n733), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n743), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(KEYINPUT31), .B2(new_n743), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n965), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n951), .A2(new_n953), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n917), .B2(new_n946), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n927), .B1(new_n972), .B2(KEYINPUT38), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n964), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n969), .A2(new_n966), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT40), .B1(new_n926), .B2(new_n927), .ZN(new_n976));
  INV_X1    g0776(.A(new_n965), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n450), .A2(new_n975), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n759), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n980), .B2(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n963), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n255), .B2(new_n777), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n963), .A2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n909), .B1(new_n984), .B2(new_n985), .ZN(G367));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n591), .A2(new_n586), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n587), .A2(new_n700), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n988), .A2(new_n989), .B1(new_n675), .B2(new_n700), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT107), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n987), .B1(new_n991), .B2(new_n715), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT110), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n990), .B(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n715), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT109), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT110), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n987), .C1(new_n991), .C2(new_n715), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT109), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n995), .A2(new_n996), .A3(new_n1001), .A4(KEYINPUT44), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n993), .A2(new_n998), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n995), .A2(new_n996), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n711), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1003), .A2(new_n1005), .A3(new_n711), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n713), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n712), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1011), .B1(new_n710), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(new_n705), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n776), .B2(new_n1013), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n774), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT111), .B1(new_n1010), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1015), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n773), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT111), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1019), .A2(new_n1020), .A3(new_n1009), .A4(new_n1008), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n773), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n718), .B(KEYINPUT41), .Z(new_n1023));
  OAI21_X1  g0823(.A(new_n778), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n591), .B1(new_n995), .B2(new_n542), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT108), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n701), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n995), .A2(new_n1011), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT42), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n478), .A2(new_n701), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n664), .A2(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n654), .A2(new_n1032), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1029), .A2(new_n1031), .B1(KEYINPUT43), .B2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(KEYINPUT43), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n711), .A2(new_n995), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1024), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n788), .B1(new_n229), .B2(new_n394), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n241), .B2(new_n792), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n820), .A2(new_n859), .B1(new_n810), .B2(new_n860), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n506), .B(new_n1044), .C1(G50), .C2(new_n844), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n865), .A2(G68), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G159), .A2(new_n817), .B1(new_n846), .B2(G58), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G143), .A2(new_n825), .B1(new_n863), .B2(G77), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n828), .A2(new_n210), .B1(new_n805), .B2(new_n569), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G311), .B2(new_n825), .ZN(new_n1051));
  INV_X1    g0851(.A(G317), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n820), .A2(new_n618), .B1(new_n810), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n844), .B2(new_n875), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n846), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n337), .B1(G294), .B2(new_n817), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT46), .B1(new_n846), .B2(G116), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT112), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n1049), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n782), .B(new_n1043), .C1(new_n1062), .C2(new_n784), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1033), .A2(new_n787), .A3(new_n1034), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1041), .A2(new_n1065), .ZN(G387));
  NAND2_X1  g0866(.A1(new_n773), .A2(new_n1018), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1016), .A2(new_n718), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT116), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n782), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n797), .A2(new_n721), .B1(G107), .B2(new_n229), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n238), .A2(G45), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n277), .A2(G50), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT50), .ZN(new_n1074));
  AOI211_X1 g0874(.A(G45), .B(new_n720), .C1(G68), .C2(G77), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n793), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1071), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1070), .B1(new_n1077), .B2(new_n789), .ZN(new_n1078));
  INV_X1    g0878(.A(G159), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n826), .A2(new_n1079), .B1(new_n394), .B2(new_n828), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n844), .A2(G68), .B1(G50), .B2(new_n819), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n859), .B2(new_n810), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n858), .A2(new_n277), .B1(new_n806), .B2(new_n208), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n337), .B1(new_n569), .B2(new_n805), .ZN(new_n1084));
  NOR4_X1   g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT114), .Z(new_n1086));
  AOI21_X1  g0886(.A(new_n337), .B1(G326), .B2(new_n811), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n828), .A2(new_n874), .B1(new_n806), .B2(new_n837), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n844), .A2(G303), .B1(G317), .B2(new_n819), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n817), .A2(G311), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(new_n842), .C2(new_n826), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT48), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1092), .B2(new_n1091), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT49), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1087), .B1(new_n454), .B2(new_n805), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1086), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1078), .B1(new_n1098), .B2(new_n784), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n710), .B2(new_n851), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT115), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1015), .B2(new_n779), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1068), .A2(new_n1069), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1067), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n718), .B1(new_n773), .B2(new_n1018), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT116), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1103), .A2(new_n1107), .ZN(G393));
  NAND2_X1  g0908(.A1(new_n995), .A2(new_n787), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n789), .B1(G97), .B2(new_n717), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n250), .A2(new_n792), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n825), .A2(G317), .B1(G311), .B2(new_n819), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT52), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n506), .B1(new_n821), .B2(new_n837), .C1(new_n842), .C2(new_n810), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n858), .A2(new_n618), .B1(new_n805), .B2(new_n210), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n828), .A2(new_n454), .B1(new_n874), .B2(new_n806), .ZN(new_n1117));
  OR4_X1    g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n828), .A2(new_n208), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G87), .B2(new_n863), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n201), .B2(new_n858), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n615), .B(new_n1123), .C1(new_n360), .C2(new_n844), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n825), .A2(G150), .B1(G159), .B2(new_n819), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT51), .Z(new_n1126));
  AOI22_X1  g0926(.A1(new_n846), .A2(G68), .B1(new_n811), .B2(G143), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT117), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1120), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n782), .B(new_n1112), .C1(new_n1131), .C2(new_n784), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1109), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1010), .B2(new_n778), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n719), .B1(new_n1010), .B2(new_n1016), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(G390));
  NAND3_X1  g0938(.A1(new_n975), .A2(new_n977), .A3(G330), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT120), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT38), .B1(new_n947), .B2(new_n954), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n942), .B1(new_n1142), .B2(new_n945), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n937), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n891), .B(new_n701), .C1(new_n766), .C2(new_n769), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n884), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT119), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n884), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n937), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT119), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1149), .A2(new_n973), .A3(new_n1150), .A4(new_n942), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n910), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n942), .B1(new_n1153), .B2(new_n1144), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n944), .B1(new_n956), .B2(KEYINPUT39), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1141), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n891), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n754), .B2(new_n760), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(new_n937), .C1(KEYINPUT120), .C2(new_n1139), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1157), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1155), .A2(new_n785), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n855), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1070), .B1(new_n360), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n805), .A2(new_n201), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n858), .A2(new_n860), .B1(new_n1079), .B2(new_n828), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(G128), .C2(new_n825), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n835), .A2(G125), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n821), .A2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n506), .B(new_n1172), .C1(G132), .C2(new_n819), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n806), .A2(new_n859), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1169), .A2(new_n1170), .A3(new_n1173), .A4(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n834), .A2(new_n837), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n506), .B1(new_n821), .B2(new_n569), .C1(new_n820), .C2(new_n454), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n327), .A2(new_n805), .B1(new_n806), .B2(new_n467), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1121), .B1(G107), .B2(new_n817), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n838), .C2(new_n826), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT122), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(new_n803), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1177), .A2(KEYINPUT122), .A3(new_n1183), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1166), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1163), .A2(new_n779), .B1(new_n1164), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n450), .A2(G330), .A3(new_n975), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n961), .A2(new_n1189), .A3(new_n692), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1139), .B1(new_n1161), .B2(new_n937), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n910), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n761), .A2(new_n891), .A3(new_n937), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n975), .A2(G330), .A3(new_n891), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1148), .B1(new_n1194), .B2(new_n1144), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1190), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n718), .B1(new_n1163), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n753), .B1(new_n752), .B2(G330), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n758), .A2(KEYINPUT93), .A3(new_n759), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n891), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1140), .B1(new_n1201), .B2(new_n1144), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1196), .B1(new_n1202), .B2(new_n1153), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1190), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1141), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1158), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1162), .A2(new_n1152), .A3(new_n1156), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1188), .B1(new_n1198), .B2(new_n1210), .ZN(G378));
  OAI21_X1  g1011(.A(G330), .B1(new_n974), .B2(new_n978), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n305), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n698), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n298), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n305), .A2(new_n1215), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  OR3_X1    g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1212), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1223), .B(G330), .C1(new_n974), .C2(new_n978), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n960), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1225), .A2(new_n960), .A3(new_n1226), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1224), .A2(new_n785), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1070), .B1(G50), .B2(new_n1165), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n835), .A2(G283), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n337), .A2(G41), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n844), .A2(new_n474), .B1(G107), .B2(new_n819), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1234), .A2(new_n1046), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n826), .A2(new_n454), .B1(new_n806), .B2(new_n208), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n863), .A2(G58), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n858), .B2(new_n569), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT58), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1235), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n825), .A2(G125), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n858), .B2(new_n867), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n844), .A2(G137), .B1(G128), .B2(new_n819), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n806), .B2(new_n1171), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1247), .B(new_n1249), .C1(G150), .C2(new_n865), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(KEYINPUT59), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(KEYINPUT59), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n863), .A2(G159), .ZN(new_n1254));
  AOI211_X1 g1054(.A(G33), .B(G41), .C1(new_n811), .C2(G124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1245), .B1(KEYINPUT58), .B2(new_n1241), .C1(new_n1252), .C2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1233), .B1(new_n1257), .B2(new_n784), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1231), .A2(new_n779), .B1(new_n1232), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1190), .B1(new_n1163), .B2(new_n1197), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1225), .A2(new_n960), .A3(new_n1226), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n960), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT57), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n718), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1191), .A2(new_n910), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1204), .B1(new_n1209), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT57), .B1(new_n1266), .B2(new_n1231), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1259), .B1(new_n1264), .B2(new_n1267), .ZN(G375));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1190), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1023), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1205), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1070), .B1(G68), .B2(new_n1165), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n826), .A2(new_n837), .B1(new_n806), .B2(new_n569), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G116), .B2(new_n817), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n835), .A2(G303), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n506), .B1(new_n821), .B2(new_n210), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(G283), .B2(new_n819), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n865), .A2(new_n474), .B1(new_n863), .B2(G77), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1274), .A2(new_n1275), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n337), .B1(new_n859), .B2(new_n821), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1239), .B1(new_n1079), .B2(new_n806), .C1(new_n201), .C2(new_n828), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(G128), .C2(new_n835), .ZN(new_n1282));
  XOR2_X1   g1082(.A(new_n1282), .B(KEYINPUT123), .Z(new_n1283));
  NAND2_X1  g1083(.A1(new_n825), .A2(G132), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1284), .B1(new_n860), .B2(new_n820), .C1(new_n858), .C2(new_n1171), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1279), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1272), .B1(new_n1286), .B2(new_n784), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n937), .B2(new_n786), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1271), .B(new_n1288), .C1(new_n778), .C2(new_n1265), .ZN(G381));
  INV_X1    g1089(.A(G375), .ZN(new_n1290));
  INV_X1    g1090(.A(G387), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1164), .A2(new_n1187), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1209), .B2(new_n778), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n719), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1163), .A2(new_n1197), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G396), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1103), .A2(new_n1107), .A3(new_n1297), .ZN(new_n1298));
  NOR4_X1   g1098(.A1(G390), .A2(G381), .A3(new_n1298), .A4(G384), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1290), .A2(new_n1291), .A3(new_n1296), .A4(new_n1299), .ZN(G407));
  INV_X1    g1100(.A(G213), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(G343), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1296), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G407), .B(G213), .C1(G375), .C2(new_n1303), .ZN(G409));
  NAND2_X1  g1104(.A1(G387), .A2(KEYINPUT127), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1041), .A2(new_n1306), .A3(new_n1065), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1297), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(G390), .A2(new_n1309), .A3(new_n1298), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1298), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1137), .B1(new_n1311), .B2(new_n1308), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1305), .A2(new_n1307), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1306), .B1(new_n1041), .B2(new_n1065), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1065), .ZN(new_n1316));
  AOI211_X1 g1116(.A(KEYINPUT127), .B(new_n1316), .C1(new_n1024), .C2(new_n1040), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1314), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1313), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G378), .B(new_n1259), .C1(new_n1264), .C2(new_n1267), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1266), .A2(new_n1270), .A3(new_n1231), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1259), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1296), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1302), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT60), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1269), .B1(new_n1197), .B2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1265), .A2(KEYINPUT60), .A3(new_n1190), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n718), .A3(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT124), .ZN(new_n1330));
  OAI221_X1 g1130(.A(new_n1288), .B1(G384), .B2(new_n1330), .C1(new_n1265), .C2(new_n778), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G384), .A2(new_n1330), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1329), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1333), .B1(new_n1329), .B2(new_n1332), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT125), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1335), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1326), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n718), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1328), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1332), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1333), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT125), .B1(new_n1345), .B2(new_n1334), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1325), .B1(new_n1338), .B2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(KEYINPUT62), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT62), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1325), .B(new_n1349), .C1(new_n1338), .C2(new_n1346), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT61), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1302), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1302), .A2(G2897), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1345), .A2(new_n1357), .A3(new_n1334), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1337), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1345), .A2(KEYINPUT125), .A3(new_n1334), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1357), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1352), .B1(new_n1359), .B2(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1320), .B1(new_n1351), .B2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1347), .A2(KEYINPUT63), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT63), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1325), .B(new_n1366), .C1(new_n1338), .C2(new_n1346), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1365), .A2(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(KEYINPUT61), .B1(new_n1313), .B2(new_n1318), .ZN(new_n1369));
  OAI21_X1  g1169(.A(KEYINPUT126), .B1(new_n1359), .B2(new_n1362), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1356), .B1(new_n1338), .B2(new_n1346), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT126), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1371), .A2(new_n1372), .A3(new_n1355), .A4(new_n1358), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1368), .A2(new_n1369), .A3(new_n1370), .A4(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1364), .A2(new_n1374), .ZN(G405));
  NAND2_X1  g1175(.A1(G375), .A2(new_n1296), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1376), .A2(new_n1321), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1377), .A2(new_n1361), .A3(new_n1360), .ZN(new_n1378));
  OAI211_X1 g1178(.A(new_n1376), .B(new_n1321), .C1(new_n1336), .C2(new_n1335), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1380));
  XNOR2_X1  g1180(.A(new_n1319), .B(new_n1380), .ZN(G402));
endmodule


