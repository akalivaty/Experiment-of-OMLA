

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594;

  NOR2_X1 U326 ( .A1(n589), .A2(n393), .ZN(n394) );
  XNOR2_X1 U327 ( .A(n454), .B(n453), .ZN(n455) );
  OR2_X1 U328 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U329 ( .A(n331), .B(n330), .ZN(n334) );
  XNOR2_X1 U330 ( .A(n329), .B(n328), .ZN(n330) );
  NOR2_X1 U331 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U332 ( .A(n490), .B(KEYINPUT107), .ZN(n491) );
  XNOR2_X1 U333 ( .A(n456), .B(n455), .ZN(n459) );
  XOR2_X1 U334 ( .A(G211GAT), .B(G78GAT), .Z(n294) );
  XOR2_X1 U335 ( .A(n449), .B(n448), .Z(n295) );
  XOR2_X1 U336 ( .A(n349), .B(n348), .Z(n296) );
  XOR2_X1 U337 ( .A(G1GAT), .B(G64GAT), .Z(n297) );
  XNOR2_X1 U338 ( .A(n338), .B(n297), .ZN(n341) );
  XNOR2_X1 U339 ( .A(n341), .B(n340), .ZN(n343) );
  XOR2_X1 U340 ( .A(G50GAT), .B(G162GAT), .Z(n438) );
  INV_X1 U341 ( .A(KEYINPUT87), .ZN(n453) );
  AND2_X1 U342 ( .A1(n578), .A2(n479), .ZN(n447) );
  INV_X1 U343 ( .A(KEYINPUT37), .ZN(n490) );
  XNOR2_X1 U344 ( .A(n492), .B(n491), .ZN(n534) );
  XOR2_X1 U345 ( .A(n336), .B(n335), .Z(n556) );
  XNOR2_X1 U346 ( .A(n461), .B(n460), .ZN(n544) );
  XNOR2_X1 U347 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U348 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U349 ( .A(n472), .B(n471), .ZN(G1349GAT) );
  XNOR2_X1 U350 ( .A(n498), .B(n497), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(G8GAT), .B(KEYINPUT81), .Z(n338) );
  XOR2_X1 U352 ( .A(G211GAT), .B(KEYINPUT21), .Z(n299) );
  XNOR2_X1 U353 ( .A(G197GAT), .B(G218GAT), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n435) );
  XOR2_X1 U355 ( .A(n338), .B(n435), .Z(n301) );
  NAND2_X1 U356 ( .A1(G226GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(G176GAT), .B(G64GAT), .Z(n360) );
  XOR2_X1 U359 ( .A(n302), .B(n360), .Z(n304) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G92GAT), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n314) );
  XOR2_X1 U362 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n306) );
  XNOR2_X1 U363 ( .A(G190GAT), .B(KEYINPUT89), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U365 ( .A(n307), .B(KEYINPUT17), .Z(n309) );
  XNOR2_X1 U366 ( .A(G169GAT), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n461) );
  XOR2_X1 U368 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n311) );
  XNOR2_X1 U369 ( .A(G204GAT), .B(KEYINPUT101), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U371 ( .A(n461), .B(n312), .Z(n313) );
  XOR2_X1 U372 ( .A(n314), .B(n313), .Z(n537) );
  INV_X1 U373 ( .A(n537), .ZN(n399) );
  INV_X1 U374 ( .A(KEYINPUT36), .ZN(n337) );
  XOR2_X1 U375 ( .A(KEYINPUT10), .B(KEYINPUT78), .Z(n316) );
  XNOR2_X1 U376 ( .A(G99GAT), .B(KEYINPUT9), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U378 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n318) );
  XNOR2_X1 U379 ( .A(G190GAT), .B(G106GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n336) );
  XOR2_X1 U382 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n322) );
  XNOR2_X1 U383 ( .A(G36GAT), .B(G29GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U385 ( .A(KEYINPUT7), .B(n323), .Z(n389) );
  INV_X1 U386 ( .A(n389), .ZN(n327) );
  XOR2_X1 U387 ( .A(KEYINPUT79), .B(n438), .Z(n325) );
  XOR2_X1 U388 ( .A(G43GAT), .B(G134GAT), .Z(n449) );
  XNOR2_X1 U389 ( .A(n449), .B(G218GAT), .ZN(n324) );
  XNOR2_X1 U390 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n331) );
  NAND2_X1 U392 ( .A1(G232GAT), .A2(G233GAT), .ZN(n329) );
  INV_X1 U393 ( .A(KEYINPUT65), .ZN(n328) );
  XNOR2_X1 U394 ( .A(G85GAT), .B(G92GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n332), .B(KEYINPUT74), .ZN(n368) );
  XNOR2_X1 U396 ( .A(KEYINPUT80), .B(n368), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n337), .B(n556), .ZN(n488) );
  XNOR2_X1 U399 ( .A(G183GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n294), .B(n339), .ZN(n340) );
  XNOR2_X1 U401 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n342), .B(KEYINPUT13), .ZN(n359) );
  XOR2_X1 U403 ( .A(n343), .B(n359), .Z(n345) );
  XOR2_X1 U404 ( .A(G15GAT), .B(G127GAT), .Z(n457) );
  XOR2_X1 U405 ( .A(G22GAT), .B(G155GAT), .Z(n432) );
  XNOR2_X1 U406 ( .A(n457), .B(n432), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U408 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n347) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U411 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n351) );
  XNOR2_X1 U412 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n352), .B(KEYINPUT15), .ZN(n353) );
  XOR2_X1 U415 ( .A(n296), .B(n353), .Z(n570) );
  NOR2_X1 U416 ( .A1(n488), .A2(n570), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n354), .B(KEYINPUT45), .ZN(n391) );
  XNOR2_X1 U418 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n355), .B(KEYINPUT73), .ZN(n356) );
  XOR2_X1 U420 ( .A(n356), .B(G204GAT), .Z(n358) );
  XNOR2_X1 U421 ( .A(G78GAT), .B(G106GAT), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n443) );
  XOR2_X1 U423 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n362) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n443), .B(n363), .ZN(n372) );
  XOR2_X1 U427 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n365) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U430 ( .A(n366), .B(KEYINPUT33), .Z(n370) );
  XNOR2_X1 U431 ( .A(G99GAT), .B(G71GAT), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n367), .B(G120GAT), .ZN(n452) );
  XNOR2_X1 U433 ( .A(n452), .B(n368), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U435 ( .A(n372), .B(n371), .Z(n586) );
  XOR2_X1 U436 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n374) );
  XNOR2_X1 U437 ( .A(G8GAT), .B(KEYINPUT67), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n387) );
  XOR2_X1 U439 ( .A(G22GAT), .B(G197GAT), .Z(n376) );
  XNOR2_X1 U440 ( .A(G43GAT), .B(G50GAT), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U442 ( .A(G113GAT), .B(G15GAT), .Z(n378) );
  XNOR2_X1 U443 ( .A(G169GAT), .B(G141GAT), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U445 ( .A(n380), .B(n379), .Z(n385) );
  XOR2_X1 U446 ( .A(KEYINPUT68), .B(G1GAT), .Z(n382) );
  NAND2_X1 U447 ( .A1(G229GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U449 ( .A(KEYINPUT70), .B(n383), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U451 ( .A(n387), .B(n386), .Z(n388) );
  XOR2_X1 U452 ( .A(n389), .B(n388), .Z(n581) );
  INV_X1 U453 ( .A(n581), .ZN(n564) );
  AND2_X1 U454 ( .A1(n586), .A2(n564), .ZN(n390) );
  AND2_X1 U455 ( .A1(n391), .A2(n390), .ZN(n397) );
  INV_X1 U456 ( .A(n556), .ZN(n574) );
  INV_X1 U457 ( .A(n570), .ZN(n589) );
  XOR2_X1 U458 ( .A(n586), .B(KEYINPUT41), .Z(n566) );
  NOR2_X1 U459 ( .A1(n564), .A2(n566), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n392), .B(KEYINPUT46), .ZN(n393) );
  NAND2_X1 U461 ( .A1(n574), .A2(n394), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n395), .B(KEYINPUT47), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n398), .B(KEYINPUT48), .ZN(n561) );
  NOR2_X1 U464 ( .A1(n399), .A2(n561), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n400), .B(KEYINPUT54), .ZN(n427) );
  XOR2_X1 U466 ( .A(G85GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U467 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n401), .B(KEYINPUT86), .ZN(n448) );
  XNOR2_X1 U469 ( .A(G134GAT), .B(n448), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U471 ( .A(G29GAT), .B(n404), .ZN(n426) );
  XOR2_X1 U472 ( .A(KEYINPUT98), .B(KEYINPUT1), .Z(n406) );
  XNOR2_X1 U473 ( .A(KEYINPUT97), .B(KEYINPUT6), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U475 ( .A(KEYINPUT96), .B(n407), .Z(n409) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U478 ( .A(n410), .B(KEYINPUT4), .Z(n416) );
  XOR2_X1 U479 ( .A(KEYINPUT93), .B(KEYINPUT2), .Z(n412) );
  XNOR2_X1 U480 ( .A(KEYINPUT3), .B(KEYINPUT94), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U482 ( .A(G141GAT), .B(n413), .Z(n444) );
  INV_X1 U483 ( .A(n444), .ZN(n414) );
  XOR2_X1 U484 ( .A(n414), .B(KEYINPUT5), .Z(n415) );
  XNOR2_X1 U485 ( .A(n416), .B(n415), .ZN(n424) );
  XOR2_X1 U486 ( .A(KEYINPUT95), .B(G57GAT), .Z(n418) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(G127GAT), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U489 ( .A(KEYINPUT80), .B(G155GAT), .Z(n420) );
  XNOR2_X1 U490 ( .A(G120GAT), .B(G148GAT), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U492 ( .A(n422), .B(n421), .Z(n423) );
  XNOR2_X1 U493 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U494 ( .A(n426), .B(n425), .Z(n507) );
  NAND2_X1 U495 ( .A1(n427), .A2(n507), .ZN(n429) );
  INV_X1 U496 ( .A(KEYINPUT64), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n429), .B(n428), .ZN(n578) );
  XOR2_X1 U498 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n431) );
  XNOR2_X1 U499 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n430) );
  XNOR2_X1 U500 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U501 ( .A(n433), .B(n432), .Z(n441) );
  INV_X1 U502 ( .A(KEYINPUT91), .ZN(n434) );
  XNOR2_X1 U503 ( .A(n435), .B(n434), .ZN(n437) );
  NAND2_X1 U504 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U505 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U506 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U507 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U508 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U509 ( .A(n445), .B(n444), .Z(n479) );
  XNOR2_X1 U510 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n446) );
  XNOR2_X1 U511 ( .A(n447), .B(n446), .ZN(n463) );
  NAND2_X1 U512 ( .A1(G227GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n295), .B(n450), .ZN(n451) );
  XOR2_X1 U514 ( .A(n451), .B(G176GAT), .Z(n456) );
  XNOR2_X1 U515 ( .A(n452), .B(KEYINPUT88), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT20), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U518 ( .A(n544), .ZN(n462) );
  XNOR2_X2 U519 ( .A(n464), .B(KEYINPUT119), .ZN(n576) );
  NAND2_X1 U520 ( .A1(n576), .A2(n581), .ZN(n466) );
  XNOR2_X1 U521 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(G1348GAT) );
  XNOR2_X1 U523 ( .A(KEYINPUT111), .B(n566), .ZN(n549) );
  NAND2_X1 U524 ( .A1(n549), .A2(n576), .ZN(n472) );
  XOR2_X1 U525 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n468) );
  XNOR2_X1 U526 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n467) );
  XOR2_X1 U527 ( .A(n468), .B(n467), .Z(n470) );
  XOR2_X1 U528 ( .A(G176GAT), .B(KEYINPUT56), .Z(n469) );
  NOR2_X1 U529 ( .A1(n544), .A2(n479), .ZN(n473) );
  XNOR2_X1 U530 ( .A(KEYINPUT26), .B(n473), .ZN(n579) );
  XOR2_X1 U531 ( .A(KEYINPUT27), .B(n537), .Z(n482) );
  INV_X1 U532 ( .A(n482), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n579), .A2(n474), .ZN(n560) );
  NAND2_X1 U534 ( .A1(n537), .A2(n544), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n479), .A2(n475), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT25), .B(n476), .Z(n477) );
  NAND2_X1 U537 ( .A1(n560), .A2(n477), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n478), .A2(n507), .ZN(n486) );
  XOR2_X1 U539 ( .A(n544), .B(KEYINPUT90), .Z(n483) );
  XNOR2_X1 U540 ( .A(KEYINPUT66), .B(KEYINPUT28), .ZN(n480) );
  XOR2_X1 U541 ( .A(n480), .B(n479), .Z(n540) );
  OR2_X1 U542 ( .A1(n507), .A2(n540), .ZN(n481) );
  NOR2_X1 U543 ( .A1(n482), .A2(n481), .ZN(n545) );
  NAND2_X1 U544 ( .A1(n483), .A2(n545), .ZN(n484) );
  XNOR2_X1 U545 ( .A(KEYINPUT102), .B(n484), .ZN(n485) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT103), .B(n487), .Z(n504) );
  NOR2_X1 U548 ( .A1(n589), .A2(n488), .ZN(n489) );
  AND2_X1 U549 ( .A1(n504), .A2(n489), .ZN(n492) );
  NAND2_X1 U550 ( .A1(n581), .A2(n586), .ZN(n506) );
  NOR2_X1 U551 ( .A1(n534), .A2(n506), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT108), .B(KEYINPUT38), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n522) );
  NAND2_X1 U554 ( .A1(n522), .A2(n544), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n496) );
  INV_X1 U556 ( .A(G43GAT), .ZN(n495) );
  NAND2_X1 U557 ( .A1(n576), .A2(n556), .ZN(n500) );
  XOR2_X1 U558 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n502) );
  INV_X1 U560 ( .A(G190GAT), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1351GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT34), .Z(n509) );
  NOR2_X1 U563 ( .A1(n556), .A2(n570), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT16), .ZN(n505) );
  NAND2_X1 U565 ( .A1(n505), .A2(n504), .ZN(n524) );
  NOR2_X1 U566 ( .A1(n506), .A2(n524), .ZN(n516) );
  INV_X1 U567 ( .A(n507), .ZN(n562) );
  NAND2_X1 U568 ( .A1(n516), .A2(n562), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U570 ( .A(G1GAT), .B(n510), .Z(G1324GAT) );
  NAND2_X1 U571 ( .A1(n516), .A2(n537), .ZN(n511) );
  XNOR2_X1 U572 ( .A(n511), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT35), .Z(n513) );
  NAND2_X1 U574 ( .A1(n516), .A2(n544), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(n515) );
  XOR2_X1 U576 ( .A(G15GAT), .B(KEYINPUT105), .Z(n514) );
  XNOR2_X1 U577 ( .A(n515), .B(n514), .ZN(G1326GAT) );
  NAND2_X1 U578 ( .A1(n516), .A2(n540), .ZN(n517) );
  XNOR2_X1 U579 ( .A(n517), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U580 ( .A1(n562), .A2(n522), .ZN(n520) );
  XNOR2_X1 U581 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1328GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n537), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U586 ( .A1(n522), .A2(n540), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U588 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n526) );
  NAND2_X1 U589 ( .A1(n549), .A2(n564), .ZN(n533) );
  NOR2_X1 U590 ( .A1(n533), .A2(n524), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n530), .A2(n562), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1332GAT) );
  NAND2_X1 U593 ( .A1(n530), .A2(n537), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U595 ( .A1(n544), .A2(n530), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(KEYINPUT112), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G71GAT), .B(n529), .ZN(G1334GAT) );
  XOR2_X1 U598 ( .A(G78GAT), .B(KEYINPUT43), .Z(n532) );
  NAND2_X1 U599 ( .A1(n530), .A2(n540), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(G1335GAT) );
  XOR2_X1 U601 ( .A(G85GAT), .B(KEYINPUT113), .Z(n536) );
  NOR2_X1 U602 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n541), .A2(n562), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1336GAT) );
  NAND2_X1 U605 ( .A1(n541), .A2(n537), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n538), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U607 ( .A1(n544), .A2(n541), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n539), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(KEYINPUT44), .ZN(n543) );
  XNOR2_X1 U611 ( .A(G106GAT), .B(n543), .ZN(G1339GAT) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U613 ( .A1(n561), .A2(n546), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n557), .A2(n581), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT114), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G113GAT), .B(n548), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n551) );
  NAND2_X1 U618 ( .A1(n557), .A2(n549), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U620 ( .A(G120GAT), .B(n552), .Z(G1341GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n554) );
  NAND2_X1 U622 ( .A1(n557), .A2(n589), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U624 ( .A(G127GAT), .B(n555), .Z(G1342GAT) );
  XOR2_X1 U625 ( .A(G134GAT), .B(KEYINPUT51), .Z(n559) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1343GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n573) );
  NOR2_X1 U630 ( .A1(n564), .A2(n573), .ZN(n565) );
  XOR2_X1 U631 ( .A(G141GAT), .B(n565), .Z(G1344GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n573), .ZN(n568) );
  XNOR2_X1 U633 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G148GAT), .B(n569), .ZN(G1345GAT) );
  NOR2_X1 U636 ( .A1(n570), .A2(n573), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1346GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G162GAT), .B(n575), .Z(G1347GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n589), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n579), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(n580), .Z(n592) );
  INV_X1 U645 ( .A(n592), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n590), .A2(n581), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  OR2_X1 U652 ( .A1(n592), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U656 ( .A1(n488), .A2(n592), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

