//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G219), .A2(G218), .A3(G221), .A4(G220), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n454), .A2(new_n448), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT71), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n463), .B2(new_n465), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n471), .A2(KEYINPUT72), .A3(G101), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT72), .B1(new_n471), .B2(G101), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(KEYINPUT70), .A2(G113), .A3(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n469), .A2(new_n481), .A3(G125), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n469), .A2(new_n481), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT69), .A3(G125), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n467), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n474), .A2(new_n486), .ZN(G160));
  INV_X1    g062(.A(KEYINPUT73), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n466), .A2(new_n469), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n469), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT71), .B(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(KEYINPUT3), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT73), .A3(new_n467), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G136), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n489), .A2(new_n467), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n467), .A2(G112), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n497), .A2(G124), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G162));
  NAND2_X1  g078(.A1(new_n469), .A2(new_n481), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n467), .A3(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G2105), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n466), .A2(new_n469), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n510), .B2(KEYINPUT4), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n512));
  OR2_X1    g087(.A1(G102), .A2(G2105), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n513), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n511), .A2(new_n515), .ZN(G164));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT74), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(new_n521), .B1(KEYINPUT6), .B2(new_n517), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G62), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n524), .A2(G50), .B1(new_n531), .B2(G651), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n518), .A2(new_n521), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n533), .B1(new_n536), .B2(new_n529), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n522), .A2(KEYINPUT75), .A3(new_n528), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G88), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n532), .B1(new_n539), .B2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND3_X1  g117(.A1(new_n537), .A2(G89), .A3(new_n538), .ZN(new_n543));
  XOR2_X1   g118(.A(KEYINPUT76), .B(G51), .Z(new_n544));
  NAND3_X1  g119(.A1(new_n522), .A2(G543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n548));
  AND2_X1   g123(.A1(G63), .A2(G651), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n547), .A2(new_n548), .B1(new_n528), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(G168));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n529), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n524), .A2(G52), .B1(new_n556), .B2(G651), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n537), .A2(G90), .A3(new_n538), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  INV_X1    g135(.A(new_n539), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G81), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n529), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n524), .A2(G43), .B1(new_n565), .B2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n562), .A2(G860), .A3(new_n566), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND3_X1  g146(.A1(new_n522), .A2(G53), .A3(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n537), .A2(G91), .A3(new_n538), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n517), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(G299));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n552), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n543), .A2(KEYINPUT77), .A3(new_n551), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G286));
  OAI21_X1  g157(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n583));
  INV_X1    g158(.A(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n523), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n561), .B2(G87), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G288));
  NAND3_X1  g162(.A1(new_n537), .A2(G86), .A3(new_n538), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n537), .A2(KEYINPUT79), .A3(G86), .A4(new_n538), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n522), .A2(G48), .A3(G543), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n526), .B2(new_n527), .ZN(new_n595));
  AND2_X1   g170(.A1(G73), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT78), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n599), .B(G651), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n593), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n590), .A2(new_n591), .A3(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n517), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n537), .A2(G85), .A3(new_n538), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n524), .A2(G47), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n605), .A2(KEYINPUT80), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT80), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G301), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n529), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n524), .A2(G54), .B1(new_n614), .B2(G651), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n539), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .A4(new_n538), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT81), .Z(new_n622));
  AOI21_X1  g197(.A(new_n611), .B1(new_n622), .B2(new_n610), .ZN(G321));
  XNOR2_X1  g198(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NOR2_X1   g199(.A1(G299), .A2(G868), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n581), .B2(G868), .ZN(G297));
  AOI21_X1  g201(.A(new_n625), .B1(new_n581), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n562), .A2(new_n566), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n628), .ZN(new_n631));
  MUX2_X1   g206(.A(new_n630), .B(new_n631), .S(G868), .Z(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n471), .A2(new_n484), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT83), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n495), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n497), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n467), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  OAI211_X1 g219(.A(new_n638), .B(new_n644), .C1(G2100), .C2(new_n636), .ZN(G156));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2438), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n660), .B(G14), .C1(new_n658), .C2(new_n657), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT86), .ZN(G401));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT17), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2084), .B(G2090), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n665), .B2(new_n663), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT87), .ZN(new_n671));
  INV_X1    g246(.A(new_n668), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n665), .A3(new_n663), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n665), .A2(new_n668), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n664), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT88), .B(G2096), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n683), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G229));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n495), .A2(G131), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n467), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n497), .A2(G119), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT89), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n700), .B1(new_n708), .B2(new_n699), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(KEYINPUT90), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G22), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G166), .B2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G1971), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(G6), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G305), .B2(new_n713), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n713), .A2(G23), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n586), .B2(new_n713), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT33), .B(G1976), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n717), .A2(new_n721), .A3(new_n722), .A4(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n729));
  MUX2_X1   g304(.A(G24), .B(G290), .S(G16), .Z(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1986), .Z(new_n731));
  NAND4_X1  g306(.A1(new_n712), .A2(new_n728), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G19), .B(new_n630), .S(G16), .Z(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  XOR2_X1   g311(.A(KEYINPUT94), .B(KEYINPUT23), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n713), .A2(G20), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G299), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n713), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT95), .B(G1956), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n699), .A2(G26), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT28), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n495), .A2(G140), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n467), .A2(G116), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n497), .A2(G128), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2067), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n699), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n699), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT29), .B(G2090), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n736), .A2(new_n743), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n713), .A2(G4), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n622), .B2(new_n713), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n758), .B1(G1348), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G1348), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n699), .A2(G33), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(new_n467), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT91), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n765), .A2(KEYINPUT91), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n495), .A2(G139), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n763), .B1(new_n772), .B2(new_n699), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2072), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n699), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n699), .ZN(new_n776));
  INV_X1    g351(.A(G2078), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G34), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(KEYINPUT24), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n779), .B2(KEYINPUT24), .ZN(new_n781));
  AOI22_X1  g356(.A1(G160), .A2(G29), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n778), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n713), .A2(G21), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G168), .B2(new_n713), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G1966), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT30), .B(G28), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n699), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n792), .B1(new_n782), .B2(G2084), .C1(new_n643), .C2(new_n699), .ZN(new_n793));
  NOR4_X1   g368(.A1(new_n774), .A2(new_n785), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n699), .A2(G32), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n495), .A2(G141), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT92), .Z(new_n797));
  NAND3_X1  g372(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT26), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n471), .A2(G105), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n799), .B(new_n800), .C1(new_n497), .C2(G129), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n795), .B1(new_n803), .B2(new_n699), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT27), .B(G1996), .Z(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n713), .A2(G5), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G171), .B2(new_n713), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1961), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G1966), .B2(new_n787), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n794), .A2(new_n806), .A3(new_n807), .A4(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n762), .B1(new_n812), .B2(KEYINPUT93), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n732), .A2(new_n733), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n812), .A2(KEYINPUT93), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n734), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND2_X1  g392(.A1(G80), .A2(G543), .ZN(new_n818));
  INV_X1    g393(.A(G67), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n529), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n524), .A2(G55), .B1(new_n820), .B2(G651), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n537), .A2(G93), .A3(new_n538), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n821), .B2(new_n822), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n630), .B1(new_n824), .B2(new_n825), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n562), .A2(new_n566), .A3(new_n822), .A4(new_n821), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n622), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT97), .ZN(new_n837));
  AOI21_X1  g412(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n828), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT98), .ZN(G145));
  XNOR2_X1  g415(.A(G162), .B(new_n643), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G160), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n515), .A2(KEYINPUT100), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n512), .A2(new_n845), .A3(new_n514), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n505), .B1(new_n493), .B2(new_n509), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(new_n507), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n511), .A2(KEYINPUT99), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n751), .B(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n853), .A2(new_n772), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n772), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n854), .A2(new_n855), .A3(new_n802), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n495), .A2(G142), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n467), .A2(G118), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n497), .A2(G130), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n706), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n635), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n701), .A2(KEYINPUT101), .A3(new_n705), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  INV_X1    g446(.A(new_n862), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n802), .B1(new_n854), .B2(new_n855), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n856), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n874), .B1(new_n856), .B2(new_n875), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n856), .A2(KEYINPUT102), .A3(new_n874), .A4(new_n875), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n843), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n877), .A2(new_n842), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n883), .B2(new_n876), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g461(.A1(new_n826), .A2(new_n610), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n605), .A2(new_n606), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT80), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n605), .A2(KEYINPUT80), .A3(new_n606), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n586), .B1(new_n893), .B2(new_n604), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n586), .B(new_n604), .C1(new_n607), .C2(new_n608), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n888), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(G290), .A2(G288), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(KEYINPUT104), .A3(new_n895), .ZN(new_n899));
  XNOR2_X1  g474(.A(G305), .B(G303), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n900), .A2(KEYINPUT104), .A3(new_n898), .A4(new_n895), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(KEYINPUT105), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n829), .A2(new_n830), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n631), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n621), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n740), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT103), .B1(new_n621), .B2(G299), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n621), .A2(G299), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT41), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n917), .A2(new_n918), .A3(new_n922), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n914), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n914), .A2(new_n920), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n912), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(new_n909), .A3(new_n911), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n887), .B1(new_n930), .B2(new_n610), .ZN(G295));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n932), .B(new_n887), .C1(new_n930), .C2(new_n610), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n610), .B1(new_n927), .B2(new_n929), .ZN(new_n934));
  INV_X1    g509(.A(new_n887), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT106), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n933), .A2(new_n936), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(G168), .B2(G301), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n581), .B2(G301), .ZN(new_n941));
  NAND4_X1  g516(.A1(G171), .A2(new_n579), .A3(new_n939), .A4(new_n580), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n913), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n831), .A2(new_n941), .A3(new_n942), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n921), .A2(new_n944), .A3(new_n923), .A4(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n945), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n831), .B1(new_n941), .B2(new_n942), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n920), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n906), .A3(new_n907), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n951), .A2(KEYINPUT108), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT108), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n902), .A2(KEYINPUT105), .A3(new_n903), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT105), .B1(new_n902), .B2(new_n903), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(new_n950), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n908), .A2(KEYINPUT109), .A3(new_n949), .A4(new_n946), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n938), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT43), .B1(new_n960), .B2(new_n961), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n951), .A2(new_n952), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n963), .A2(new_n967), .A3(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(new_n966), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT110), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n962), .A2(new_n971), .A3(new_n966), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(KEYINPUT43), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n955), .A2(new_n964), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n968), .B1(new_n975), .B2(KEYINPUT44), .ZN(G397));
  AOI211_X1 g551(.A(new_n848), .B(new_n507), .C1(KEYINPUT4), .C2(new_n510), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n978));
  INV_X1    g553(.A(new_n507), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT99), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n981), .B2(new_n847), .ZN(new_n982));
  INV_X1    g557(.A(new_n486), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n472), .A2(new_n473), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n984), .A3(G40), .A4(new_n470), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n982), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  OR3_X1    g562(.A1(new_n987), .A2(G1986), .A3(G290), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(G1986), .A3(G290), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n990), .B(KEYINPUT111), .Z(new_n991));
  NOR2_X1   g566(.A1(new_n802), .A2(G1996), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G2067), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n751), .B(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(G1996), .B2(new_n802), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n987), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n706), .B(new_n710), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n999), .B1(new_n987), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n991), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n590), .A2(new_n1003), .A3(new_n601), .A4(new_n591), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n588), .A2(new_n597), .A3(new_n592), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G1981), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT113), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT112), .B(G8), .Z(new_n1012));
  INV_X1    g587(.A(G40), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n474), .A2(new_n486), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n982), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1010), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G288), .A2(G1976), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1005), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n852), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n511), .B2(new_n515), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT50), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1029), .A2(new_n1014), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(G2090), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n985), .B1(new_n1033), .B2(new_n1028), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n1026), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1971), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(G8), .B(new_n1024), .C1(new_n1032), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n982), .A2(new_n1014), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1012), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n586), .A2(G1976), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1015), .A2(new_n1044), .A3(new_n1040), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1011), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1015), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1042), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1020), .A2(new_n1021), .B1(new_n1037), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1025), .B1(new_n852), .B2(new_n1026), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n985), .ZN(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  OAI211_X1 g628(.A(KEYINPUT115), .B(new_n1014), .C1(new_n982), .C2(new_n1025), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1028), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1025), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1036), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1024), .B1(new_n1059), .B2(new_n1039), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1037), .A2(new_n1016), .A3(new_n1045), .A4(new_n1042), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1055), .A2(KEYINPUT45), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1014), .B(new_n1063), .C1(new_n982), .C2(KEYINPUT45), .ZN(new_n1064));
  INV_X1    g639(.A(G1966), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1029), .A2(new_n1014), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n982), .B2(new_n1025), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n784), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1012), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(G286), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1062), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1062), .A2(new_n1076), .A3(new_n1072), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1037), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(new_n1048), .ZN(new_n1080));
  OAI21_X1  g655(.A(G8), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1024), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1075), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1072), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1049), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n1070), .B2(new_n552), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n552), .A2(new_n1039), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1064), .A2(new_n1065), .B1(new_n1068), .B2(new_n784), .ZN(new_n1089));
  INV_X1    g664(.A(G8), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1086), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1087), .A2(new_n1091), .B1(new_n1071), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1094), .A2(KEYINPUT62), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1059), .A2(new_n1039), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1082), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1031), .A2(KEYINPUT118), .ZN(new_n1098));
  INV_X1    g673(.A(G1961), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1027), .A2(new_n1030), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(G2078), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n850), .A2(new_n851), .ZN(new_n1106));
  INV_X1    g681(.A(new_n846), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n845), .B1(new_n512), .B2(new_n514), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1026), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n985), .B1(new_n1110), .B2(new_n1033), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1111), .A2(KEYINPUT53), .A3(new_n777), .A4(new_n1063), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1102), .A2(new_n1105), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1097), .A2(new_n1114), .A3(new_n1080), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1966), .B1(new_n1111), .B2(new_n1063), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1031), .A2(G2084), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n552), .B(new_n1039), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1091), .A2(KEYINPUT51), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1071), .A2(new_n1093), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT62), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1095), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT123), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT124), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1113), .A2(G171), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1060), .A2(new_n1061), .A3(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(new_n1123), .C1(KEYINPUT62), .C2(new_n1094), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1094), .A2(KEYINPUT62), .ZN(new_n1130));
  AND4_X1   g705(.A1(KEYINPUT124), .A2(new_n1129), .A3(new_n1125), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1085), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1111), .A2(KEYINPUT53), .A3(new_n777), .A4(new_n1035), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1102), .A2(new_n1105), .A3(new_n1133), .ZN(new_n1134));
  OR3_X1    g709(.A1(new_n1134), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT122), .B1(new_n1134), .B2(G171), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1135), .B(new_n1136), .C1(new_n1114), .C2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1134), .B2(G171), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(G171), .B2(new_n1113), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1138), .A2(new_n1094), .A3(new_n1062), .A4(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(G299), .B(KEYINPUT57), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1056), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n985), .B1(new_n1110), .B2(KEYINPUT50), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(KEYINPUT115), .ZN(new_n1145));
  AOI21_X1  g720(.A(G1956), .B1(new_n1145), .B2(new_n1052), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1104), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT56), .B(G2072), .Z(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT117), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1142), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1052), .A2(new_n1056), .A3(new_n1054), .ZN(new_n1153));
  INV_X1    g728(.A(G1956), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1142), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n1150), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1152), .A2(KEYINPUT61), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT120), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1152), .A2(new_n1163), .A3(new_n1157), .A4(KEYINPUT61), .ZN(new_n1164));
  XOR2_X1   g739(.A(KEYINPUT58), .B(G1341), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1038), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(G1996), .B2(new_n1104), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n630), .A2(KEYINPUT119), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1159), .A2(new_n1162), .A3(new_n1164), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT121), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1161), .B2(new_n1160), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n1164), .A4(new_n1159), .ZN(new_n1177));
  INV_X1    g752(.A(G1348), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1098), .A2(new_n1178), .A3(new_n1101), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n982), .A2(new_n994), .A3(new_n1014), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT60), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(new_n621), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(KEYINPUT60), .B2(new_n1181), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1174), .A2(new_n1177), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1152), .B1(new_n915), .B2(new_n1181), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1157), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1141), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1002), .B1(new_n1132), .B2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n988), .B(KEYINPUT48), .Z(new_n1190));
  NOR2_X1   g765(.A1(new_n1001), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT46), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n803), .B1(new_n1192), .B2(G1996), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n986), .B1(new_n1193), .B2(new_n996), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1192), .B1(new_n987), .B2(G1996), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT47), .Z(new_n1199));
  NAND2_X1  g774(.A1(new_n708), .A2(new_n710), .ZN(new_n1200));
  OAI22_X1  g775(.A1(new_n998), .A2(new_n1200), .B1(G2067), .B2(new_n751), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n987), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n1191), .B(new_n1199), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1189), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1208));
  INV_X1    g782(.A(KEYINPUT108), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n951), .A2(KEYINPUT108), .A3(new_n952), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n962), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI22_X1  g786(.A1(new_n1212), .A2(KEYINPUT43), .B1(new_n966), .B2(new_n964), .ZN(new_n1213));
  NOR3_X1   g787(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1214));
  INV_X1    g788(.A(new_n884), .ZN(new_n1215));
  OAI211_X1 g789(.A(new_n661), .B(new_n1214), .C1(new_n1215), .C2(new_n881), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1208), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n661), .A2(new_n1214), .ZN(new_n1218));
  AOI21_X1  g792(.A(new_n1218), .B1(new_n882), .B2(new_n884), .ZN(new_n1219));
  OAI211_X1 g793(.A(new_n1219), .B(KEYINPUT127), .C1(new_n963), .C2(new_n967), .ZN(new_n1220));
  AND2_X1   g794(.A1(new_n1217), .A2(new_n1220), .ZN(G308));
  NAND2_X1  g795(.A1(new_n1217), .A2(new_n1220), .ZN(G225));
endmodule


