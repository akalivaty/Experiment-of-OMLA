//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT3), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n187), .A2(KEYINPUT3), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n188), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n192), .B2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n196), .A2(G104), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n188), .B2(new_n190), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n195), .B1(new_n203), .B2(new_n197), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(KEYINPUT4), .A3(new_n205), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT2), .B(G113), .Z(new_n207));
  XNOR2_X1  g021(.A(G116), .B(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G116), .ZN(new_n211));
  INV_X1    g025(.A(G116), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT2), .B(G113), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(KEYINPUT67), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n207), .A2(new_n208), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n214), .A2(new_n215), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(G101), .C1(new_n192), .C2(new_n198), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n206), .A2(new_n217), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT5), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n210), .A3(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT81), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n228), .A2(new_n225), .A3(new_n210), .A4(G116), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G113), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n208), .B2(KEYINPUT5), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n220), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n190), .B2(new_n200), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n205), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n224), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n224), .A2(KEYINPUT82), .A3(new_n235), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n238), .A2(new_n239), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n224), .A2(KEYINPUT82), .A3(new_n235), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT82), .B1(new_n224), .B2(new_n235), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n244), .A2(new_n245), .A3(new_n241), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n221), .A2(new_n217), .A3(new_n223), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n199), .A2(KEYINPUT4), .A3(new_n205), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n235), .B(new_n241), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT6), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT83), .B(new_n243), .C1(new_n246), .C2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n238), .A2(new_n239), .A3(new_n242), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT6), .A4(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT0), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT0), .B(G128), .Z(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G125), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n256), .A2(new_n263), .A3(G128), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  INV_X1    g079(.A(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G143), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G146), .ZN(new_n269));
  AOI21_X1  g083(.A(G128), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n263), .A2(new_n266), .A3(G143), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n266), .A2(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT1), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(KEYINPUT66), .C1(new_n256), .C2(G128), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n264), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n262), .B1(new_n276), .B2(G125), .ZN(new_n277));
  INV_X1    g091(.A(G224), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n279), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n262), .B(new_n281), .C1(new_n276), .C2(G125), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n255), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n280), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n256), .A2(new_n263), .A3(G128), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n268), .A2(G146), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n258), .B1(new_n292), .B2(new_n273), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT66), .B1(new_n293), .B2(new_n274), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n270), .A2(new_n265), .A3(new_n271), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G125), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n298), .A2(new_n288), .A3(new_n281), .A4(new_n262), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n205), .A2(new_n234), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n208), .A2(KEYINPUT5), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(G113), .A3(new_n227), .A4(new_n229), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n209), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n205), .A2(new_n234), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n233), .B1(new_n306), .B2(KEYINPUT84), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n241), .B(KEYINPUT8), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n290), .A2(new_n249), .A3(new_n299), .A4(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n287), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n280), .A2(new_n282), .A3(new_n289), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n299), .A2(new_n249), .A3(new_n309), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n287), .B(new_n311), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n285), .A2(new_n286), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n286), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n283), .B1(new_n251), .B2(new_n254), .ZN(new_n320));
  INV_X1    g134(.A(new_n316), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(new_n312), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(G221), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT9), .B(G234), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n326), .B1(new_n328), .B2(new_n311), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n205), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n296), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n206), .A2(new_n261), .A3(new_n223), .ZN(new_n332));
  INV_X1    g146(.A(G131), .ZN(new_n333));
  INV_X1    g147(.A(G137), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(G134), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT64), .ZN(new_n337));
  INV_X1    g151(.A(G134), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n337), .B(KEYINPUT11), .C1(new_n338), .C2(G137), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n334), .A2(G134), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT11), .B1(new_n341), .B2(new_n337), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n336), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT65), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n337), .B1(new_n338), .B2(G137), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT11), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n339), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT65), .A3(new_n336), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n338), .A2(G137), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n340), .B2(new_n342), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n345), .A2(new_n350), .B1(G131), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n291), .A2(new_n293), .A3(new_n274), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n205), .A3(new_n234), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n331), .A2(new_n332), .A3(new_n353), .A4(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G140), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT75), .ZN(new_n360));
  INV_X1    g174(.A(G227), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G953), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n360), .B(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n331), .A2(new_n332), .A3(new_n357), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n353), .B1(new_n365), .B2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n331), .A2(new_n332), .A3(new_n357), .A4(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n364), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n355), .B1(new_n296), .B2(new_n300), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n352), .A2(G131), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT65), .B1(new_n349), .B2(new_n336), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n344), .B(new_n335), .C1(new_n348), .C2(new_n339), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(KEYINPUT77), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT12), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(KEYINPUT78), .A3(new_n374), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT12), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n276), .A2(new_n306), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n345), .A2(new_n350), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n381), .A2(new_n355), .B1(new_n382), .B2(new_n371), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT78), .B1(new_n383), .B2(KEYINPUT77), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n377), .B(new_n358), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n363), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n369), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G469), .B1(new_n387), .B2(G902), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n377), .B1(new_n380), .B2(new_n384), .ZN(new_n389));
  INV_X1    g203(.A(new_n358), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n366), .B2(new_n368), .ZN(new_n391));
  OAI22_X1  g205(.A1(new_n389), .A2(new_n364), .B1(new_n391), .B2(new_n363), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT80), .B(G469), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n311), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n329), .B1(new_n388), .B2(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n324), .A2(new_n325), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n221), .A2(new_n217), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n374), .A2(new_n261), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n341), .A2(new_n351), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G131), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n382), .A2(new_n296), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n400), .B2(new_n403), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n403), .A3(new_n398), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(G237), .A2(G953), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G210), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT27), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G101), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n400), .A2(new_n403), .A3(new_n398), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n398), .B1(new_n400), .B2(new_n403), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT28), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT68), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n417), .C2(new_n418), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT28), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n415), .B1(new_n408), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n400), .A2(new_n403), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n399), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT69), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n408), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(KEYINPUT69), .A3(new_n399), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(KEYINPUT28), .A3(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n424), .A2(KEYINPUT29), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G472), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n408), .A2(new_n423), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n421), .A2(new_n422), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n415), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n407), .A2(new_n408), .A3(new_n414), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT31), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n407), .A2(KEYINPUT31), .A3(new_n408), .A4(new_n414), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(G472), .A2(G902), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT32), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  AOI211_X1 g263(.A(G472), .B(G902), .C1(new_n439), .C2(new_n444), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n436), .B(new_n449), .C1(new_n450), .C2(KEYINPUT32), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT71), .B1(new_n210), .B2(G128), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n258), .A3(G119), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n452), .B(new_n454), .C1(G119), .C2(new_n258), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT24), .B(G110), .ZN(new_n456));
  OR3_X1    g270(.A1(new_n455), .A2(KEYINPUT72), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT72), .B1(new_n455), .B2(new_n456), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G125), .B(G140), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT16), .ZN(new_n461));
  INV_X1    g275(.A(G140), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G125), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n463), .A2(KEYINPUT16), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n266), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(G146), .A3(new_n464), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT23), .B1(new_n258), .B2(G119), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT73), .B1(new_n210), .B2(G128), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n469), .B(new_n470), .Z(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G110), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n459), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n455), .A2(new_n456), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n471), .B2(G110), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n460), .A2(new_n266), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n467), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT22), .B(G137), .ZN(new_n479));
  INV_X1    g293(.A(G234), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n326), .A2(new_n480), .A3(G953), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n479), .B(new_n481), .Z(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n473), .A2(new_n477), .A3(new_n482), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n311), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT25), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n484), .A2(KEYINPUT25), .A3(new_n311), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G217), .B1(new_n480), .B2(G902), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT70), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n484), .A2(KEYINPUT74), .A3(new_n485), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT74), .B1(new_n484), .B2(new_n485), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(G128), .B(G143), .Z(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT91), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n501), .A2(new_n338), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT88), .B(G122), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n503), .A2(new_n212), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT14), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n212), .A2(G122), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n503), .A2(new_n212), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n505), .B(G107), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n504), .B(new_n506), .C1(KEYINPUT14), .C2(new_n196), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(new_n338), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n502), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G953), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n328), .A2(G217), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n504), .A2(new_n196), .A3(new_n506), .ZN(new_n516));
  OAI21_X1  g330(.A(G107), .B1(new_n508), .B2(new_n507), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n519), .A2(KEYINPUT13), .B1(new_n268), .B2(G128), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n519), .A2(KEYINPUT13), .ZN(new_n521));
  OAI21_X1  g335(.A(G134), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(new_n500), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n518), .B2(new_n523), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n512), .B(new_n515), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n518), .A2(new_n523), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT90), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n525), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n515), .B1(new_n532), .B2(new_n512), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n311), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n410), .A2(G143), .A3(G214), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G143), .B1(new_n410), .B2(G214), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT18), .B(G131), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n297), .A2(G140), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n463), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G146), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n476), .ZN(new_n545));
  INV_X1    g359(.A(new_n540), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT18), .A2(G131), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n538), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n541), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n541), .A2(new_n548), .A3(new_n545), .A4(KEYINPUT86), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n546), .A2(new_n333), .A3(new_n538), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n557), .A3(new_n555), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n556), .A2(new_n558), .A3(new_n466), .A4(new_n467), .ZN(new_n559));
  XNOR2_X1  g373(.A(G113), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(new_n189), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n553), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n563));
  INV_X1    g377(.A(new_n467), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT19), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n543), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n460), .A2(KEYINPUT19), .ZN(new_n567));
  AOI21_X1  g381(.A(G146), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n563), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n467), .B(KEYINPUT87), .C1(new_n570), .C2(G146), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n554), .A2(new_n557), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n561), .B1(new_n573), .B2(new_n553), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n562), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G475), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT20), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT20), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n579), .B(new_n576), .C1(new_n562), .C2(new_n574), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI221_X1 g395(.A(new_n311), .B1(KEYINPUT15), .B2(new_n535), .C1(new_n529), .C2(new_n533), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n561), .B1(new_n553), .B2(new_n559), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n311), .B1(new_n562), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G475), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n537), .A2(new_n581), .A3(new_n582), .A4(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G952), .ZN(new_n587));
  AOI211_X1 g401(.A(G953), .B(new_n587), .C1(G234), .C2(G237), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n311), .B(new_n513), .C1(G234), .C2(G237), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT21), .B(G898), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n499), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n397), .A2(new_n451), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  AOI22_X1  g408(.A1(new_n438), .A2(new_n415), .B1(new_n442), .B2(new_n443), .ZN(new_n595));
  OAI21_X1  g409(.A(G472), .B1(new_n595), .B2(G902), .ZN(new_n596));
  INV_X1    g410(.A(G472), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n445), .A2(new_n597), .A3(new_n311), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n325), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n600), .B(new_n591), .C1(new_n318), .C2(new_n323), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n388), .A2(new_n395), .ZN(new_n602));
  INV_X1    g416(.A(new_n329), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n499), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n535), .A2(G902), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n532), .A2(new_n512), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n514), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n528), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT92), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n528), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n609), .B(new_n528), .C1(new_n612), .C2(new_n611), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n607), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT93), .B(G478), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n610), .B2(new_n311), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n581), .A2(new_n585), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n599), .A2(new_n601), .A3(new_n605), .A4(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  AND2_X1   g439(.A1(new_n537), .A2(new_n582), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n620), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n599), .A2(new_n601), .A3(new_n605), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  OR2_X1    g444(.A1(new_n483), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n478), .B(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n490), .A2(new_n492), .B1(new_n494), .B2(new_n633), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n586), .A2(new_n634), .A3(new_n591), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n596), .A2(new_n635), .A3(new_n598), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n397), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n600), .B1(new_n318), .B2(new_n323), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n436), .A2(new_n449), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n439), .B2(new_n444), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT32), .B1(new_n643), .B2(new_n597), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n641), .B(new_n396), .C1(new_n642), .C2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n589), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n588), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n627), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n634), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n640), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n650), .A2(new_n634), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n397), .A2(new_n451), .A3(new_n655), .A4(KEYINPUT94), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XNOR2_X1  g472(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n324), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n649), .B(KEYINPUT39), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n396), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT40), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n447), .B1(new_n439), .B2(new_n444), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n409), .A2(new_n414), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n430), .A2(new_n431), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n665), .B(new_n311), .C1(new_n414), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT96), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n670), .A3(G472), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n664), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT32), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n598), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n621), .A2(new_n626), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n325), .A3(new_n634), .ZN(new_n677));
  OR4_X1    g491(.A1(new_n660), .A2(new_n663), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  OAI211_X1 g493(.A(new_n620), .B(new_n649), .C1(new_n616), .C2(new_n618), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n645), .A2(new_n634), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n266), .ZN(G48));
  AOI21_X1  g496(.A(new_n664), .B1(G472), .B2(new_n435), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n499), .B1(new_n683), .B2(new_n674), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n392), .A2(new_n311), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n603), .A3(new_n395), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n684), .A2(new_n622), .A3(new_n601), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT97), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n689), .B(new_n691), .ZN(G15));
  INV_X1    g506(.A(new_n591), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n641), .A2(new_n693), .A3(new_n627), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n684), .A2(new_n694), .A3(new_n688), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AND2_X1   g510(.A1(new_n688), .A2(new_n641), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n451), .A3(new_n635), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  AND2_X1   g513(.A1(new_n432), .A2(new_n437), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n444), .B1(new_n414), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n446), .ZN(new_n702));
  INV_X1    g516(.A(new_n499), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n596), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n686), .A2(new_n603), .A3(new_n395), .A4(new_n693), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT98), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n641), .A2(new_n707), .A3(new_n676), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n707), .B1(new_n641), .B2(new_n676), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  INV_X1    g525(.A(new_n680), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n688), .A2(new_n641), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n596), .A2(new_n702), .A3(new_n652), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT99), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n596), .A2(new_n702), .A3(KEYINPUT99), .A4(new_n652), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n297), .ZN(G27));
  NAND3_X1  g533(.A1(new_n318), .A2(new_n323), .A3(new_n325), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n604), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n712), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT100), .B1(new_n595), .B2(new_n447), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT100), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n445), .A2(new_n726), .A3(new_n448), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT101), .B1(new_n728), .B2(new_n644), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n674), .A2(new_n730), .A3(new_n725), .A4(new_n727), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n731), .A3(new_n436), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n724), .A2(new_n732), .A3(new_n703), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n684), .A2(new_n721), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n723), .B1(new_n734), .B2(new_n680), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT102), .B(G131), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G33));
  NAND4_X1  g552(.A1(new_n451), .A2(new_n721), .A3(new_n651), .A4(new_n703), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n619), .B2(new_n620), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n621), .B(new_n742), .C1(new_n616), .C2(new_n618), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n599), .B2(new_n634), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n596), .A2(new_n598), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(KEYINPUT104), .A3(new_n652), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n744), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  OR3_X1    g563(.A1(new_n749), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n750));
  NAND2_X1  g564(.A1(G469), .A2(G902), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n387), .A2(KEYINPUT45), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n387), .B2(KEYINPUT45), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n395), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n329), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n661), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT103), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT105), .B1(new_n749), .B2(KEYINPUT44), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n720), .B1(new_n749), .B2(KEYINPUT44), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n750), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  NOR4_X1   g579(.A1(new_n451), .A2(new_n703), .A3(new_n680), .A4(new_n720), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT106), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n660), .A2(new_n600), .A3(new_n688), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n741), .A2(new_n588), .A3(new_n743), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n741), .A2(new_n776), .A3(new_n588), .A4(new_n743), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n704), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n773), .B(new_n778), .C1(KEYINPUT112), .C2(KEYINPUT50), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n687), .B(new_n720), .C1(new_n775), .C2(new_n777), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n716), .A2(new_n717), .ZN(new_n785));
  INV_X1    g599(.A(new_n720), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n499), .A2(new_n648), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n675), .A2(new_n688), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n619), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n620), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n784), .A2(new_n785), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n783), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n686), .A2(new_n395), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n603), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n769), .A2(new_n768), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n778), .A2(new_n786), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n772), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n732), .A2(new_n703), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n784), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n788), .A2(new_n622), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n587), .B(G953), .C1(new_n778), .C2(new_n697), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n800), .A2(new_n801), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n798), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n783), .A2(new_n791), .A3(KEYINPUT51), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n795), .A2(KEYINPUT113), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n796), .B1(new_n795), .B2(KEYINPUT113), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n689), .A2(new_n710), .A3(new_n695), .A4(new_n698), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n733), .B2(new_n735), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n593), .A2(new_n623), .A3(new_n628), .A4(new_n637), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n722), .B1(new_n716), .B2(new_n717), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n634), .B(new_n586), .C1(new_n648), .C2(new_n647), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n451), .A2(new_n721), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n739), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n324), .A2(new_n325), .A3(new_n676), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n641), .A2(new_n707), .A3(new_n676), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n396), .A2(new_n634), .A3(new_n649), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n672), .B2(new_n674), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n286), .B1(new_n285), .B2(new_n317), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n320), .A2(new_n322), .A3(new_n319), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n396), .B(new_n325), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n674), .B2(new_n683), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n680), .A2(new_n634), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n825), .A2(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n718), .ZN(new_n834));
  AND4_X1   g648(.A1(KEYINPUT52), .A2(new_n657), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n718), .B1(new_n654), .B2(new_n656), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(new_n836), .B2(new_n833), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n815), .B(new_n821), .C1(new_n835), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n657), .A2(new_n833), .A3(new_n834), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(KEYINPUT52), .A3(new_n833), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n689), .A2(new_n710), .A3(new_n695), .A4(new_n698), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n821), .A2(new_n736), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT54), .B1(new_n840), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n835), .A2(new_n837), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n821), .A2(KEYINPUT53), .A3(new_n736), .A4(new_n846), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT110), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n815), .A2(new_n821), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n839), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT110), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n845), .A2(new_n855), .A3(new_n856), .A4(new_n815), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n852), .A2(new_n854), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n813), .A2(new_n849), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n587), .A2(new_n513), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n789), .A2(new_n621), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n703), .A2(new_n325), .A3(new_n603), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n863), .B(new_n864), .C1(KEYINPUT49), .C2(new_n793), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT107), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n660), .A3(new_n867), .A4(new_n675), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT108), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT115), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n862), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n513), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n852), .A2(new_n854), .A3(new_n857), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(G210), .A3(G902), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n255), .B(new_n284), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT55), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n876), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT56), .B1(new_n878), .B2(KEYINPUT116), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(KEYINPUT116), .B2(new_n878), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(new_n881), .ZN(G51));
  NAND2_X1  g700(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n888), .A3(new_n859), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n877), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n751), .B(KEYINPUT117), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n392), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n752), .A2(new_n753), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n877), .A2(G902), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n875), .B1(new_n894), .B2(new_n896), .ZN(G54));
  NAND4_X1  g711(.A1(new_n877), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n898), .A2(new_n575), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n575), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n875), .ZN(G60));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT59), .Z(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n849), .B2(new_n859), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n614), .A2(new_n615), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n876), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n889), .A2(new_n890), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n614), .B2(new_n615), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT60), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n877), .A2(new_n633), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n851), .B1(new_n843), .B2(new_n844), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n914), .A2(new_n855), .B1(new_n838), .B2(new_n839), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n915), .B2(new_n852), .ZN(new_n916));
  INV_X1    g730(.A(new_n498), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n876), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(KEYINPUT119), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(KEYINPUT119), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n877), .A2(new_n912), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n875), .B1(new_n923), .B2(new_n498), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n924), .A2(KEYINPUT119), .A3(new_n919), .A4(new_n913), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(G66));
  OAI21_X1  g740(.A(G953), .B1(new_n590), .B2(new_n278), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n814), .A2(new_n816), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n251), .B(new_n254), .C1(G898), .C2(new_n513), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT120), .Z(new_n931));
  XNOR2_X1  g745(.A(new_n929), .B(new_n931), .ZN(G69));
  OR2_X1    g746(.A1(new_n405), .A2(new_n406), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n570), .B(KEYINPUT121), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n764), .A2(new_n770), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n761), .A2(new_n825), .A3(new_n799), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n736), .A2(new_n739), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n718), .B(new_n681), .C1(new_n654), .C2(new_n656), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n942), .A3(KEYINPUT125), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n936), .B2(new_n941), .ZN(new_n945));
  AOI21_X1  g759(.A(G953), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n513), .A2(G900), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n935), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n940), .A2(new_n678), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n661), .B1(new_n622), .B2(new_n627), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n734), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT123), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n937), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n513), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n935), .B(KEYINPUT122), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n361), .B2(new_n646), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n948), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n948), .B2(new_n958), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(G72));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  INV_X1    g779(.A(new_n928), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n955), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n665), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n876), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n943), .A2(new_n945), .A3(new_n928), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n414), .B(new_n409), .C1(new_n971), .C2(new_n965), .ZN(new_n972));
  INV_X1    g786(.A(new_n440), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n414), .B1(new_n407), .B2(new_n408), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT126), .Z(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n840), .B2(new_n848), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT127), .Z(new_n978));
  NOR3_X1   g792(.A1(new_n970), .A2(new_n972), .A3(new_n978), .ZN(G57));
endmodule


