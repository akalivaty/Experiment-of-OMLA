

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n516, n517, n518, n519, n520, n521, n522, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778;

  NOR2_X1 U367 ( .A1(n613), .A2(KEYINPUT89), .ZN(n373) );
  AND2_X1 U368 ( .A1(n561), .A2(n602), .ZN(n612) );
  NOR2_X1 U369 ( .A1(n557), .A2(n534), .ZN(n559) );
  AND2_X1 U370 ( .A1(n401), .A2(n733), .ZN(n347) );
  XNOR2_X1 U371 ( .A(n541), .B(n540), .ZN(n745) );
  XNOR2_X1 U372 ( .A(n526), .B(KEYINPUT114), .ZN(n734) );
  XNOR2_X1 U373 ( .A(n522), .B(G478), .ZN(n590) );
  XNOR2_X1 U374 ( .A(n348), .B(n513), .ZN(n520) );
  XNOR2_X1 U375 ( .A(n514), .B(n349), .ZN(n348) );
  INV_X1 U376 ( .A(KEYINPUT110), .ZN(n349) );
  XNOR2_X1 U377 ( .A(G116), .B(KEYINPUT9), .ZN(n511) );
  XNOR2_X1 U378 ( .A(G104), .B(G122), .ZN(n500) );
  NAND2_X1 U379 ( .A1(G234), .A2(G237), .ZN(n438) );
  INV_X1 U380 ( .A(G104), .ZN(n430) );
  XNOR2_X2 U381 ( .A(n476), .B(n475), .ZN(n553) );
  NAND2_X4 U382 ( .A1(n651), .A2(G953), .ZN(n686) );
  XNOR2_X2 U383 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n546) );
  XNOR2_X2 U384 ( .A(n565), .B(KEYINPUT30), .ZN(n566) );
  XNOR2_X2 U385 ( .A(n346), .B(KEYINPUT111), .ZN(n591) );
  NOR2_X2 U386 ( .A1(n589), .A2(n590), .ZN(n346) );
  NAND2_X1 U387 ( .A1(n584), .A2(n347), .ZN(n557) );
  XOR2_X2 U388 ( .A(n434), .B(KEYINPUT86), .Z(n383) );
  XOR2_X2 U389 ( .A(KEYINPUT62), .B(n648), .Z(n649) );
  XNOR2_X2 U390 ( .A(n378), .B(n655), .ZN(n657) );
  XNOR2_X2 U391 ( .A(n379), .B(n663), .ZN(n665) );
  XNOR2_X2 U392 ( .A(n380), .B(n671), .ZN(n673) );
  XNOR2_X2 U393 ( .A(n382), .B(n383), .ZN(n560) );
  AND2_X2 U394 ( .A1(n374), .A2(n371), .ZN(n370) );
  OR2_X2 U395 ( .A1(n405), .A2(n603), .ZN(n404) );
  XNOR2_X1 U396 ( .A(G113), .B(G143), .ZN(n506) );
  INV_X1 U397 ( .A(G953), .ZN(n755) );
  BUF_X1 U398 ( .A(G107), .Z(n413) );
  XNOR2_X2 U399 ( .A(KEYINPUT79), .B(n491), .ZN(n505) );
  NAND2_X2 U400 ( .A1(n356), .A2(n355), .ZN(n354) );
  XNOR2_X2 U401 ( .A(n414), .B(n361), .ZN(n525) );
  NOR2_X1 U402 ( .A1(n600), .A2(n599), .ZN(n601) );
  AND2_X1 U403 ( .A1(n598), .A2(KEYINPUT47), .ZN(n599) );
  OR2_X1 U404 ( .A1(n597), .A2(n629), .ZN(n598) );
  OR2_X1 U405 ( .A1(n705), .A2(n693), .ZN(n628) );
  AND2_X1 U406 ( .A1(n576), .A2(n411), .ZN(n594) );
  XNOR2_X1 U407 ( .A(n416), .B(KEYINPUT81), .ZN(n603) );
  OR2_X1 U408 ( .A1(n573), .A2(n719), .ZN(n575) );
  XNOR2_X1 U409 ( .A(n769), .B(n420), .ZN(n419) );
  AND2_X1 U410 ( .A1(n353), .A2(n352), .ZN(n355) );
  NAND2_X1 U411 ( .A1(n610), .A2(n609), .ZN(n395) );
  INV_X1 U412 ( .A(n678), .ZN(n372) );
  NOR2_X1 U413 ( .A1(n680), .A2(n578), .ZN(n580) );
  AND2_X1 U414 ( .A1(n679), .A2(n623), .ZN(n636) );
  XNOR2_X1 U415 ( .A(n410), .B(n366), .ZN(n680) );
  NAND2_X1 U416 ( .A1(n403), .A2(n360), .ZN(n410) );
  XNOR2_X1 U417 ( .A(n529), .B(n528), .ZN(n619) );
  XNOR2_X1 U418 ( .A(n575), .B(n574), .ZN(n576) );
  AND2_X1 U419 ( .A1(n733), .A2(n731), .ZN(n570) );
  XNOR2_X1 U420 ( .A(n602), .B(KEYINPUT38), .ZN(n731) );
  XNOR2_X1 U421 ( .A(G137), .B(G110), .ZN(n453) );
  XNOR2_X2 U422 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n424) );
  XNOR2_X1 U423 ( .A(G116), .B(G113), .ZN(n432) );
  XNOR2_X2 U424 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n425) );
  INV_X2 U425 ( .A(G237), .ZN(n433) );
  XNOR2_X2 U426 ( .A(G146), .B(G125), .ZN(n460) );
  XNOR2_X2 U427 ( .A(KEYINPUT3), .B(G119), .ZN(n431) );
  XNOR2_X1 U428 ( .A(G137), .B(G131), .ZN(n480) );
  XOR2_X1 U429 ( .A(KEYINPUT106), .B(KEYINPUT11), .Z(n501) );
  AND2_X1 U430 ( .A1(n754), .A2(n638), .ZN(n421) );
  XNOR2_X1 U431 ( .A(n357), .B(KEYINPUT72), .ZN(n356) );
  NAND2_X1 U432 ( .A1(n637), .A2(KEYINPUT44), .ZN(n352) );
  NAND2_X1 U433 ( .A1(n527), .A2(n350), .ZN(n627) );
  INV_X1 U434 ( .A(n724), .ZN(n350) );
  XNOR2_X1 U435 ( .A(n527), .B(KEYINPUT100), .ZN(n396) );
  XNOR2_X2 U436 ( .A(n449), .B(n351), .ZN(n527) );
  INV_X1 U437 ( .A(n448), .ZN(n351) );
  AND2_X1 U438 ( .A1(n633), .A2(n632), .ZN(n353) );
  XNOR2_X2 U439 ( .A(n354), .B(KEYINPUT45), .ZN(n754) );
  NAND2_X1 U440 ( .A1(n624), .A2(n636), .ZN(n357) );
  XNOR2_X1 U441 ( .A(n395), .B(n611), .ZN(n358) );
  BUF_X1 U442 ( .A(n595), .Z(n359) );
  XNOR2_X1 U443 ( .A(KEYINPUT15), .B(G902), .ZN(n468) );
  NOR2_X1 U444 ( .A1(n626), .A2(n538), .ZN(n539) );
  INV_X1 U445 ( .A(KEYINPUT78), .ZN(n420) );
  INV_X1 U446 ( .A(KEYINPUT89), .ZN(n376) );
  NOR2_X1 U447 ( .A1(n608), .A2(n699), .ZN(n609) );
  XOR2_X1 U448 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n461) );
  INV_X1 U449 ( .A(KEYINPUT71), .ZN(n452) );
  XNOR2_X2 U450 ( .A(KEYINPUT105), .B(KEYINPUT12), .ZN(n502) );
  INV_X1 U451 ( .A(KEYINPUT87), .ZN(n417) );
  INV_X1 U452 ( .A(G902), .ZN(n521) );
  INV_X1 U453 ( .A(G472), .ZN(n384) );
  NAND2_X1 U454 ( .A1(n369), .A2(n376), .ZN(n368) );
  INV_X1 U455 ( .A(KEYINPUT8), .ZN(n456) );
  XNOR2_X1 U456 ( .A(n413), .B(G122), .ZN(n514) );
  INV_X1 U457 ( .A(G134), .ZN(n387) );
  AND2_X1 U458 ( .A1(n556), .A2(n555), .ZN(n584) );
  INV_X1 U459 ( .A(G469), .ZN(n412) );
  XNOR2_X1 U460 ( .A(n591), .B(KEYINPUT115), .ZN(n556) );
  INV_X1 U461 ( .A(G140), .ZN(n562) );
  INV_X1 U462 ( .A(n597), .ZN(n700) );
  BUF_X1 U463 ( .A(n556), .Z(n702) );
  AND2_X1 U464 ( .A1(n408), .A2(n569), .ZN(n360) );
  XOR2_X1 U465 ( .A(KEYINPUT13), .B(G475), .Z(n361) );
  XOR2_X1 U466 ( .A(KEYINPUT113), .B(KEYINPUT6), .Z(n362) );
  AND2_X1 U467 ( .A1(n715), .A2(n527), .ZN(n363) );
  AND2_X2 U468 ( .A1(n553), .A2(n715), .ZN(n713) );
  XOR2_X1 U469 ( .A(n579), .B(KEYINPUT46), .Z(n365) );
  XNOR2_X1 U470 ( .A(KEYINPUT117), .B(KEYINPUT40), .ZN(n366) );
  XNOR2_X2 U471 ( .A(n367), .B(n496), .ZN(n647) );
  XNOR2_X1 U472 ( .A(n367), .B(n488), .ZN(n656) );
  XNOR2_X2 U473 ( .A(n764), .B(n483), .ZN(n367) );
  NAND2_X2 U474 ( .A1(n370), .A2(n368), .ZN(n769) );
  INV_X1 U475 ( .A(n358), .ZN(n369) );
  NOR2_X1 U476 ( .A1(n373), .A2(n372), .ZN(n371) );
  NAND2_X1 U477 ( .A1(n377), .A2(n375), .ZN(n374) );
  NOR2_X1 U478 ( .A1(n612), .A2(n376), .ZN(n375) );
  XNOR2_X1 U479 ( .A(n395), .B(n611), .ZN(n377) );
  XNOR2_X1 U480 ( .A(n453), .B(n452), .ZN(n454) );
  BUF_X1 U481 ( .A(n656), .Z(n378) );
  BUF_X1 U482 ( .A(n664), .Z(n379) );
  BUF_X1 U483 ( .A(n672), .Z(n380) );
  XNOR2_X1 U484 ( .A(n502), .B(n503), .ZN(n381) );
  NOR2_X1 U485 ( .A1(n672), .A2(n638), .ZN(n382) );
  XNOR2_X2 U486 ( .A(n385), .B(n384), .ZN(n564) );
  NOR2_X2 U487 ( .A1(n647), .A2(G902), .ZN(n385) );
  NAND2_X1 U488 ( .A1(n388), .A2(n389), .ZN(n518) );
  NAND2_X1 U489 ( .A1(n386), .A2(n387), .ZN(n389) );
  NAND2_X1 U490 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U491 ( .A1(n423), .A2(G134), .ZN(n388) );
  INV_X1 U492 ( .A(n423), .ZN(n386) );
  XNOR2_X1 U493 ( .A(n390), .B(KEYINPUT68), .ZN(n624) );
  NOR2_X2 U494 ( .A1(n616), .A2(KEYINPUT44), .ZN(n390) );
  INV_X1 U495 ( .A(n568), .ZN(n406) );
  NAND2_X1 U496 ( .A1(n568), .A2(n409), .ZN(n407) );
  BUF_X1 U497 ( .A(n616), .Z(n634) );
  XNOR2_X2 U498 ( .A(n484), .B(n391), .ZN(n400) );
  XNOR2_X2 U499 ( .A(n393), .B(n392), .ZN(n391) );
  XNOR2_X2 U500 ( .A(G122), .B(KEYINPUT74), .ZN(n392) );
  XNOR2_X2 U501 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n393) );
  XNOR2_X2 U502 ( .A(n394), .B(n430), .ZN(n484) );
  XNOR2_X2 U503 ( .A(G110), .B(G107), .ZN(n394) );
  NAND2_X1 U504 ( .A1(n396), .A2(n745), .ZN(n543) );
  AND2_X1 U505 ( .A1(n396), .A2(n499), .ZN(n693) );
  XNOR2_X1 U506 ( .A(n427), .B(n429), .ZN(n398) );
  XNOR2_X1 U507 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U508 ( .A(n426), .B(n460), .ZN(n397) );
  XNOR2_X1 U509 ( .A(n399), .B(n751), .ZN(n672) );
  XNOR2_X2 U510 ( .A(n400), .B(n494), .ZN(n751) );
  NAND2_X1 U511 ( .A1(n401), .A2(n402), .ZN(n581) );
  NAND2_X1 U512 ( .A1(n539), .A2(n401), .ZN(n541) );
  NOR2_X1 U513 ( .A1(n617), .A2(n401), .ZN(n618) );
  NOR2_X1 U514 ( .A1(n536), .A2(n401), .ZN(n537) );
  XNOR2_X2 U515 ( .A(n719), .B(n362), .ZN(n401) );
  INV_X1 U516 ( .A(n602), .ZN(n402) );
  NAND2_X1 U517 ( .A1(n403), .A2(n408), .ZN(n615) );
  AND2_X2 U518 ( .A1(n404), .A2(n407), .ZN(n403) );
  NAND2_X1 U519 ( .A1(n406), .A2(KEYINPUT39), .ZN(n405) );
  NAND2_X1 U520 ( .A1(n603), .A2(n409), .ZN(n408) );
  INV_X1 U521 ( .A(KEYINPUT39), .ZN(n409) );
  NOR2_X1 U522 ( .A1(n530), .A2(n563), .ZN(n415) );
  OR2_X1 U523 ( .A1(n538), .A2(n530), .ZN(n498) );
  INV_X1 U524 ( .A(n530), .ZN(n411) );
  XNOR2_X2 U525 ( .A(n489), .B(n412), .ZN(n530) );
  XNOR2_X1 U526 ( .A(n504), .B(n381), .ZN(n509) );
  NOR2_X2 U527 ( .A1(n664), .A2(G902), .ZN(n414) );
  NAND2_X1 U528 ( .A1(n415), .A2(n713), .ZN(n567) );
  NOR2_X2 U529 ( .A1(n566), .A2(n567), .ZN(n416) );
  XNOR2_X2 U530 ( .A(G143), .B(G128), .ZN(n423) );
  NAND2_X1 U531 ( .A1(n421), .A2(n419), .ZN(n418) );
  XNOR2_X2 U532 ( .A(n518), .B(n481), .ZN(n764) );
  XNOR2_X1 U533 ( .A(n418), .B(n417), .ZN(n640) );
  NAND2_X1 U534 ( .A1(n594), .A2(n359), .ZN(n597) );
  AND2_X2 U535 ( .A1(n688), .A2(G478), .ZN(n689) );
  BUF_X1 U536 ( .A(n683), .Z(n688) );
  XNOR2_X1 U537 ( .A(n547), .B(n546), .ZN(n616) );
  XOR2_X1 U538 ( .A(KEYINPUT66), .B(KEYINPUT19), .Z(n422) );
  INV_X1 U539 ( .A(KEYINPUT48), .ZN(n611) );
  XNOR2_X1 U540 ( .A(n455), .B(n454), .ZN(n459) );
  INV_X1 U541 ( .A(KEYINPUT65), .ZN(n641) );
  XNOR2_X2 U542 ( .A(KEYINPUT67), .B(G101), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n423), .B(n482), .ZN(n427) );
  XNOR2_X1 U544 ( .A(n425), .B(n424), .ZN(n426) );
  NAND2_X1 U545 ( .A1(n755), .A2(G224), .ZN(n428) );
  XNOR2_X1 U546 ( .A(n428), .B(KEYINPUT83), .ZN(n429) );
  XNOR2_X1 U547 ( .A(n432), .B(n431), .ZN(n494) );
  INV_X1 U548 ( .A(n468), .ZN(n638) );
  NAND2_X1 U549 ( .A1(n521), .A2(n433), .ZN(n435) );
  NAND2_X1 U550 ( .A1(n435), .A2(G210), .ZN(n434) );
  NAND2_X1 U551 ( .A1(n435), .A2(G214), .ZN(n436) );
  XNOR2_X1 U552 ( .A(n436), .B(KEYINPUT96), .ZN(n733) );
  INV_X1 U553 ( .A(n733), .ZN(n582) );
  NOR2_X2 U554 ( .A1(n560), .A2(n582), .ZN(n437) );
  XNOR2_X1 U555 ( .A(n437), .B(n422), .ZN(n595) );
  XNOR2_X1 U556 ( .A(n438), .B(KEYINPUT14), .ZN(n443) );
  NAND2_X1 U557 ( .A1(n443), .A2(G902), .ZN(n439) );
  XNOR2_X1 U558 ( .A(n439), .B(KEYINPUT99), .ZN(n548) );
  INV_X1 U559 ( .A(G898), .ZN(n440) );
  NAND2_X1 U560 ( .A1(n440), .A2(G953), .ZN(n442) );
  INV_X1 U561 ( .A(KEYINPUT98), .ZN(n441) );
  XNOR2_X1 U562 ( .A(n442), .B(n441), .ZN(n752) );
  NAND2_X1 U563 ( .A1(n548), .A2(n752), .ZN(n445) );
  NAND2_X1 U564 ( .A1(G952), .A2(n443), .ZN(n743) );
  NOR2_X1 U565 ( .A1(G953), .A2(n743), .ZN(n444) );
  XNOR2_X1 U566 ( .A(n444), .B(KEYINPUT97), .ZN(n552) );
  NAND2_X1 U567 ( .A1(n445), .A2(n552), .ZN(n446) );
  NAND2_X1 U568 ( .A1(n595), .A2(n446), .ZN(n449) );
  INV_X1 U569 ( .A(KEYINPUT93), .ZN(n447) );
  XNOR2_X1 U570 ( .A(n447), .B(KEYINPUT0), .ZN(n448) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n451) );
  XNOR2_X1 U572 ( .A(G119), .B(G128), .ZN(n450) );
  XNOR2_X1 U573 ( .A(n451), .B(n450), .ZN(n455) );
  NAND2_X1 U574 ( .A1(n755), .A2(G234), .ZN(n457) );
  XNOR2_X1 U575 ( .A(n457), .B(n456), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n516), .A2(G221), .ZN(n458) );
  XNOR2_X1 U577 ( .A(n459), .B(n458), .ZN(n465) );
  INV_X1 U578 ( .A(n465), .ZN(n464) );
  XNOR2_X1 U579 ( .A(n460), .B(n562), .ZN(n462) );
  XNOR2_X1 U580 ( .A(n462), .B(n461), .ZN(n767) );
  INV_X1 U581 ( .A(n767), .ZN(n463) );
  NAND2_X1 U582 ( .A1(n464), .A2(n463), .ZN(n467) );
  NAND2_X1 U583 ( .A1(n465), .A2(n767), .ZN(n466) );
  NAND2_X1 U584 ( .A1(n467), .A2(n466), .ZN(n681) );
  NAND2_X1 U585 ( .A1(n681), .A2(n521), .ZN(n476) );
  NAND2_X1 U586 ( .A1(n468), .A2(G234), .ZN(n469) );
  XNOR2_X1 U587 ( .A(n469), .B(KEYINPUT102), .ZN(n470) );
  XNOR2_X1 U588 ( .A(KEYINPUT20), .B(n470), .ZN(n477) );
  NAND2_X1 U589 ( .A1(G217), .A2(n477), .ZN(n474) );
  XOR2_X1 U590 ( .A(KEYINPUT25), .B(KEYINPUT82), .Z(n472) );
  XNOR2_X1 U591 ( .A(KEYINPUT101), .B(KEYINPUT103), .ZN(n471) );
  XNOR2_X1 U592 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U593 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U594 ( .A1(n477), .A2(G221), .ZN(n479) );
  INV_X1 U595 ( .A(KEYINPUT21), .ZN(n478) );
  XNOR2_X1 U596 ( .A(n479), .B(n478), .ZN(n715) );
  XNOR2_X1 U597 ( .A(n480), .B(KEYINPUT4), .ZN(n481) );
  XNOR2_X1 U598 ( .A(n482), .B(G146), .ZN(n483) );
  INV_X1 U599 ( .A(n484), .ZN(n487) );
  NAND2_X1 U600 ( .A1(n755), .A2(G227), .ZN(n485) );
  XNOR2_X1 U601 ( .A(n485), .B(G140), .ZN(n486) );
  XNOR2_X1 U602 ( .A(n487), .B(n486), .ZN(n488) );
  OR2_X2 U603 ( .A1(n656), .A2(G902), .ZN(n489) );
  INV_X1 U604 ( .A(G953), .ZN(n490) );
  NAND2_X1 U605 ( .A1(n490), .A2(n433), .ZN(n491) );
  NAND2_X1 U606 ( .A1(n505), .A2(G210), .ZN(n493) );
  XNOR2_X1 U607 ( .A(KEYINPUT77), .B(KEYINPUT5), .ZN(n492) );
  XNOR2_X1 U608 ( .A(n493), .B(n492), .ZN(n495) );
  XNOR2_X1 U609 ( .A(n495), .B(n494), .ZN(n496) );
  BUF_X1 U610 ( .A(n564), .Z(n497) );
  NOR2_X1 U611 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U612 ( .A(n501), .B(n500), .ZN(n504) );
  XNOR2_X2 U613 ( .A(G131), .B(KEYINPUT107), .ZN(n503) );
  NAND2_X1 U614 ( .A1(n505), .A2(G214), .ZN(n507) );
  XNOR2_X1 U615 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n510), .B(n767), .ZN(n664) );
  XNOR2_X1 U618 ( .A(n525), .B(KEYINPUT108), .ZN(n589) );
  XOR2_X1 U619 ( .A(KEYINPUT109), .B(KEYINPUT7), .Z(n512) );
  XNOR2_X1 U620 ( .A(n512), .B(n511), .ZN(n513) );
  NAND2_X1 U621 ( .A1(n516), .A2(G217), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U623 ( .A(n520), .B(n519), .ZN(n690) );
  NAND2_X1 U624 ( .A1(n690), .A2(n521), .ZN(n522) );
  NAND2_X1 U625 ( .A1(n693), .A2(n702), .ZN(n524) );
  XNOR2_X1 U626 ( .A(n524), .B(G104), .ZN(G6) );
  INV_X1 U627 ( .A(n525), .ZN(n544) );
  NOR2_X2 U628 ( .A1(n544), .A2(n590), .ZN(n526) );
  NAND2_X1 U629 ( .A1(n734), .A2(n363), .ZN(n529) );
  XNOR2_X1 U630 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n528) );
  XNOR2_X2 U631 ( .A(n530), .B(KEYINPUT1), .ZN(n626) );
  INV_X1 U632 ( .A(n553), .ZN(n535) );
  INV_X1 U633 ( .A(n535), .ZN(n716) );
  NOR2_X1 U634 ( .A1(n497), .A2(n716), .ZN(n531) );
  AND2_X1 U635 ( .A1(n626), .A2(n531), .ZN(n532) );
  NAND2_X1 U636 ( .A1(n619), .A2(n532), .ZN(n623) );
  XOR2_X1 U637 ( .A(G110), .B(KEYINPUT119), .Z(n533) );
  XNOR2_X1 U638 ( .A(n623), .B(n533), .ZN(G12) );
  INV_X1 U639 ( .A(n626), .ZN(n534) );
  OR2_X1 U640 ( .A1(n534), .A2(n535), .ZN(n536) );
  INV_X1 U641 ( .A(n564), .ZN(n719) );
  NAND2_X1 U642 ( .A1(n619), .A2(n537), .ZN(n632) );
  XNOR2_X1 U643 ( .A(n632), .B(G101), .ZN(G3) );
  INV_X1 U644 ( .A(n713), .ZN(n538) );
  XNOR2_X1 U645 ( .A(KEYINPUT94), .B(KEYINPUT33), .ZN(n540) );
  INV_X1 U646 ( .A(KEYINPUT34), .ZN(n542) );
  XNOR2_X1 U647 ( .A(n543), .B(n542), .ZN(n545) );
  AND2_X1 U648 ( .A1(n590), .A2(n544), .ZN(n606) );
  NAND2_X1 U649 ( .A1(n545), .A2(n606), .ZN(n547) );
  XOR2_X1 U650 ( .A(n634), .B(G122), .Z(G24) );
  INV_X1 U651 ( .A(G900), .ZN(n550) );
  AND2_X1 U652 ( .A1(G953), .A2(n548), .ZN(n549) );
  NAND2_X1 U653 ( .A1(n550), .A2(n549), .ZN(n551) );
  AND2_X1 U654 ( .A1(n552), .A2(n551), .ZN(n563) );
  NOR2_X1 U655 ( .A1(n563), .A2(n553), .ZN(n554) );
  NAND2_X1 U656 ( .A1(n715), .A2(n554), .ZN(n573) );
  INV_X1 U657 ( .A(n573), .ZN(n555) );
  INV_X1 U658 ( .A(KEYINPUT43), .ZN(n558) );
  XNOR2_X1 U659 ( .A(n559), .B(n558), .ZN(n561) );
  BUF_X2 U660 ( .A(n560), .Z(n602) );
  XNOR2_X1 U661 ( .A(n612), .B(n562), .ZN(G42) );
  NAND2_X1 U662 ( .A1(n564), .A2(n733), .ZN(n565) );
  INV_X1 U663 ( .A(n731), .ZN(n568) );
  INV_X1 U664 ( .A(n591), .ZN(n569) );
  NAND2_X1 U665 ( .A1(n570), .A2(n734), .ZN(n572) );
  XNOR2_X1 U666 ( .A(KEYINPUT118), .B(KEYINPUT41), .ZN(n571) );
  XNOR2_X2 U667 ( .A(n572), .B(n571), .ZN(n744) );
  INV_X1 U668 ( .A(KEYINPUT28), .ZN(n574) );
  NAND2_X2 U669 ( .A1(n744), .A2(n594), .ZN(n577) );
  XNOR2_X2 U670 ( .A(n577), .B(KEYINPUT42), .ZN(n778) );
  INV_X1 U671 ( .A(n778), .ZN(n578) );
  INV_X1 U672 ( .A(KEYINPUT64), .ZN(n579) );
  XNOR2_X1 U673 ( .A(n580), .B(n365), .ZN(n610) );
  NOR2_X1 U674 ( .A1(n582), .A2(n581), .ZN(n583) );
  AND2_X1 U675 ( .A1(n584), .A2(n583), .ZN(n587) );
  INV_X1 U676 ( .A(KEYINPUT90), .ZN(n585) );
  XOR2_X1 U677 ( .A(n585), .B(KEYINPUT36), .Z(n586) );
  XNOR2_X1 U678 ( .A(n587), .B(n586), .ZN(n588) );
  NAND2_X1 U679 ( .A1(n588), .A2(n534), .ZN(n707) );
  AND2_X1 U680 ( .A1(n590), .A2(n589), .ZN(n704) );
  INV_X1 U681 ( .A(n704), .ZN(n614) );
  AND2_X1 U682 ( .A1(n591), .A2(n614), .ZN(n629) );
  XOR2_X1 U683 ( .A(KEYINPUT69), .B(KEYINPUT47), .Z(n592) );
  NOR2_X1 U684 ( .A1(n629), .A2(n592), .ZN(n593) );
  XNOR2_X1 U685 ( .A(KEYINPUT76), .B(n593), .ZN(n596) );
  AND2_X1 U686 ( .A1(n596), .A2(n700), .ZN(n600) );
  NAND2_X1 U687 ( .A1(n707), .A2(n601), .ZN(n608) );
  OR2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n605) );
  INV_X1 U689 ( .A(KEYINPUT116), .ZN(n604) );
  XNOR2_X1 U690 ( .A(n605), .B(n604), .ZN(n607) );
  AND2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n699) );
  INV_X1 U692 ( .A(n612), .ZN(n613) );
  OR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n678) );
  OR2_X1 U694 ( .A1(n626), .A2(n716), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n622) );
  INV_X1 U696 ( .A(KEYINPUT85), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n620), .B(KEYINPUT32), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n622), .B(n621), .ZN(n679) );
  NAND2_X1 U699 ( .A1(n713), .A2(n497), .ZN(n625) );
  OR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n724) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT31), .ZN(n705) );
  XNOR2_X1 U702 ( .A(n628), .B(KEYINPUT104), .ZN(n630) );
  INV_X1 U703 ( .A(n629), .ZN(n728) );
  NAND2_X1 U704 ( .A1(n630), .A2(n728), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n631), .B(KEYINPUT112), .ZN(n633) );
  INV_X1 U706 ( .A(n634), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n638), .A2(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n642), .B(n641), .ZN(n646) );
  INV_X1 U710 ( .A(n769), .ZN(n643) );
  AND2_X1 U711 ( .A1(n754), .A2(n643), .ZN(n709) );
  NAND2_X1 U712 ( .A1(n709), .A2(KEYINPUT2), .ZN(n644) );
  XOR2_X1 U713 ( .A(KEYINPUT80), .B(n644), .Z(n711) );
  INV_X1 U714 ( .A(n711), .ZN(n645) );
  AND2_X2 U715 ( .A1(n646), .A2(n645), .ZN(n683) );
  NAND2_X1 U716 ( .A1(n683), .A2(G472), .ZN(n650) );
  BUF_X1 U717 ( .A(n647), .Z(n648) );
  XNOR2_X1 U718 ( .A(n650), .B(n649), .ZN(n652) );
  INV_X1 U719 ( .A(G952), .ZN(n651) );
  NAND2_X1 U720 ( .A1(n652), .A2(n686), .ZN(n654) );
  XOR2_X1 U721 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(G57) );
  NAND2_X1 U723 ( .A1(n683), .A2(G469), .ZN(n658) );
  XNOR2_X1 U724 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n659), .A2(n686), .ZN(n661) );
  INV_X1 U727 ( .A(KEYINPUT122), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n661), .B(n660), .ZN(G54) );
  NAND2_X1 U729 ( .A1(n683), .A2(G475), .ZN(n666) );
  XNOR2_X1 U730 ( .A(KEYINPUT95), .B(KEYINPUT123), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT59), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U733 ( .A1(n667), .A2(n686), .ZN(n669) );
  INV_X1 U734 ( .A(KEYINPUT60), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n669), .B(n668), .ZN(G60) );
  NAND2_X1 U736 ( .A1(n683), .A2(G210), .ZN(n674) );
  XNOR2_X1 U737 ( .A(KEYINPUT92), .B(KEYINPUT54), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n670), .B(KEYINPUT55), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U740 ( .A1(n675), .A2(n686), .ZN(n677) );
  INV_X1 U741 ( .A(KEYINPUT56), .ZN(n676) );
  XNOR2_X1 U742 ( .A(n677), .B(n676), .ZN(G51) );
  XNOR2_X1 U743 ( .A(n678), .B(G134), .ZN(G36) );
  XNOR2_X1 U744 ( .A(n679), .B(G119), .ZN(G21) );
  XOR2_X1 U745 ( .A(n680), .B(G131), .Z(G33) );
  BUF_X1 U746 ( .A(n681), .Z(n682) );
  INV_X1 U747 ( .A(n682), .ZN(n685) );
  NAND2_X1 U748 ( .A1(n688), .A2(G217), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n685), .B(n684), .ZN(n687) );
  INV_X1 U750 ( .A(n686), .ZN(n691) );
  NOR2_X1 U751 ( .A1(n687), .A2(n691), .ZN(G66) );
  XNOR2_X1 U752 ( .A(n689), .B(n690), .ZN(n692) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(G63) );
  NAND2_X1 U754 ( .A1(n693), .A2(n704), .ZN(n695) );
  XOR2_X1 U755 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n694) );
  XNOR2_X1 U756 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U757 ( .A(n413), .B(n696), .ZN(G9) );
  XOR2_X1 U758 ( .A(G128), .B(KEYINPUT29), .Z(n698) );
  NAND2_X1 U759 ( .A1(n700), .A2(n704), .ZN(n697) );
  XNOR2_X1 U760 ( .A(n698), .B(n697), .ZN(G30) );
  XOR2_X1 U761 ( .A(G143), .B(n699), .Z(G45) );
  NAND2_X1 U762 ( .A1(n702), .A2(n700), .ZN(n701) );
  XNOR2_X1 U763 ( .A(n701), .B(G146), .ZN(G48) );
  NAND2_X1 U764 ( .A1(n705), .A2(n702), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n703), .B(G113), .ZN(G15) );
  NAND2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U767 ( .A(n706), .B(G116), .ZN(G18) );
  XOR2_X1 U768 ( .A(n707), .B(G125), .Z(n708) );
  XNOR2_X1 U769 ( .A(n708), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U770 ( .A1(n709), .A2(KEYINPUT2), .ZN(n710) );
  NOR2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U772 ( .A1(n712), .A2(G953), .ZN(n749) );
  NOR2_X1 U773 ( .A1(n534), .A2(n713), .ZN(n714) );
  XNOR2_X1 U774 ( .A(n714), .B(KEYINPUT50), .ZN(n722) );
  NOR2_X1 U775 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U776 ( .A(KEYINPUT120), .B(KEYINPUT49), .ZN(n717) );
  XNOR2_X1 U777 ( .A(n718), .B(n717), .ZN(n720) );
  NAND2_X1 U778 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U780 ( .A(n723), .B(KEYINPUT121), .ZN(n725) );
  NAND2_X1 U781 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U782 ( .A(KEYINPUT51), .B(n726), .Z(n727) );
  NAND2_X1 U783 ( .A1(n727), .A2(n744), .ZN(n740) );
  INV_X1 U784 ( .A(n734), .ZN(n730) );
  NAND2_X1 U785 ( .A1(n728), .A2(n733), .ZN(n729) );
  NAND2_X1 U786 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U787 ( .A1(n732), .A2(n406), .ZN(n737) );
  AND2_X1 U788 ( .A1(n734), .A2(n733), .ZN(n735) );
  INV_X1 U789 ( .A(n735), .ZN(n736) );
  NAND2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U791 ( .A1(n745), .A2(n738), .ZN(n739) );
  NAND2_X1 U792 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U793 ( .A(KEYINPUT52), .B(n741), .Z(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n747) );
  AND2_X1 U795 ( .A1(n744), .A2(n745), .ZN(n746) );
  NOR2_X1 U796 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U798 ( .A(KEYINPUT53), .B(n750), .Z(G75) );
  XNOR2_X1 U799 ( .A(n751), .B(G101), .ZN(n753) );
  NOR2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n763) );
  BUF_X1 U801 ( .A(n754), .Z(n756) );
  NAND2_X1 U802 ( .A1(n756), .A2(n755), .ZN(n761) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n757) );
  XNOR2_X1 U804 ( .A(KEYINPUT61), .B(n757), .ZN(n758) );
  NAND2_X1 U805 ( .A1(n758), .A2(G898), .ZN(n759) );
  XNOR2_X1 U806 ( .A(n759), .B(KEYINPUT124), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U808 ( .A(n763), .B(n762), .ZN(G69) );
  INV_X1 U809 ( .A(n764), .ZN(n765) );
  INV_X1 U810 ( .A(n765), .ZN(n766) );
  XOR2_X1 U811 ( .A(n767), .B(n766), .Z(n771) );
  XNOR2_X1 U812 ( .A(n771), .B(KEYINPUT125), .ZN(n768) );
  XNOR2_X1 U813 ( .A(n769), .B(n768), .ZN(n770) );
  NOR2_X1 U814 ( .A1(G953), .A2(n770), .ZN(n776) );
  XNOR2_X1 U815 ( .A(n771), .B(G227), .ZN(n772) );
  NAND2_X1 U816 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U817 ( .A1(G953), .A2(n773), .ZN(n774) );
  XOR2_X1 U818 ( .A(KEYINPUT126), .B(n774), .Z(n775) );
  NOR2_X1 U819 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U820 ( .A(KEYINPUT127), .B(n777), .ZN(G72) );
  XNOR2_X1 U821 ( .A(n778), .B(G137), .ZN(G39) );
endmodule

