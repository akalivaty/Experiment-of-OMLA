

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X2 U325 ( .A(n454), .B(KEYINPUT122), .ZN(n565) );
  NOR2_X2 U326 ( .A1(n453), .A2(n537), .ZN(n454) );
  XOR2_X1 U327 ( .A(KEYINPUT36), .B(n544), .Z(n583) );
  INV_X1 U328 ( .A(KEYINPUT68), .ZN(n326) );
  NOR2_X1 U329 ( .A1(n394), .A2(n563), .ZN(n395) );
  XNOR2_X1 U330 ( .A(n414), .B(n293), .ZN(n433) );
  XNOR2_X1 U331 ( .A(n347), .B(n346), .ZN(n504) );
  XNOR2_X1 U332 ( .A(n345), .B(n344), .ZN(n346) );
  BUF_X1 U333 ( .A(n391), .Z(n544) );
  XNOR2_X1 U334 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U336 ( .A(n367), .B(n366), .ZN(n387) );
  XNOR2_X1 U337 ( .A(n392), .B(KEYINPUT45), .ZN(n393) );
  INV_X1 U338 ( .A(KEYINPUT67), .ZN(n338) );
  XNOR2_X1 U339 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U340 ( .A(n380), .B(n340), .ZN(n341) );
  INV_X1 U341 ( .A(n521), .ZN(n432) );
  XNOR2_X1 U342 ( .A(n327), .B(n326), .ZN(n328) );
  NAND2_X1 U343 ( .A1(n433), .A2(n432), .ZN(n434) );
  XNOR2_X1 U344 ( .A(n329), .B(n328), .ZN(n345) );
  XNOR2_X1 U345 ( .A(n434), .B(KEYINPUT64), .ZN(n568) );
  XOR2_X1 U346 ( .A(KEYINPUT94), .B(n472), .Z(n521) );
  XNOR2_X1 U347 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U348 ( .A(G78GAT), .B(KEYINPUT87), .Z(n295) );
  XNOR2_X1 U349 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U351 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n297) );
  XNOR2_X1 U352 ( .A(KEYINPUT86), .B(KEYINPUT91), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U354 ( .A(n299), .B(n298), .Z(n311) );
  XNOR2_X1 U355 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n300), .B(KEYINPUT3), .ZN(n301) );
  XOR2_X1 U357 ( .A(n301), .B(KEYINPUT90), .Z(n303) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(G148GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n431) );
  XOR2_X1 U360 ( .A(G162GAT), .B(G106GAT), .Z(n305) );
  XNOR2_X1 U361 ( .A(G50GAT), .B(G218GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(KEYINPUT88), .B(n306), .Z(n308) );
  NAND2_X1 U364 ( .A1(G228GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n431), .B(n309), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U368 ( .A(KEYINPUT21), .B(G211GAT), .Z(n313) );
  XNOR2_X1 U369 ( .A(KEYINPUT89), .B(G204GAT), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(n314), .ZN(n412) );
  XNOR2_X1 U372 ( .A(n315), .B(n412), .ZN(n475) );
  XOR2_X1 U373 ( .A(G190GAT), .B(G218GAT), .Z(n401) );
  AND2_X1 U374 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n401), .B(n316), .ZN(n318) );
  XNOR2_X1 U376 ( .A(G134GAT), .B(G162GAT), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n317), .B(KEYINPUT77), .ZN(n421) );
  XNOR2_X1 U378 ( .A(n318), .B(n421), .ZN(n319) );
  XOR2_X1 U379 ( .A(n319), .B(KEYINPUT78), .Z(n323) );
  XOR2_X1 U380 ( .A(G85GAT), .B(G92GAT), .Z(n321) );
  XNOR2_X1 U381 ( .A(G99GAT), .B(G106GAT), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n351) );
  XNOR2_X1 U383 ( .A(n351), .B(KEYINPUT10), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n334) );
  XOR2_X1 U385 ( .A(G43GAT), .B(G29GAT), .Z(n325) );
  XNOR2_X1 U386 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n329) );
  XNOR2_X1 U388 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n327) );
  XOR2_X1 U389 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n331) );
  XNOR2_X1 U390 ( .A(KEYINPUT76), .B(KEYINPUT65), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U392 ( .A(n345), .B(n332), .Z(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n561) );
  XOR2_X1 U394 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n336) );
  XNOR2_X1 U395 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U397 ( .A(G169GAT), .B(G8GAT), .Z(n409) );
  XNOR2_X1 U398 ( .A(n337), .B(n409), .ZN(n342) );
  XOR2_X1 U399 ( .A(G15GAT), .B(G22GAT), .Z(n380) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U402 ( .A(G113GAT), .B(G1GAT), .Z(n418) );
  XOR2_X1 U403 ( .A(n343), .B(n418), .Z(n347) );
  XNOR2_X1 U404 ( .A(G197GAT), .B(G141GAT), .ZN(n344) );
  INV_X1 U405 ( .A(n504), .ZN(n569) );
  XOR2_X1 U406 ( .A(G176GAT), .B(G64GAT), .Z(n408) );
  XOR2_X1 U407 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n349) );
  XNOR2_X1 U408 ( .A(G71GAT), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n368) );
  XNOR2_X1 U410 ( .A(n408), .B(n368), .ZN(n350) );
  XOR2_X1 U411 ( .A(G120GAT), .B(G57GAT), .Z(n417) );
  XNOR2_X1 U412 ( .A(n350), .B(n417), .ZN(n355) );
  XOR2_X1 U413 ( .A(n351), .B(KEYINPUT33), .Z(n353) );
  NAND2_X1 U414 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n363) );
  XOR2_X1 U417 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n357) );
  XNOR2_X1 U418 ( .A(G204GAT), .B(G148GAT), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U420 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n359) );
  XNOR2_X1 U421 ( .A(KEYINPUT32), .B(KEYINPUT74), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U423 ( .A(n361), .B(n360), .Z(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n573) );
  XNOR2_X1 U425 ( .A(n573), .B(KEYINPUT41), .ZN(n555) );
  NAND2_X1 U426 ( .A1(n569), .A2(n555), .ZN(n367) );
  XOR2_X1 U427 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n365) );
  INV_X1 U428 ( .A(KEYINPUT114), .ZN(n364) );
  XOR2_X1 U429 ( .A(n368), .B(KEYINPUT81), .Z(n370) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n386) );
  XOR2_X1 U432 ( .A(KEYINPUT82), .B(G57GAT), .Z(n372) );
  XNOR2_X1 U433 ( .A(G1GAT), .B(G64GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U435 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n374) );
  XNOR2_X1 U436 ( .A(KEYINPUT12), .B(KEYINPUT83), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n384) );
  XOR2_X1 U439 ( .A(G155GAT), .B(G211GAT), .Z(n378) );
  XNOR2_X1 U440 ( .A(G183GAT), .B(G127GAT), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U442 ( .A(n379), .B(KEYINPUT80), .Z(n382) );
  XNOR2_X1 U443 ( .A(G8GAT), .B(n380), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n492) );
  INV_X1 U447 ( .A(n492), .ZN(n577) );
  NOR2_X1 U448 ( .A1(n387), .A2(n577), .ZN(n388) );
  XOR2_X1 U449 ( .A(KEYINPUT116), .B(n388), .Z(n389) );
  NOR2_X1 U450 ( .A1(n561), .A2(n389), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n390), .B(KEYINPUT47), .ZN(n397) );
  XOR2_X1 U452 ( .A(KEYINPUT79), .B(n561), .Z(n391) );
  NOR2_X1 U453 ( .A1(n583), .A2(n492), .ZN(n392) );
  NAND2_X1 U454 ( .A1(n393), .A2(n573), .ZN(n394) );
  XNOR2_X1 U455 ( .A(KEYINPUT70), .B(n569), .ZN(n563) );
  XNOR2_X1 U456 ( .A(n395), .B(KEYINPUT117), .ZN(n396) );
  NAND2_X1 U457 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X2 U458 ( .A(n398), .B(KEYINPUT48), .ZN(n550) );
  XOR2_X1 U459 ( .A(G183GAT), .B(KEYINPUT17), .Z(n400) );
  XNOR2_X1 U460 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n438) );
  XOR2_X1 U462 ( .A(n401), .B(n438), .Z(n403) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U465 ( .A(KEYINPUT80), .B(KEYINPUT95), .Z(n405) );
  XNOR2_X1 U466 ( .A(G36GAT), .B(G92GAT), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U468 ( .A(n407), .B(n406), .Z(n411) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n524) );
  NAND2_X1 U472 ( .A1(n550), .A2(n524), .ZN(n414) );
  XOR2_X1 U473 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n416) );
  XNOR2_X1 U474 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n429) );
  XOR2_X1 U476 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n420) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n425) );
  XOR2_X1 U479 ( .A(KEYINPUT0), .B(G127GAT), .Z(n439) );
  XOR2_X1 U480 ( .A(n421), .B(n439), .Z(n423) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U483 ( .A(n425), .B(n424), .Z(n427) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(G85GAT), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U486 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n472) );
  NOR2_X1 U488 ( .A1(n475), .A2(n568), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n435), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n437) );
  XNOR2_X1 U491 ( .A(G190GAT), .B(G134GAT), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n452) );
  XOR2_X1 U493 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G99GAT), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT85), .B(G120GAT), .Z(n443) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n450) );
  XOR2_X1 U500 ( .A(G71GAT), .B(G176GAT), .Z(n447) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(G15GAT), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U503 ( .A(G113GAT), .B(n448), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n537) );
  NAND2_X1 U506 ( .A1(n565), .A2(n544), .ZN(n458) );
  XOR2_X1 U507 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n456) );
  INV_X1 U508 ( .A(G190GAT), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  NAND2_X1 U510 ( .A1(n565), .A2(n555), .ZN(n462) );
  XOR2_X1 U511 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n460) );
  XOR2_X1 U512 ( .A(G176GAT), .B(KEYINPUT56), .Z(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n462), .B(n461), .ZN(G1349GAT) );
  XNOR2_X1 U515 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(KEYINPUT34), .ZN(n464) );
  XOR2_X1 U517 ( .A(KEYINPUT98), .B(n464), .Z(n481) );
  NAND2_X1 U518 ( .A1(n573), .A2(n563), .ZN(n495) );
  NOR2_X1 U519 ( .A1(n544), .A2(n492), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n465), .B(KEYINPUT16), .ZN(n479) );
  INV_X1 U521 ( .A(n537), .ZN(n528) );
  AND2_X1 U522 ( .A1(n528), .A2(n524), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n475), .A2(n466), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT25), .ZN(n471) );
  XNOR2_X1 U525 ( .A(n524), .B(KEYINPUT27), .ZN(n474) );
  XOR2_X1 U526 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n469) );
  NAND2_X1 U527 ( .A1(n475), .A2(n537), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(n567) );
  INV_X1 U529 ( .A(n567), .ZN(n549) );
  NAND2_X1 U530 ( .A1(n474), .A2(n549), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n472), .ZN(n478) );
  NAND2_X1 U533 ( .A1(n521), .A2(n474), .ZN(n552) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT28), .ZN(n532) );
  NOR2_X1 U535 ( .A1(n552), .A2(n532), .ZN(n535) );
  XNOR2_X1 U536 ( .A(n535), .B(KEYINPUT96), .ZN(n476) );
  NAND2_X1 U537 ( .A1(n476), .A2(n537), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n478), .A2(n477), .ZN(n491) );
  NAND2_X1 U539 ( .A1(n479), .A2(n491), .ZN(n506) );
  NOR2_X1 U540 ( .A1(n495), .A2(n506), .ZN(n487) );
  NAND2_X1 U541 ( .A1(n487), .A2(n521), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n487), .A2(n524), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(KEYINPUT100), .ZN(n483) );
  XNOR2_X1 U545 ( .A(G8GAT), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U547 ( .A1(n487), .A2(n528), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U549 ( .A(G15GAT), .B(n486), .Z(G1326GAT) );
  NAND2_X1 U550 ( .A1(n532), .A2(n487), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n490) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n498) );
  NAND2_X1 U555 ( .A1(n492), .A2(n491), .ZN(n493) );
  NOR2_X1 U556 ( .A1(n493), .A2(n583), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n494), .B(KEYINPUT37), .ZN(n519) );
  NOR2_X1 U558 ( .A1(n495), .A2(n519), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT38), .ZN(n502) );
  NAND2_X1 U560 ( .A1(n502), .A2(n521), .ZN(n497) );
  XOR2_X1 U561 ( .A(n498), .B(n497), .Z(G1328GAT) );
  NAND2_X1 U562 ( .A1(n502), .A2(n524), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U564 ( .A1(n502), .A2(n528), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(KEYINPUT40), .ZN(n501) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U567 ( .A1(n502), .A2(n532), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U569 ( .A1(n555), .A2(n504), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(KEYINPUT104), .ZN(n520) );
  NOR2_X1 U571 ( .A1(n520), .A2(n506), .ZN(n507) );
  XOR2_X1 U572 ( .A(KEYINPUT105), .B(n507), .Z(n514) );
  NAND2_X1 U573 ( .A1(n521), .A2(n514), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(KEYINPUT42), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n524), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(KEYINPUT106), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(n511), .ZN(G1333GAT) );
  XOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT107), .Z(n513) );
  NAND2_X1 U580 ( .A1(n514), .A2(n528), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U583 ( .A1(n514), .A2(n532), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT109), .Z(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n523) );
  NOR2_X1 U588 ( .A1(n520), .A2(n519), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n531), .A2(n521), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(G1336GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n526) );
  NAND2_X1 U592 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  XOR2_X1 U595 ( .A(G99GAT), .B(KEYINPUT113), .Z(n530) );
  NAND2_X1 U596 ( .A1(n531), .A2(n528), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n550), .A2(n535), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n563), .A2(n545), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT118), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U607 ( .A1(n545), .A2(n555), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n545), .A2(n577), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n547) );
  NAND2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT120), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n569), .A2(n560), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n560), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n577), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n565), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n577), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n578), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U639 ( .A(n578), .ZN(n582) );
  OR2_X1 U640 ( .A1(n582), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n581) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n585) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(n585), .B(n584), .Z(G1355GAT) );
endmodule

