//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G148gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(G148gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(KEYINPUT74), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n205), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT75), .B(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n202), .B1(new_n204), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(new_n218), .B2(new_n204), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n211), .B2(new_n208), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n214), .A2(new_n217), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT67), .B(G120gat), .Z(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT68), .B(G113gat), .ZN(new_n228));
  INV_X1    g027(.A(G120gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n226), .A2(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(G127gat), .A2(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(G127gat), .A2(G134gat), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT1), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT1), .B1(new_n227), .B2(new_n229), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n227), .B2(new_n229), .ZN(new_n236));
  INV_X1    g035(.A(G127gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT66), .B(G134gat), .Z(new_n238));
  OAI211_X1 g037(.A(new_n236), .B(new_n231), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n223), .A2(new_n224), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n234), .A2(new_n239), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n223), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT77), .B1(new_n247), .B2(KEYINPUT4), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n214), .A2(new_n217), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n220), .A2(new_n222), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(new_n240), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n253));
  OAI21_X1  g052(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n247), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n245), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G225gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n247), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n253), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n252), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n260), .B(new_n262), .C1(new_n242), .C2(new_n241), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n263), .B2(new_n244), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n251), .A2(new_n240), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n247), .A2(KEYINPUT78), .A3(new_n266), .ZN(new_n267));
  OR3_X1    g066(.A1(new_n246), .A2(KEYINPUT78), .A3(new_n223), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n257), .A2(new_n244), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G1gat), .B(G29gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT0), .ZN(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G85gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n271), .B1(new_n256), .B2(new_n264), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT6), .B1(new_n280), .B2(new_n277), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(KEYINPUT6), .A3(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G211gat), .A2(G218gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT22), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G197gat), .ZN(new_n288));
  INV_X1    g087(.A(G204gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G211gat), .B(G218gat), .Z(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n294), .A2(new_n295), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G226gat), .ZN(new_n300));
  INV_X1    g099(.A(G233gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT27), .B(G183gat), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT26), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n316), .A2(new_n311), .A3(KEYINPUT26), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(KEYINPUT23), .B2(new_n311), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n325));
  MUX2_X1   g124(.A(G183gat), .B(new_n325), .S(G190gat), .Z(new_n326));
  INV_X1    g125(.A(new_n310), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(KEYINPUT24), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT24), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(KEYINPUT65), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT65), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n310), .B1(new_n333), .B2(KEYINPUT24), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n326), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n323), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT64), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n320), .B(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n321), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n304), .B1(new_n330), .B2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n309), .A2(new_n318), .B1(new_n324), .B2(new_n328), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n320), .B(KEYINPUT64), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT25), .B1(new_n343), .B2(new_n336), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(KEYINPUT72), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n303), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n302), .A2(KEYINPUT29), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n330), .B2(new_n340), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n299), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n341), .A2(new_n347), .A3(new_n345), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n330), .A2(new_n340), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n302), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n350), .A2(new_n357), .A3(new_n361), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(KEYINPUT30), .A3(new_n364), .ZN(new_n365));
  OR3_X1    g164(.A1(new_n358), .A2(KEYINPUT30), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n284), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n299), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n224), .B1(new_n370), .B2(KEYINPUT29), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n371), .B2(new_n251), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT29), .B1(new_n223), .B2(new_n224), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n374), .A3(new_n353), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT80), .B(G22gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n378));
  INV_X1    g177(.A(new_n292), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n379), .A2(new_n295), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n379), .B2(new_n295), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n224), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n251), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(new_n373), .B2(new_n299), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n378), .B1(new_n385), .B2(new_n369), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n378), .A3(new_n369), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n376), .B(new_n377), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G78gat), .B(G106gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT31), .B(G50gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G22gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n376), .B1(new_n388), .B2(new_n386), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(KEYINPUT81), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n385), .A2(new_n369), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT79), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n399), .A2(new_n387), .B1(new_n375), .B2(new_n372), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n394), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n377), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n393), .B1(new_n405), .B2(new_n389), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT82), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(G22gat), .B1(new_n400), .B2(new_n401), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n389), .B(new_n393), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n389), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n392), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n368), .A2(new_n407), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n246), .B1(new_n330), .B2(new_n340), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n342), .A2(new_n240), .A3(new_n344), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT34), .ZN(new_n419));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n419), .B1(new_n418), .B2(new_n420), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT69), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT69), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n421), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n416), .A2(G227gat), .A3(G233gat), .A4(new_n417), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429));
  XOR2_X1   g228(.A(G15gat), .B(G43gat), .Z(new_n430));
  XNOR2_X1  g229(.A(G71gat), .B(G99gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n428), .B(KEYINPUT32), .C1(new_n429), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(KEYINPUT32), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n428), .A2(new_n429), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n432), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n424), .A2(new_n427), .A3(new_n434), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n435), .A2(new_n436), .A3(new_n432), .ZN(new_n440));
  INV_X1    g239(.A(new_n434), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n426), .B(new_n439), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT36), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT83), .B1(new_n263), .B2(new_n258), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n263), .A2(KEYINPUT83), .A3(new_n258), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n269), .A2(new_n257), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n446), .A2(KEYINPUT39), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(KEYINPUT84), .B(KEYINPUT39), .Z(new_n450));
  INV_X1    g249(.A(new_n447), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n445), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n452), .A3(new_n277), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT40), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n453), .A2(KEYINPUT85), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT40), .A4(new_n277), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n456), .A2(new_n365), .A3(new_n366), .A4(new_n279), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT85), .B1(new_n453), .B2(new_n454), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n410), .A2(new_n412), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n346), .A2(new_n349), .A3(new_n299), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n354), .B1(new_n351), .B2(new_n356), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT37), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT38), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n361), .B1(new_n350), .B2(new_n357), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n361), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n463), .B(new_n464), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n363), .A2(new_n469), .B1(KEYINPUT37), .B2(new_n358), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n364), .B(new_n468), .C1(new_n470), .C2(new_n464), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n460), .B1(new_n471), .B2(new_n284), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n415), .B(new_n444), .C1(new_n459), .C2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n367), .B(new_n443), .C1(new_n403), .C2(new_n406), .ZN(new_n474));
  INV_X1    g273(.A(new_n284), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT35), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n410), .A2(new_n412), .B1(new_n442), .B2(new_n438), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n284), .A3(new_n367), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(KEYINPUT87), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n474), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n284), .A4(new_n478), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n473), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(G43gat), .A2(G50gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(G43gat), .A2(G50gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT90), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G43gat), .ZN(new_n490));
  INV_X1    g289(.A(G50gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G43gat), .A2(G50gat), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n492), .A2(KEYINPUT90), .A3(new_n488), .A4(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT14), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT15), .B1(new_n485), .B2(new_n486), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n508), .A2(new_n501), .A3(new_n499), .A4(new_n502), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n496), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT91), .B1(new_n503), .B2(new_n504), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n488), .A3(new_n493), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n494), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n512), .B1(new_n516), .B2(new_n509), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n511), .A2(KEYINPUT92), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n511), .A2(new_n517), .A3(KEYINPUT92), .A4(KEYINPUT17), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT16), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(G1gat), .B2(new_n523), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G8gat), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n526), .B(new_n529), .C1(G1gat), .C2(new_n523), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(KEYINPUT93), .Z(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n511), .A3(new_n517), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G169gat), .B(G197gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT12), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n535), .B(KEYINPUT13), .Z(new_n546));
  INV_X1    g345(.A(new_n536), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n531), .B1(new_n511), .B2(new_n517), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n531), .B1(new_n520), .B2(new_n521), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n535), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n545), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n539), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT94), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT89), .Z(new_n561));
  AND3_X1   g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n554), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n484), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  INV_X1    g367(.A(G78gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(G57gat), .A2(G64gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G57gat), .A2(G64gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n574), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n571), .A3(new_n572), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n576), .A3(new_n570), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(new_n237), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(KEYINPUT21), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n532), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n585), .B(G127gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n532), .A2(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n588), .A2(new_n591), .A3(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n511), .A2(new_n517), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT7), .ZN(new_n603));
  INV_X1    g402(.A(G85gat), .ZN(new_n604));
  INV_X1    g403(.A(G92gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT8), .ZN(new_n611));
  OR2_X1    g410(.A1(G85gat), .A2(G92gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n611), .B2(new_n612), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G99gat), .B(G106gat), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n611), .A2(new_n612), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT99), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n614), .ZN(new_n622));
  INV_X1    g421(.A(new_n618), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n609), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n601), .B1(new_n602), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n522), .B2(new_n625), .ZN(new_n627));
  XOR2_X1   g426(.A(G190gat), .B(G218gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT97), .ZN(new_n632));
  XOR2_X1   g431(.A(G134gat), .B(G162gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT101), .B1(new_n627), .B2(new_n629), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n627), .A2(KEYINPUT101), .A3(new_n629), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n634), .B(KEYINPUT98), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n627), .A2(new_n629), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n630), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n575), .A2(new_n577), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n576), .B1(new_n580), .B2(new_n570), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n623), .B1(new_n622), .B2(new_n609), .ZN(new_n649));
  AOI211_X1 g448(.A(new_n618), .B(new_n608), .C1(new_n621), .C2(new_n614), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n619), .A2(new_n582), .A3(new_n624), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n619), .A2(new_n582), .A3(new_n624), .A4(KEYINPUT10), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n645), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n653), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(new_n645), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT102), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n662), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n600), .A2(new_n643), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT103), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n566), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n475), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  INV_X1    g474(.A(new_n673), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n676), .A2(new_n367), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n367), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n529), .B1(new_n673), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT42), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(KEYINPUT42), .B2(new_n678), .ZN(G1325gat));
  OAI21_X1  g481(.A(G15gat), .B1(new_n676), .B2(new_n444), .ZN(new_n683));
  INV_X1    g482(.A(new_n443), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n676), .B2(new_n685), .ZN(G1326gat));
  NAND2_X1  g485(.A1(new_n407), .A2(new_n414), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(new_n600), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n666), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n565), .A2(new_n643), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n497), .A3(new_n475), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n484), .A2(new_n642), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n700));
  NAND3_X1  g499(.A1(new_n484), .A2(new_n642), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n564), .A2(KEYINPUT104), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n703), .B(new_n554), .C1(new_n562), .C2(new_n563), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n693), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n699), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n284), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n696), .A2(new_n708), .ZN(G1328gat));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n498), .A3(new_n679), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT46), .Z(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n707), .B2(new_n367), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1329gat));
  NAND3_X1  g512(.A1(new_n694), .A2(new_n490), .A3(new_n443), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT106), .ZN(new_n715));
  OAI21_X1  g514(.A(G43gat), .B1(new_n707), .B2(new_n444), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n714), .A2(KEYINPUT47), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n718), .A2(new_n719), .A3(new_n716), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n718), .B2(new_n716), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n717), .A2(KEYINPUT47), .B1(new_n720), .B2(new_n721), .ZN(G1330gat));
  NAND3_X1  g521(.A1(new_n694), .A2(new_n491), .A3(new_n688), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT109), .B1(new_n707), .B2(new_n460), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G50gat), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n707), .A2(KEYINPUT109), .A3(new_n460), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT48), .B(new_n723), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G50gat), .B1(new_n707), .B2(new_n687), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n723), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(G1331gat));
  NOR3_X1   g530(.A1(new_n692), .A2(new_n642), .A3(new_n666), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n484), .A2(new_n705), .A3(new_n732), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT110), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(KEYINPUT110), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n475), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g538(.A1(new_n736), .A2(new_n367), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n736), .B2(new_n444), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n443), .A2(new_n568), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n736), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1334gat));
  NOR2_X1   g548(.A1(new_n736), .A2(new_n687), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n569), .ZN(G1335gat));
  NAND4_X1  g550(.A1(new_n484), .A2(new_n692), .A3(new_n642), .A4(new_n705), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT51), .Z(new_n753));
  NAND4_X1  g552(.A1(new_n753), .A2(new_n604), .A3(new_n475), .A4(new_n665), .ZN(new_n754));
  INV_X1    g553(.A(new_n705), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n755), .A2(new_n600), .A3(new_n666), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n699), .A2(new_n701), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n699), .A2(KEYINPUT112), .A3(new_n701), .A4(new_n756), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(new_n475), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n754), .B1(new_n761), .B2(new_n604), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT113), .ZN(G1336gat));
  NOR3_X1   g562(.A1(new_n367), .A2(G92gat), .A3(new_n666), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n753), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI21_X1  g565(.A(G92gat), .B1(new_n757), .B2(new_n367), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n759), .A2(new_n679), .A3(new_n760), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n752), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n752), .B2(KEYINPUT114), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n769), .A2(G92gat), .B1(new_n772), .B2(new_n764), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n768), .B1(new_n773), .B2(new_n766), .ZN(G1337gat));
  INV_X1    g573(.A(new_n444), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n775), .A3(new_n760), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G99gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n684), .A2(G99gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n753), .A2(new_n665), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1338gat));
  NOR3_X1   g579(.A1(new_n460), .A2(G106gat), .A3(new_n666), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n753), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  OAI21_X1  g582(.A(G106gat), .B1(new_n757), .B2(new_n460), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n759), .A2(new_n688), .A3(new_n760), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(new_n781), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n770), .A2(new_n771), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT115), .B1(new_n791), .B2(KEYINPUT53), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n789), .B1(new_n786), .B2(G106gat), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n793), .A2(new_n794), .A3(new_n783), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n785), .B1(new_n792), .B2(new_n795), .ZN(G1339gat));
  NAND2_X1  g595(.A1(new_n654), .A2(new_n655), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n644), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n654), .A2(new_n655), .A3(new_n645), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n662), .B1(new_n656), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n664), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n802), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n702), .A2(new_n704), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n550), .A2(new_n547), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n547), .A2(new_n548), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n809), .A2(new_n535), .B1(new_n810), .B2(new_n546), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n544), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n665), .A2(new_n554), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n642), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n807), .A2(new_n642), .A3(new_n554), .A4(new_n812), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n692), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n705), .A2(new_n668), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n688), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n475), .A2(new_n367), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n684), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n227), .B1(new_n822), .B2(new_n564), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n284), .B1(new_n817), .B2(new_n818), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n481), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(new_n228), .A3(new_n705), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n823), .A2(new_n826), .ZN(G1340gat));
  AOI21_X1  g626(.A(new_n229), .B1(new_n822), .B2(new_n665), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n825), .A2(new_n226), .A3(new_n666), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT116), .ZN(G1341gat));
  NAND3_X1  g630(.A1(new_n822), .A2(G127gat), .A3(new_n600), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  INV_X1    g634(.A(new_n825), .ZN(new_n836));
  AOI21_X1  g635(.A(G127gat), .B1(new_n836), .B2(new_n600), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(G1342gat));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n238), .A3(new_n642), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n840));
  INV_X1    g639(.A(new_n822), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n841), .B2(new_n643), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n775), .A2(new_n820), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n687), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n803), .A2(new_n664), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n806), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g651(.A(KEYINPUT119), .B(new_n850), .C1(new_n800), .C2(new_n802), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n848), .B(KEYINPUT120), .C1(new_n852), .C2(new_n853), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n564), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n642), .B1(new_n858), .B2(new_n813), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n692), .B1(new_n859), .B2(new_n816), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT121), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n818), .B1(new_n860), .B2(KEYINPUT121), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT122), .B(new_n847), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n460), .B1(new_n817), .B2(new_n818), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(KEYINPUT57), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n861), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT122), .B1(new_n868), .B2(new_n847), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n845), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n564), .ZN(new_n871));
  OAI21_X1  g670(.A(G141gat), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n775), .A2(new_n460), .A3(new_n679), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n824), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n206), .A3(new_n564), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n872), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n870), .B2(new_n705), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n877), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n880), .B2(new_n873), .ZN(G1344gat));
  NOR3_X1   g680(.A1(new_n775), .A2(new_n666), .A3(new_n820), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883));
  INV_X1    g682(.A(new_n460), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n808), .A2(new_n813), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n643), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n600), .B1(new_n886), .B2(new_n815), .ZN(new_n887));
  INV_X1    g686(.A(new_n818), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT57), .B(new_n884), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n858), .A2(new_n813), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n643), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n600), .B1(new_n891), .B2(new_n815), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n669), .A2(new_n871), .A3(new_n671), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n688), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n846), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n883), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT123), .B1(new_n865), .B2(KEYINPUT57), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n882), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G148gat), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n665), .B(new_n845), .C1(new_n866), .C2(new_n869), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n210), .A2(KEYINPUT59), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n899), .A2(KEYINPUT59), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n875), .A2(G148gat), .A3(new_n666), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT124), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  INV_X1    g704(.A(new_n903), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n900), .A2(new_n901), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n898), .B2(G148gat), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n905), .B(new_n906), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n904), .A2(new_n910), .ZN(G1345gat));
  INV_X1    g710(.A(new_n215), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(new_n870), .B2(new_n692), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n876), .A2(new_n215), .A3(new_n600), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  OR3_X1    g714(.A1(new_n870), .A2(new_n216), .A3(new_n643), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n216), .B1(new_n875), .B2(new_n643), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(G1347gat));
  AOI21_X1  g717(.A(new_n475), .B1(new_n817), .B2(new_n818), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n477), .A2(new_n679), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT125), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n755), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n679), .A2(new_n284), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n684), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n819), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n564), .A2(G169gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1348gat));
  INV_X1    g727(.A(new_n926), .ZN(new_n929));
  OAI21_X1  g728(.A(G176gat), .B1(new_n929), .B2(new_n666), .ZN(new_n930));
  INV_X1    g729(.A(G176gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n922), .A2(new_n931), .A3(new_n665), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1349gat));
  NAND2_X1  g732(.A1(new_n926), .A2(new_n600), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n600), .A2(new_n305), .ZN(new_n935));
  AOI22_X1  g734(.A1(new_n934), .A2(G183gat), .B1(new_n922), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g736(.A(new_n306), .B1(new_n926), .B2(new_n642), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT61), .Z(new_n939));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n306), .A3(new_n642), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n775), .A2(new_n924), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n564), .B(new_n942), .C1(new_n896), .C2(new_n897), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G197gat), .ZN(new_n944));
  AND4_X1   g743(.A1(new_n884), .A2(new_n919), .A3(new_n679), .A4(new_n444), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n288), .A3(new_n755), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n947), .B(new_n948), .ZN(G1352gat));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n289), .A3(new_n665), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  OR2_X1    g750(.A1(new_n896), .A2(new_n897), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n665), .A3(new_n942), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G204gat), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n953), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(G1353gat));
  INV_X1    g757(.A(G211gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n945), .A2(new_n959), .A3(new_n600), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n952), .A2(new_n600), .A3(new_n942), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  INV_X1    g763(.A(G218gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n945), .A2(new_n965), .A3(new_n642), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n952), .A2(new_n642), .A3(new_n942), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n965), .ZN(G1355gat));
endmodule


