//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n461), .A3(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n458), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(new_n461), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n469), .B1(new_n460), .B2(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n467), .A2(G137), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n472));
  AND3_X1   g047(.A1(new_n465), .A2(new_n471), .A3(new_n472), .ZN(G160));
  AND4_X1   g048(.A1(G2105), .A2(new_n470), .A3(new_n466), .A4(new_n461), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(G112), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n470), .A2(new_n466), .A3(new_n468), .A4(new_n461), .ZN(new_n478));
  OR2_X1    g053(.A1(new_n478), .A2(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI221_X1 g057(.A(new_n475), .B1(new_n476), .B2(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(new_n474), .A2(G126), .ZN(new_n485));
  OR2_X1    g060(.A1(KEYINPUT70), .A2(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT70), .A2(G114), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n468), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n470), .A2(new_n466), .A3(new_n492), .A4(new_n461), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n459), .A2(new_n461), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n491), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n485), .B(new_n490), .C1(new_n494), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n500), .B1(new_n506), .B2(G651), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n503), .A2(new_n502), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n509), .A2(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n506), .A2(new_n500), .A3(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n521), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  OR2_X1    g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(new_n508), .A3(G89), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT72), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n538), .B(new_n535), .C1(new_n502), .C2(new_n503), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n524), .A2(new_n534), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  OAI211_X1 g117(.A(G52), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n513), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  OAI21_X1  g121(.A(G64), .B1(new_n502), .B2(new_n503), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n509), .A2(new_n551), .B1(new_n513), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n532), .A2(G56), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n546), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT74), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n509), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n528), .A2(new_n566), .A3(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n504), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n530), .A2(new_n531), .B1(new_n526), .B2(new_n527), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n571), .A2(G651), .B1(new_n572), .B2(G91), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n568), .A2(new_n573), .ZN(G299));
  NAND3_X1  g149(.A1(new_n532), .A2(new_n508), .A3(G90), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n543), .B(new_n575), .C1(new_n576), .C2(new_n546), .ZN(G301));
  NAND2_X1  g152(.A1(new_n516), .A2(new_n517), .ZN(G303));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n504), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n528), .B2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n572), .A2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  OAI211_X1 g158(.A(G48), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n572), .A2(G86), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n504), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(G305));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n530), .B2(new_n531), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT76), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n597), .B(new_n594), .C1(new_n504), .C2(new_n592), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(G651), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n572), .A2(G85), .B1(new_n528), .B2(G47), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n600), .B1(new_n599), .B2(new_n601), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n530), .B2(new_n531), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT78), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n613), .B(new_n610), .C1(new_n504), .C2(new_n608), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n612), .A2(G651), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n513), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n532), .A2(new_n508), .A3(KEYINPUT10), .A4(G92), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n528), .A2(G54), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n615), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n607), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n607), .B1(new_n623), .B2(G868), .ZN(G321));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(G299), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G168), .B2(new_n626), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(G168), .B2(new_n626), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n623), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND4_X1  g210(.A1(new_n470), .A2(new_n466), .A3(G2105), .A4(new_n461), .ZN(new_n636));
  INV_X1    g211(.A(G123), .ZN(new_n637));
  OAI21_X1  g212(.A(KEYINPUT79), .B1(new_n468), .B2(G111), .ZN(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(G2104), .A3(new_n639), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n468), .A2(KEYINPUT79), .A3(G111), .ZN(new_n641));
  OAI22_X1  g216(.A1(new_n636), .A2(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n481), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(G135), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(G156));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n656), .B(new_n662), .Z(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  INV_X1    g253(.A(new_n669), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n672), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2096), .B(G2100), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n692), .A2(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(KEYINPUT20), .ZN(new_n694));
  OAI221_X1 g269(.A(new_n689), .B1(new_n686), .B2(new_n690), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT87), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n703), .A2(G6), .ZN(new_n709));
  INV_X1    g284(.A(G305), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n703), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT84), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n528), .A2(G49), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n532), .A2(new_n508), .A3(G87), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT85), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n581), .A2(new_n720), .A3(new_n582), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G23), .B(new_n722), .S(G16), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT33), .B(G1976), .Z(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT86), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n708), .A2(new_n714), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n643), .A2(G131), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n734));
  INV_X1    g309(.A(G107), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n474), .B2(G119), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n731), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT35), .B(G1991), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT83), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n703), .A2(G24), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n605), .B2(new_n703), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G1986), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n745), .A2(G1986), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n743), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n729), .A2(new_n730), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT36), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G35), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G162), .B2(G29), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT29), .B(G2090), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n703), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n623), .B2(new_n703), .ZN(new_n756));
  INV_X1    g331(.A(G1348), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n703), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G299), .B2(G16), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT24), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n731), .B1(new_n765), .B2(G34), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n765), .B2(G34), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G160), .B2(G29), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n764), .A2(G1956), .B1(G2084), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n703), .A2(G19), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT88), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n557), .B2(new_n703), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1341), .ZN(new_n773));
  INV_X1    g348(.A(G1956), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n763), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n754), .A2(new_n758), .A3(new_n769), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n731), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT28), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n643), .A2(G140), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n780));
  OR3_X1    g355(.A1(KEYINPUT89), .A2(G104), .A3(G2105), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT89), .B1(G104), .B2(G2105), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n474), .B2(G128), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(new_n731), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n703), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G171), .B2(new_n703), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n768), .A2(G2084), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n731), .A2(G27), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n731), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n791), .B(new_n792), .C1(G2078), .C2(new_n794), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n788), .B(new_n795), .C1(G2078), .C2(new_n794), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT31), .B(G11), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT94), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n645), .A2(new_n731), .ZN(new_n799));
  INV_X1    g374(.A(G28), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT30), .ZN(new_n801));
  AOI21_X1  g376(.A(G29), .B1(new_n800), .B2(KEYINPUT30), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n798), .B(new_n799), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n703), .A2(G21), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G168), .B2(new_n703), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G1966), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT93), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n790), .A2(G1961), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT95), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n805), .A2(G1966), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n803), .A2(new_n807), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n776), .B(new_n796), .C1(KEYINPUT96), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n731), .A2(G33), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT25), .Z(new_n815));
  INV_X1    g390(.A(G139), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n481), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT90), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(new_n468), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n813), .B1(new_n822), .B2(new_n731), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G2072), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n812), .B(new_n824), .C1(KEYINPUT96), .C2(new_n811), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(G2072), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT91), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n731), .A2(G32), .ZN(new_n828));
  NAND3_X1  g403(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT26), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G129), .B2(new_n474), .ZN(new_n834));
  INV_X1    g409(.A(G141), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n481), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n828), .B1(new_n838), .B2(new_n731), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT27), .ZN(new_n840));
  INV_X1    g415(.A(G1996), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n825), .A2(new_n827), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n750), .A2(new_n843), .ZN(G150));
  INV_X1    g419(.A(G150), .ZN(G311));
  NAND2_X1  g420(.A1(new_n623), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n509), .A2(new_n848), .B1(new_n513), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(G67), .B1(new_n502), .B2(new_n503), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n546), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI22_X1  g428(.A1(new_n556), .A2(new_n553), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n554), .A2(new_n555), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G651), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n572), .A2(G81), .B1(new_n528), .B2(G43), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n572), .A2(G93), .B1(new_n528), .B2(G55), .ZN(new_n858));
  INV_X1    g433(.A(new_n853), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n847), .B(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT98), .B(G860), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n866), .B1(new_n858), .B2(new_n859), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  XNOR2_X1  g445(.A(new_n836), .B(KEYINPUT92), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n498), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n838), .A2(G164), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n821), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n821), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n785), .ZN(new_n877));
  INV_X1    g452(.A(new_n785), .ZN(new_n878));
  INV_X1    g453(.A(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n874), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n474), .A2(G130), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n468), .A2(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n643), .B2(G142), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(new_n649), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n738), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n877), .A2(new_n880), .A3(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(KEYINPUT100), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(KEYINPUT100), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n877), .A2(new_n880), .ZN(new_n891));
  INV_X1    g466(.A(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(G160), .B(KEYINPUT99), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G162), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n645), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n889), .A2(new_n890), .A3(new_n893), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n888), .ZN(new_n898));
  INV_X1    g473(.A(new_n896), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g477(.A(new_n626), .B1(new_n850), .B2(new_n853), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n632), .B(new_n861), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n622), .A2(G299), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n618), .A2(new_n619), .B1(G54), .B2(new_n528), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n906), .A2(new_n615), .B1(new_n568), .B2(new_n573), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT41), .B1(new_n905), .B2(new_n907), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n622), .A2(G299), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n906), .A2(new_n568), .A3(new_n573), .A4(new_n615), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n905), .A2(new_n907), .A3(KEYINPUT41), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT101), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n909), .B1(new_n919), .B2(new_n904), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n710), .A2(new_n722), .ZN(new_n921));
  NAND3_X1  g496(.A1(G305), .A2(new_n719), .A3(new_n721), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n599), .A2(new_n601), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT77), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n925), .A2(G303), .A3(new_n602), .ZN(new_n926));
  AOI21_X1  g501(.A(G303), .B1(new_n925), .B2(new_n602), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(G166), .B1(new_n603), .B2(new_n604), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n925), .A2(G303), .A3(new_n602), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n929), .A2(new_n930), .A3(new_n922), .A4(new_n921), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n920), .B(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n903), .B1(new_n935), .B2(new_n626), .ZN(G295));
  OAI21_X1  g511(.A(new_n903), .B1(new_n935), .B2(new_n626), .ZN(G331));
  NAND4_X1  g512(.A1(G171), .A2(new_n524), .A3(new_n534), .A4(new_n540), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n538), .B1(new_n532), .B2(new_n535), .ZN(new_n939));
  INV_X1    g514(.A(new_n539), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n533), .B(new_n529), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT7), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n520), .B2(new_n522), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(G301), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n861), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n861), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n908), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(KEYINPUT104), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n946), .A2(new_n938), .B1(new_n854), .B2(new_n860), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n948), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n932), .B(new_n951), .C1(new_n919), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT105), .ZN(new_n958));
  INV_X1    g533(.A(G37), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n947), .A2(new_n954), .A3(new_n861), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n954), .B1(new_n947), .B2(new_n861), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n949), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n918), .A3(new_n916), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n932), .A4(new_n951), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n958), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n967));
  INV_X1    g542(.A(new_n932), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n917), .A2(new_n969), .B1(new_n948), .B2(new_n953), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT106), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n949), .B(new_n908), .C1(new_n960), .C2(new_n961), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n970), .A2(KEYINPUT106), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n966), .A2(new_n967), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n963), .A2(new_n951), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n968), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n966), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n979), .B2(new_n967), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  AOI21_X1  g558(.A(G37), .B1(new_n957), .B2(KEYINPUT105), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(new_n965), .A3(new_n975), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n985), .B2(KEYINPUT43), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n984), .A2(new_n967), .A3(new_n978), .A4(new_n965), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n983), .B(new_n986), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n966), .A2(KEYINPUT107), .A3(new_n967), .A4(new_n978), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n987), .A2(new_n988), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n983), .B1(new_n995), .B2(new_n986), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n982), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT109), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(new_n982), .C1(new_n992), .C2(new_n996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(G397));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n493), .A2(KEYINPUT4), .B1(new_n495), .B2(new_n496), .ZN(new_n1003));
  INV_X1    g578(.A(G126), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n636), .A2(new_n1004), .B1(new_n488), .B2(new_n489), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n465), .A2(new_n471), .A3(G40), .A4(new_n472), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n785), .B(new_n787), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n871), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n841), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT46), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n871), .A2(G1996), .A3(new_n1010), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT110), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n871), .A2(G1996), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1010), .B1(new_n1011), .B2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n738), .A2(new_n742), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n738), .A2(new_n742), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1010), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G290), .A2(G1986), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n1010), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT48), .Z(new_n1029));
  OAI21_X1  g604(.A(new_n1017), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(G2067), .B2(new_n878), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1030), .B1(new_n1010), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT124), .ZN(new_n1034));
  AND2_X1   g609(.A1(G290), .A2(G1986), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1010), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1022), .A2(new_n1036), .A3(new_n1025), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n719), .A2(G1976), .A3(new_n721), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1038), .A2(KEYINPUT112), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1976), .B1(new_n581), .B2(new_n582), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1039), .B(new_n1041), .C1(KEYINPUT52), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1042), .B(G8), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(KEYINPUT112), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(new_n1045), .C1(new_n1046), .C2(new_n1040), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n590), .A2(new_n586), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT75), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n584), .B(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT49), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n590), .B2(KEYINPUT113), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n585), .A2(new_n1054), .A3(new_n586), .A4(new_n590), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1053), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1043), .A2(new_n1047), .B1(new_n1041), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G303), .A2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(new_n1002), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT111), .ZN(new_n1067));
  INV_X1    g642(.A(G2090), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1009), .B1(new_n1006), .B2(KEYINPUT50), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1065), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  AND4_X1   g647(.A1(G40), .A2(new_n465), .A3(new_n471), .A4(new_n472), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1007), .A2(G1384), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1008), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n707), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1063), .A2(new_n1078), .A3(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1058), .A2(new_n1041), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G288), .A2(G1976), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1080), .A2(new_n1081), .B1(new_n1052), .B2(new_n710), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1060), .A2(new_n1079), .B1(new_n1082), .B2(new_n1040), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1059), .A2(new_n1079), .ZN(new_n1084));
  INV_X1    g659(.A(G1966), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT45), .B1(new_n498), .B2(new_n1002), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT116), .ZN(new_n1089));
  INV_X1    g664(.A(G2084), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1067), .A2(new_n1090), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1076), .A2(new_n1092), .A3(new_n1085), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1094), .A2(G8), .A3(G168), .ZN(new_n1095));
  INV_X1    g670(.A(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1069), .A2(KEYINPUT114), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1065), .B1(new_n1069), .B2(KEYINPUT114), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1006), .A2(KEYINPUT50), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1073), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n1097), .A4(new_n1065), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n1068), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1096), .B1(new_n1107), .B2(new_n1077), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1084), .B(new_n1095), .C1(new_n1108), .C2(new_n1063), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1078), .A2(G8), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1063), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1084), .A2(new_n1095), .A3(KEYINPUT63), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1083), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n774), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1117));
  XOR2_X1   g692(.A(G299), .B(KEYINPUT57), .Z(new_n1118));
  NOR2_X1   g693(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1118), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1124), .A2(new_n757), .B1(new_n787), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(new_n622), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1122), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT117), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1130), .B(new_n1122), .C1(new_n1123), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1118), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1066), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1956), .B1(new_n1134), .B2(new_n1097), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1121), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n1122), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT61), .B1(new_n1123), .B2(KEYINPUT119), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n623), .B2(KEYINPUT120), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n623), .A2(KEYINPUT120), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1126), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT118), .B(new_n1146), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1149), .B(new_n1150), .C1(new_n1076), .C2(G1996), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n557), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(KEYINPUT59), .A3(new_n557), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1145), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1137), .A2(KEYINPUT61), .A3(new_n1122), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1144), .B1(new_n1126), .B2(new_n1143), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(KEYINPUT60), .B2(new_n1126), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1132), .B1(new_n1141), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(G1961), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1124), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT53), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1076), .B2(G2078), .ZN(new_n1165));
  INV_X1    g740(.A(G2078), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1119), .A2(KEYINPUT53), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1163), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(G171), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1008), .A2(new_n1073), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1075), .A2(KEYINPUT53), .A3(new_n1166), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1177), .A2(G301), .A3(new_n1165), .A4(new_n1163), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1171), .A2(new_n1172), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1059), .A2(new_n1079), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1107), .A2(new_n1077), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(G8), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1182), .B1(new_n1184), .B2(new_n1113), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1177), .A2(new_n1165), .A3(new_n1163), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(G171), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1187), .B(KEYINPUT54), .C1(G171), .C2(new_n1168), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1009), .B1(new_n498), .B2(new_n1074), .ZN(new_n1189));
  AOI211_X1 g764(.A(KEYINPUT116), .B(G1966), .C1(new_n1189), .C2(new_n1008), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1092), .B1(new_n1076), .B2(new_n1085), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(G168), .B1(new_n1192), .B2(new_n1091), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1089), .A2(G168), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(G8), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT51), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1194), .A2(G8), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT51), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1181), .A2(new_n1185), .A3(new_n1188), .A4(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1116), .B1(new_n1161), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1196), .A2(new_n1199), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1204), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1084), .B1(new_n1108), .B2(new_n1063), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1172), .ZN(new_n1210));
  AOI21_X1  g785(.A(KEYINPUT121), .B1(new_n1168), .B2(G171), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1207), .A2(new_n1208), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1094), .A2(G286), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1198), .B1(new_n1197), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1195), .A2(KEYINPUT51), .ZN(new_n1217));
  OAI21_X1  g792(.A(KEYINPUT62), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1196), .A2(new_n1199), .A3(new_n1204), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1213), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1220), .A2(KEYINPUT123), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1214), .A2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g797(.A(new_n1034), .B(new_n1037), .C1(new_n1203), .C2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g798(.A1(new_n1141), .A2(new_n1157), .A3(new_n1159), .A4(new_n1156), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1224), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1225));
  AND3_X1   g800(.A1(new_n1188), .A2(new_n1185), .A3(new_n1200), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1225), .A2(new_n1226), .A3(new_n1181), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1208), .B1(new_n1207), .B2(new_n1213), .ZN(new_n1228));
  AND4_X1   g803(.A1(new_n1208), .A2(new_n1213), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1229));
  OAI211_X1 g804(.A(new_n1227), .B(new_n1116), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1037), .ZN(new_n1231));
  AOI21_X1  g806(.A(KEYINPUT124), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1033), .B1(new_n1223), .B2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g808(.A(G319), .ZN(new_n1235));
  NOR2_X1   g809(.A1(G227), .A2(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g810(.A(new_n1236), .B(KEYINPUT126), .ZN(new_n1237));
  OAI211_X1 g811(.A(new_n1237), .B(new_n701), .C1(new_n667), .C2(new_n666), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n897), .B2(new_n900), .ZN(new_n1239));
  AND3_X1   g813(.A1(new_n1239), .A2(KEYINPUT127), .A3(new_n980), .ZN(new_n1240));
  AOI21_X1  g814(.A(KEYINPUT127), .B1(new_n1239), .B2(new_n980), .ZN(new_n1241));
  NOR2_X1   g815(.A1(new_n1240), .A2(new_n1241), .ZN(G308));
  NAND2_X1  g816(.A1(new_n1239), .A2(new_n980), .ZN(G225));
endmodule


