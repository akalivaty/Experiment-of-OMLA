//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT76), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT11), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G134), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT65), .B1(new_n200), .B2(G134), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n197), .A3(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n202), .A2(G131), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n203), .A2(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n198), .A2(new_n201), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G104), .B(G107), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT78), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G107), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G104), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n216), .B(G101), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n220), .A2(G101), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT77), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(new_n219), .A3(KEYINPUT3), .A4(G104), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT64), .A2(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT64), .A2(G143), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(G146), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G146), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT64), .A2(G143), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT64), .A2(G143), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n239), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT1), .B1(new_n233), .B2(G146), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n242), .A2(new_n244), .B1(G128), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n229), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n224), .A2(new_n219), .A3(G104), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n226), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n215), .A2(new_n221), .B1(new_n252), .B2(new_n223), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n236), .B1(new_n242), .B2(KEYINPUT1), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n240), .A2(new_n241), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n234), .B1(new_n256), .B2(G146), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n212), .B1(new_n248), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT80), .A2(KEYINPUT12), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT10), .ZN(new_n267));
  AND2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n232), .A2(new_n235), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n230), .A2(new_n231), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n243), .B1(new_n270), .B2(new_n239), .ZN(new_n271));
  NOR2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n269), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G101), .ZN(new_n277));
  INV_X1    g091(.A(new_n220), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n252), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n220), .B1(new_n251), .B2(new_n226), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n228), .B(KEYINPUT4), .C1(new_n281), .C2(new_n214), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n267), .A2(new_n259), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT10), .B1(new_n238), .B2(new_n246), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n229), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n245), .A2(G128), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n254), .B1(new_n271), .B2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n253), .A2(new_n288), .A3(KEYINPUT79), .A4(KEYINPUT10), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n283), .A2(new_n290), .A3(new_n212), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n196), .B1(new_n266), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n212), .B1(new_n283), .B2(new_n290), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n283), .A2(new_n290), .A3(new_n212), .ZN(new_n295));
  INV_X1    g109(.A(new_n196), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT81), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n292), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(G469), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n265), .A2(new_n295), .A3(new_n296), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n196), .B1(new_n291), .B2(new_n293), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(G469), .A2(G902), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n191), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G475), .ZN(new_n311));
  INV_X1    g125(.A(G237), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n312), .A2(new_n192), .A3(G214), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G143), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n314), .B(new_n208), .C1(new_n270), .C2(new_n313), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT18), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n314), .B(new_n316), .C1(new_n270), .C2(new_n313), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT88), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT88), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G125), .B(G140), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n323), .A2(new_n239), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n239), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n314), .B1(new_n270), .B2(new_n313), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G131), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n328), .B2(new_n316), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n323), .A2(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n333), .A2(KEYINPUT16), .A3(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n239), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(G146), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n327), .A2(KEYINPUT17), .A3(G131), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n328), .A2(new_n315), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n339), .B(new_n340), .C1(KEYINPUT17), .C2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G113), .B(G122), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(new_n217), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT90), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n331), .A2(new_n342), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n344), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n311), .B1(new_n348), .B2(new_n190), .ZN(new_n349));
  INV_X1    g163(.A(new_n346), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n337), .A2(KEYINPUT74), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(KEYINPUT74), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n323), .B(KEYINPUT19), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n239), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n341), .A2(new_n351), .A3(new_n352), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n331), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n344), .B1(new_n356), .B2(KEYINPUT89), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT89), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n331), .A2(new_n358), .A3(new_n355), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n350), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(G475), .A2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT20), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n329), .B1(new_n321), .B2(new_n320), .ZN(new_n364));
  INV_X1    g178(.A(new_n355), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT89), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n344), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n359), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n346), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT20), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n361), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n349), .B1(new_n363), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT92), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n256), .A2(G128), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n236), .A2(G143), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n197), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n197), .B1(new_n374), .B2(new_n375), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT91), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n376), .ZN(new_n382));
  INV_X1    g196(.A(G116), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n383), .A2(G122), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n219), .B1(new_n384), .B2(KEYINPUT14), .ZN(new_n385));
  XNOR2_X1  g199(.A(G116), .B(G122), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n379), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n386), .B(new_n219), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n374), .A2(KEYINPUT13), .A3(new_n375), .ZN(new_n390));
  OAI21_X1  g204(.A(G134), .B1(new_n374), .B2(KEYINPUT13), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n376), .B(new_n389), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G217), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n188), .A2(new_n394), .A3(G953), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n388), .A2(new_n392), .A3(new_n395), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT15), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G478), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n190), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(G902), .B1(new_n397), .B2(new_n398), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(new_n401), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n373), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n404), .A2(new_n401), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT92), .A3(new_n402), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n192), .A2(G952), .ZN(new_n410));
  INV_X1    g224(.A(G234), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(new_n312), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n190), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n372), .A2(new_n409), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n310), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G214), .B1(G237), .B2(G902), .ZN(new_n420));
  OAI21_X1  g234(.A(G210), .B1(G237), .B2(G902), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n383), .A2(G119), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT66), .ZN(new_n423));
  INV_X1    g237(.A(G119), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(G116), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n383), .A2(KEYINPUT66), .A3(G119), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT5), .ZN(new_n428));
  INV_X1    g242(.A(G113), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT5), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n429), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT2), .B(G113), .Z(new_n432));
  AOI22_X1  g246(.A1(new_n428), .A2(new_n431), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n253), .ZN(new_n434));
  XNOR2_X1  g248(.A(G110), .B(G122), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n228), .A2(KEYINPUT4), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n281), .A2(new_n214), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n427), .A2(new_n432), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n427), .A2(new_n432), .ZN(new_n440));
  OAI22_X1  g254(.A1(new_n439), .A2(new_n440), .B1(new_n281), .B2(new_n277), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n434), .B(new_n435), .C1(new_n438), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT6), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n427), .B(new_n432), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n282), .B(new_n444), .C1(new_n281), .C2(new_n277), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n435), .B1(new_n445), .B2(new_n434), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT82), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n434), .B1(new_n438), .B2(new_n441), .ZN(new_n448));
  INV_X1    g262(.A(new_n435), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT6), .A4(new_n442), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n275), .A2(G125), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n247), .A2(new_n333), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n275), .A2(new_n457), .A3(G125), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G224), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n455), .A2(new_n456), .A3(new_n463), .A4(new_n458), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n450), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n453), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT85), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n447), .B2(new_n452), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n465), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n463), .A2(KEYINPUT7), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n459), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n459), .B2(new_n476), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n433), .B(new_n229), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n435), .B(KEYINPUT8), .Z(new_n482));
  INV_X1    g296(.A(KEYINPUT7), .ZN(new_n483));
  OAI221_X1 g297(.A(new_n442), .B1(new_n481), .B2(new_n482), .C1(new_n464), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n190), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n421), .B1(new_n474), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n421), .ZN(new_n488));
  AOI211_X1 g302(.A(new_n488), .B(new_n485), .C1(new_n470), .C2(new_n473), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n420), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n420), .ZN(new_n493));
  AND4_X1   g307(.A1(new_n472), .A2(new_n453), .A3(new_n465), .A4(new_n468), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n472), .B1(new_n471), .B2(new_n465), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n486), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n488), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n474), .A2(new_n421), .A3(new_n486), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n236), .A2(G119), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n236), .A2(G119), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT24), .B(G110), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n504), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g324(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n511), .A2(new_n509), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n512), .B2(new_n501), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n508), .B1(new_n513), .B2(G110), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n352), .A3(new_n351), .A4(new_n325), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(G110), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n338), .B(new_n516), .C1(new_n507), .C2(new_n506), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n187), .A2(new_n411), .A3(G953), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n519), .B(new_n520), .Z(new_n521));
  XNOR2_X1  g335(.A(new_n518), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n190), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n523), .A2(KEYINPUT25), .ZN(new_n524));
  OAI21_X1  g338(.A(G217), .B1(new_n411), .B2(G902), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n523), .B2(KEYINPUT25), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(G902), .B1(new_n411), .B2(G217), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n242), .A2(new_n244), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n273), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n534), .B(new_n269), .C1(new_n207), .C2(new_n211), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n200), .A2(G134), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n197), .A2(G137), .ZN(new_n538));
  OAI21_X1  g352(.A(G131), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n209), .A2(new_n208), .A3(new_n210), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n539), .B(new_n540), .C1(new_n238), .C2(new_n246), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n536), .B1(new_n535), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n444), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n439), .A2(new_n440), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n541), .B(new_n545), .C1(new_n212), .C2(new_n275), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n312), .A2(new_n192), .A3(G210), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(G101), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT68), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(KEYINPUT68), .A3(new_n551), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n544), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n544), .A2(new_n554), .A3(KEYINPUT31), .A4(new_n555), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n546), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n545), .B1(new_n535), .B2(new_n541), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT28), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n535), .A2(new_n564), .A3(new_n541), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n535), .B2(new_n541), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n566), .A2(new_n567), .A3(new_n444), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n563), .B1(new_n568), .B2(KEYINPUT28), .ZN(new_n569));
  INV_X1    g383(.A(new_n551), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n560), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(G472), .A2(G902), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n558), .A2(new_n559), .B1(new_n569), .B2(new_n570), .ZN(new_n576));
  INV_X1    g390(.A(new_n573), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT29), .ZN(new_n580));
  INV_X1    g394(.A(new_n543), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n561), .B1(new_n583), .B2(new_n444), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n580), .B1(new_n584), .B2(new_n551), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n567), .A2(new_n444), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT28), .B1(new_n586), .B2(new_n565), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT28), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n535), .A2(new_n541), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n444), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n590), .B2(new_n546), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n587), .A2(new_n591), .A3(new_n570), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n190), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n551), .A2(KEYINPUT29), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT71), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n562), .A2(KEYINPUT71), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT70), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n546), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n546), .A2(new_n598), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n596), .B(new_n597), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n594), .B(new_n587), .C1(new_n601), .C2(KEYINPUT28), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n593), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n532), .B1(new_n579), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n419), .A2(new_n492), .A3(new_n500), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  INV_X1    g420(.A(new_n310), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n572), .A2(new_n573), .ZN(new_n608));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n560), .B2(new_n571), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n607), .A2(new_n532), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n190), .A2(G478), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n399), .A2(KEYINPUT33), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n397), .A2(new_n615), .A3(new_n398), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT93), .B1(new_n404), .B2(G478), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n619), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n372), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n499), .A2(new_n417), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n612), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT94), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  OAI211_X1 g442(.A(new_n420), .B(new_n417), .C1(new_n487), .C2(new_n489), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n370), .B1(new_n369), .B2(new_n361), .ZN(new_n630));
  AOI211_X1 g444(.A(KEYINPUT20), .B(new_n362), .C1(new_n368), .C2(new_n346), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n348), .A2(new_n190), .ZN(new_n632));
  OAI22_X1  g446(.A1(new_n630), .A2(new_n631), .B1(new_n311), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n409), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT95), .B1(new_n629), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n499), .A2(new_n637), .A3(new_n417), .A4(new_n634), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n612), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT97), .B(G107), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n521), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n518), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n528), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n611), .B1(new_n527), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n419), .A2(new_n492), .A3(new_n500), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n650), .B(new_n652), .ZN(G12));
  NAND2_X1  g467(.A1(new_n499), .A2(new_n310), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT99), .B(G900), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n414), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n412), .B1(new_n656), .B2(KEYINPUT100), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(KEYINPUT100), .B2(new_n656), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT101), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n633), .A2(new_n409), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n603), .A2(new_n574), .A3(new_n578), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n527), .A2(new_n648), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n654), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n236), .ZN(G30));
  NAND2_X1  g479(.A1(new_n497), .A2(new_n498), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT38), .Z(new_n667));
  XOR2_X1   g481(.A(new_n659), .B(KEYINPUT39), .Z(new_n668));
  AND2_X1   g482(.A1(new_n310), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n601), .A2(new_n570), .ZN(new_n673));
  INV_X1    g487(.A(new_n556), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n190), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G472), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n574), .A2(new_n578), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n662), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n372), .A2(new_n409), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n420), .A3(new_n680), .ZN(new_n681));
  OR4_X1    g495(.A1(new_n667), .A2(new_n671), .A3(new_n672), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n270), .ZN(G45));
  INV_X1    g497(.A(new_n659), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n622), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n661), .A2(new_n662), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n499), .A3(new_n310), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n305), .B2(new_n306), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n303), .A2(new_n304), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n190), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n690), .A3(G469), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n191), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n532), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n661), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n623), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT41), .B(G113), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  INV_X1    g516(.A(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n639), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT103), .B(G116), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G18));
  NAND2_X1  g520(.A1(new_n499), .A2(new_n697), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n418), .A2(new_n661), .A3(new_n662), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n424), .ZN(G21));
  AND3_X1   g524(.A1(new_n666), .A2(new_n697), .A3(new_n420), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n601), .A2(KEYINPUT28), .ZN(new_n712));
  INV_X1    g526(.A(new_n587), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n570), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n577), .B1(new_n715), .B2(new_n560), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n610), .B2(new_n609), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n718), .B(G472), .C1(new_n576), .C2(G902), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n698), .ZN(new_n721));
  INV_X1    g535(.A(new_n680), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n416), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n711), .A2(new_n721), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n720), .A2(new_n698), .A3(new_n417), .A4(new_n680), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT105), .B1(new_n726), .B2(new_n707), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  INV_X1    g543(.A(new_n685), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n717), .A2(new_n719), .ZN(new_n732));
  INV_X1    g546(.A(new_n716), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n662), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n731), .B1(new_n720), .B2(new_n662), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n730), .B(new_n711), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n578), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(KEYINPUT109), .B(new_n739), .C1(new_n579), .C2(new_n738), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n738), .B1(new_n574), .B2(new_n578), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT108), .B1(new_n608), .B2(new_n575), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n744), .A3(new_n603), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n622), .A2(KEYINPUT42), .A3(new_n684), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n308), .B(KEYINPUT107), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n307), .B(new_n747), .C1(new_n306), .C2(new_n298), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n191), .A2(new_n493), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n497), .A2(new_n498), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n745), .A2(new_n698), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n497), .A2(new_n498), .A3(new_n748), .A4(new_n749), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n604), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n753), .B1(new_n755), .B2(new_n685), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  NAND3_X1  g572(.A1(new_n754), .A2(new_n604), .A3(new_n660), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n754), .A2(new_n604), .A3(new_n761), .A4(new_n660), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  NAND3_X1  g578(.A1(new_n497), .A2(new_n498), .A3(new_n420), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n621), .A2(new_n633), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT43), .B1(new_n766), .B2(KEYINPUT111), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n611), .A2(new_n662), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT112), .Z(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n765), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT45), .B1(new_n299), .B2(new_n301), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  OAI21_X1  g590(.A(G469), .B1(new_n298), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n747), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n307), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n191), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n668), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n769), .A2(new_n771), .A3(KEYINPUT44), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n774), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  NOR3_X1   g602(.A1(new_n685), .A2(new_n661), .A3(new_n698), .ZN(new_n789));
  INV_X1    g603(.A(new_n765), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(KEYINPUT113), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(KEYINPUT113), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n782), .A2(KEYINPUT47), .A3(new_n783), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT47), .B1(new_n782), .B2(new_n783), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n792), .B(new_n793), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  AND2_X1   g612(.A1(new_n697), .A2(new_n493), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n667), .A2(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n769), .A2(new_n413), .A3(new_n721), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n695), .A2(new_n696), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n497), .A3(new_n498), .A4(new_n749), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n767), .A2(new_n768), .A3(new_n808), .A4(new_n412), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n734), .B2(new_n735), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n678), .A2(new_n698), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n808), .A3(new_n412), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n372), .A3(new_n621), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n783), .B1(new_n695), .B2(new_n696), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n795), .A2(new_n796), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n802), .A2(new_n790), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT51), .B1(new_n806), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n745), .A2(new_n698), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n809), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n812), .A2(new_n622), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n802), .A2(new_n711), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n410), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n654), .A2(new_n663), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n490), .A2(new_n722), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n748), .A2(new_n783), .A3(new_n684), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n679), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n736), .A2(new_n827), .A3(new_n688), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n622), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n416), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n492), .A2(new_n835), .A3(new_n500), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT114), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n492), .A2(new_n835), .A3(new_n500), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n612), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n407), .A2(new_n402), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n372), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n416), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n492), .A2(new_n500), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n492), .A2(new_n500), .A3(new_n846), .A4(new_n843), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n612), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n650), .A2(new_n605), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n840), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n633), .A2(new_n841), .A3(new_n659), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n310), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n686), .A3(new_n765), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n732), .A2(new_n662), .A3(new_n733), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT106), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n720), .A2(new_n731), .A3(new_n662), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n685), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n858), .B2(new_n754), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n757), .A3(new_n763), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n623), .A2(new_n699), .B1(new_n707), .B2(new_n708), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n704), .A2(new_n728), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n833), .A2(new_n851), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n664), .B1(new_n858), .B2(new_n711), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT52), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n865), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n867), .A2(new_n832), .A3(new_n688), .A4(new_n830), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n752), .A2(new_n756), .B1(new_n760), .B2(new_n762), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n861), .B1(new_n725), .B2(new_n727), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n704), .A4(new_n859), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n873), .A2(new_n876), .A3(new_n850), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(KEYINPUT53), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n866), .B1(new_n868), .B2(KEYINPUT52), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n833), .A2(new_n851), .A3(new_n864), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n881), .B(new_n882), .C1(new_n877), .C2(KEYINPUT53), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n818), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n826), .A2(new_n879), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n811), .A2(new_n493), .A3(new_n766), .A4(new_n191), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n807), .B(KEYINPUT49), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n667), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n889), .ZN(G75));
  NAND2_X1  g704(.A1(new_n865), .A2(new_n866), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n190), .B1(new_n891), .B2(new_n881), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(G210), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n471), .B(KEYINPUT117), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n465), .ZN(new_n896));
  NOR2_X1   g710(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n192), .A2(G952), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G51));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n883), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n891), .A2(KEYINPUT119), .A3(new_n882), .A4(new_n881), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n881), .B1(new_n877), .B2(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n747), .B(KEYINPUT57), .Z(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n692), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n775), .A2(new_n777), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n892), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n900), .B1(new_n910), .B2(new_n912), .ZN(G54));
  AND2_X1   g727(.A1(KEYINPUT58), .A2(G475), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n905), .A2(G902), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n360), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n892), .A2(new_n369), .A3(new_n914), .ZN(new_n917));
  INV_X1    g731(.A(new_n900), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n916), .A2(new_n917), .A3(new_n921), .A4(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(G60));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n879), .B2(new_n883), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n614), .A2(new_n616), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n918), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n925), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n907), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G63));
  XNOR2_X1  g745(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n394), .A2(new_n190), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n905), .A2(new_n647), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n934), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n891), .B2(new_n881), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n935), .B(new_n918), .C1(new_n937), .C2(new_n522), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n938), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT61), .B1(new_n938), .B2(KEYINPUT121), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(G66));
  OAI21_X1  g755(.A(G953), .B1(new_n415), .B2(new_n460), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n850), .A2(new_n863), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT123), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n944), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n894), .B1(G898), .B2(new_n192), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  AND2_X1   g761(.A1(new_n797), .A2(new_n787), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n785), .A2(new_n820), .A3(new_n828), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n874), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n736), .A2(new_n827), .A3(new_n688), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n948), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n797), .A2(new_n787), .A3(new_n953), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT125), .B1(new_n955), .B2(new_n950), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n956), .A3(new_n192), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n583), .B(new_n353), .ZN(new_n958));
  NAND2_X1  g772(.A1(G900), .A2(G953), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n682), .A2(new_n953), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n834), .A2(new_n842), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n669), .A2(new_n790), .A3(new_n964), .A4(new_n604), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(KEYINPUT124), .A3(new_n948), .A4(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n961), .A2(new_n962), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT62), .B1(new_n682), .B2(new_n953), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n948), .B(new_n965), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n960), .B1(new_n972), .B2(new_n958), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT127), .Z(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n960), .B(new_n977), .C1(new_n972), .C2(new_n958), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(G72));
  NAND3_X1  g795(.A1(new_n966), .A2(new_n971), .A3(new_n944), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  AOI211_X1 g798(.A(new_n570), .B(new_n584), .C1(new_n982), .C2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n556), .B1(new_n584), .B2(new_n551), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n984), .B(new_n986), .C1(new_n870), .C2(new_n878), .ZN(new_n987));
  INV_X1    g801(.A(new_n984), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n954), .A2(new_n956), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n944), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n584), .A2(new_n570), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n987), .B(new_n918), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n985), .A2(new_n992), .ZN(G57));
endmodule


