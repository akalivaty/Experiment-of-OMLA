//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1196, new_n1197,
    new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT69), .Z(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n453), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT70), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(G112), .B2(new_n460), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT71), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n482));
  AOI22_X1  g057(.A1(G124), .A2(new_n482), .B1(new_n473), .B2(G136), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n481), .A2(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT72), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n485), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n463), .A2(new_n469), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n491), .A2(new_n493), .B1(new_n495), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  AND3_X1   g075(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT5), .B1(KEYINPUT73), .B2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n505), .A2(G651), .B1(G50), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n503), .B2(new_n508), .ZN(new_n514));
  OAI221_X1 g089(.A(KEYINPUT74), .B1(new_n506), .B2(new_n507), .C1(new_n501), .C2(new_n502), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n511), .B1(new_n512), .B2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT75), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT75), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT73), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n510), .A2(G51), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n514), .A2(new_n515), .A3(G89), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n523), .A2(new_n530), .A3(new_n531), .ZN(G168));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  INV_X1    g108(.A(G77), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n503), .A2(new_n533), .B1(new_n534), .B2(new_n509), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI221_X1 g112(.A(KEYINPUT76), .B1(new_n534), .B2(new_n509), .C1(new_n503), .C2(new_n533), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G651), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n510), .A2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n514), .A2(new_n515), .A3(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n503), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n546), .A2(G651), .B1(G43), .B2(new_n510), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n514), .A2(new_n515), .A3(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n510), .A2(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n510), .A2(new_n559), .A3(G53), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT78), .B(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n503), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n558), .A2(new_n560), .B1(G651), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n514), .A2(new_n515), .A3(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n542), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n541), .A2(new_n540), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n569), .A2(KEYINPUT79), .A3(new_n539), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G301));
  NAND3_X1  g147(.A1(new_n523), .A2(new_n531), .A3(new_n530), .ZN(G286));
  OR2_X1    g148(.A1(new_n528), .A2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G49), .B2(new_n510), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n514), .A2(new_n515), .A3(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  OAI21_X1  g152(.A(G61), .B1(new_n501), .B2(new_n502), .ZN(new_n578));
  AND3_X1   g153(.A1(KEYINPUT80), .A2(G73), .A3(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT80), .B1(G73), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n510), .B2(G48), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n514), .A2(new_n515), .A3(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n528), .A2(G60), .ZN(new_n586));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT81), .B1(new_n588), .B2(G651), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  INV_X1    g165(.A(G651), .ZN(new_n591));
  AOI211_X1 g166(.A(new_n590), .B(new_n591), .C1(new_n586), .C2(new_n587), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n510), .A2(G47), .ZN(new_n595));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n594), .B(new_n595), .C1(new_n516), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n595), .B1(new_n516), .B2(new_n596), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND3_X1  g177(.A1(new_n514), .A2(new_n515), .A3(G92), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT10), .Z(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n503), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n571), .B2(G868), .ZN(G284));
  XOR2_X1   g186(.A(G284), .B(KEYINPUT83), .Z(G321));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(G168), .A2(new_n614), .ZN(new_n615));
  AOI211_X1 g190(.A(new_n613), .B(new_n615), .C1(new_n614), .C2(G299), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n613), .B2(new_n615), .ZN(G297));
  AOI21_X1  g192(.A(new_n616), .B1(new_n613), .B2(new_n615), .ZN(G280));
  INV_X1    g193(.A(new_n609), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n549), .A2(new_n614), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n609), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g200(.A1(new_n463), .A2(new_n469), .A3(new_n474), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  AOI22_X1  g206(.A1(G123), .A2(new_n482), .B1(new_n473), .B2(G135), .ZN(new_n632));
  NOR3_X1   g207(.A1(new_n460), .A2(KEYINPUT85), .A3(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT85), .B1(new_n460), .B2(G111), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT86), .Z(G156));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT87), .ZN(G401));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT17), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT88), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n656), .A3(new_n658), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n657), .A2(new_n658), .ZN(new_n666));
  INV_X1    g241(.A(new_n656), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n660), .B1(new_n667), .B2(new_n659), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(new_n683), .B(new_n682), .S(new_n675), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n689), .B2(new_n693), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G6), .A2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G305), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G303), .B2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1971), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G23), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G288), .B2(new_n703), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT33), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n702), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT34), .Z(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT90), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n473), .A2(G131), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n482), .A2(G119), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n716), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT91), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n601), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G16), .B2(G24), .ZN(new_n727));
  INV_X1    g302(.A(G1986), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n713), .B(new_n729), .C1(new_n728), .C2(new_n727), .ZN(new_n730));
  NOR2_X1   g305(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n714), .A2(G35), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT98), .Z(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n714), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2090), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n703), .A2(G20), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT23), .Z(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G299), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT100), .Z(new_n745));
  NOR2_X1   g320(.A1(G4), .A2(G16), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT94), .Z(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n619), .B2(G16), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1348), .ZN(new_n749));
  NOR2_X1   g324(.A1(G171), .A2(new_n703), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G5), .B2(new_n703), .ZN(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G16), .A2(G19), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n550), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1341), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n751), .A2(new_n752), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n749), .A2(new_n753), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n703), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n703), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(G1966), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n714), .A2(G33), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n473), .A2(G139), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n463), .A2(new_n469), .A3(G127), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n460), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n762), .B1(new_n770), .B2(new_n714), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n761), .B1(G2072), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n714), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n714), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n772), .B1(G2072), .B2(new_n771), .C1(G2078), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n714), .A2(G32), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n473), .A2(G141), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT96), .Z(new_n778));
  AND2_X1   g353(.A1(new_n474), .A2(G105), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT26), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n779), .B(new_n781), .C1(G129), .C2(new_n482), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n776), .B1(new_n784), .B2(new_n714), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n714), .A2(KEYINPUT28), .A3(G26), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT28), .B1(new_n714), .B2(G26), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n473), .A2(G140), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n482), .A2(G128), .ZN(new_n791));
  OR2_X1    g366(.A1(G104), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n788), .B(new_n789), .C1(new_n794), .C2(G29), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT95), .B(G2067), .Z(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n795), .A2(new_n797), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT31), .B(G11), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT97), .B(G28), .Z(new_n801));
  AOI21_X1  g376(.A(G29), .B1(new_n801), .B2(KEYINPUT30), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(KEYINPUT30), .B2(new_n801), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n803), .C1(new_n636), .C2(new_n714), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n798), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT24), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n714), .B1(new_n806), .B2(G34), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n806), .B2(G34), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G160), .B2(G29), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G2084), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n760), .A2(G1966), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n787), .A2(new_n805), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n774), .A2(G2078), .ZN(new_n813));
  OAI221_X1 g388(.A(new_n813), .B1(G2084), .B2(new_n809), .C1(new_n738), .C2(G2090), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n775), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n745), .A2(new_n758), .A3(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT101), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(KEYINPUT101), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n732), .A2(new_n733), .B1(new_n817), .B2(new_n818), .ZN(G311));
  NAND2_X1  g394(.A1(new_n732), .A2(new_n733), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n818), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(G150));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n503), .B2(new_n824), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n825), .A2(G651), .B1(G55), .B2(new_n510), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n516), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G860), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT37), .Z(new_n830));
  NOR2_X1   g405(.A1(new_n609), .A2(new_n620), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT103), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n826), .B(KEYINPUT103), .C1(new_n827), .C2(new_n516), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n550), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n828), .A2(new_n834), .A3(new_n549), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n833), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  AOI21_X1  g416(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n843), .A2(KEYINPUT104), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(KEYINPUT104), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n830), .B1(new_n844), .B2(new_n845), .ZN(G145));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n847));
  INV_X1    g422(.A(new_n770), .ZN(new_n848));
  AOI22_X1  g423(.A1(G130), .A2(new_n482), .B1(new_n473), .B2(G142), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  INV_X1    g425(.A(G118), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n850), .A2(KEYINPUT105), .B1(new_n851), .B2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(KEYINPUT105), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT106), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(new_n627), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n627), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n783), .A2(new_n794), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n783), .A2(new_n794), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n721), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n721), .B1(new_n859), .B2(new_n860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n859), .A2(new_n860), .ZN(new_n865));
  INV_X1    g440(.A(new_n721), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n867), .A2(new_n857), .A3(new_n856), .A4(new_n861), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n498), .A2(new_n495), .ZN(new_n869));
  INV_X1    g444(.A(new_n490), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n864), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n864), .B2(new_n868), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n848), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n864), .A2(new_n868), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n490), .B1(new_n498), .B2(new_n495), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n770), .A3(new_n872), .ZN(new_n879));
  XOR2_X1   g454(.A(G160), .B(new_n636), .Z(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(G162), .Z(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n875), .B2(new_n879), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n847), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n875), .A2(new_n879), .ZN(new_n887));
  INV_X1    g462(.A(new_n881), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n889), .A2(KEYINPUT40), .A3(new_n883), .A4(new_n882), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n886), .A2(new_n890), .ZN(G395));
  NAND2_X1  g466(.A1(new_n609), .A2(G299), .ZN(new_n892));
  INV_X1    g467(.A(G299), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n604), .A3(new_n608), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(KEYINPUT41), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n619), .A2(new_n620), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n837), .A2(new_n838), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n623), .A2(KEYINPUT107), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n839), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n895), .A3(new_n905), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n699), .B1(new_n598), .B2(new_n600), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n915), .A2(new_n593), .A3(G305), .A4(new_n597), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G303), .B(G288), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n918), .A3(new_n916), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n908), .A2(new_n924), .A3(new_n911), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n913), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n913), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n828), .A2(new_n614), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(G295));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n929), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n914), .A2(new_n918), .A3(new_n916), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n918), .B1(new_n914), .B2(new_n916), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT109), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n920), .A2(new_n937), .A3(new_n921), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n568), .A2(G168), .A3(new_n570), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n941));
  NAND3_X1  g516(.A1(G171), .A2(new_n941), .A3(G286), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT108), .B1(G168), .B2(new_n542), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n903), .A2(new_n940), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n839), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n895), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n897), .A2(new_n944), .A3(new_n946), .A4(new_n898), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n939), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n933), .B1(new_n950), .B2(G37), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n897), .A2(new_n898), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n945), .B(new_n903), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT110), .B(new_n883), .C1(new_n954), .C2(new_n939), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n954), .B2(new_n922), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n948), .A2(new_n922), .A3(new_n949), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n883), .C1(new_n954), .C2(new_n939), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n932), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(new_n955), .A3(new_n958), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n950), .A2(G37), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n962), .A2(KEYINPUT43), .B1(new_n963), .B2(new_n956), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n961), .B1(new_n964), .B2(new_n932), .ZN(G397));
  XOR2_X1   g540(.A(KEYINPUT111), .B(G1384), .Z(new_n966));
  NAND2_X1  g541(.A1(new_n871), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n470), .A2(new_n471), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G2105), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(G40), .A3(new_n475), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT112), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n783), .B(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G2067), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n794), .B(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n721), .B(new_n723), .Z(new_n982));
  OAI21_X1  g557(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n601), .B(G1986), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n974), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT113), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  NOR3_X1   g563(.A1(G166), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n871), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT114), .B1(new_n877), .B2(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(G2090), .ZN(new_n997));
  INV_X1    g572(.A(G40), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n472), .A2(new_n476), .A3(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n485), .A2(new_n492), .A3(new_n489), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n492), .B1(new_n485), .B2(new_n489), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n869), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n993), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n996), .A2(new_n997), .A3(new_n999), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1971), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n871), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n999), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n1002), .B2(new_n993), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n991), .B1(new_n1011), .B2(new_n988), .ZN(new_n1012));
  INV_X1    g587(.A(G1966), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n994), .A2(new_n995), .A3(new_n968), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1002), .A2(new_n993), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n999), .B1(new_n1015), .B2(new_n968), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n992), .B1(new_n871), .B2(new_n993), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n877), .A2(KEYINPUT114), .A3(G1384), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1003), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n972), .B1(KEYINPUT50), .B2(new_n1015), .ZN(new_n1021));
  INV_X1    g596(.A(G2084), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n988), .B(G286), .C1(new_n1017), .C2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1021), .A3(new_n997), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n988), .B1(new_n1025), .B2(new_n1010), .ZN(new_n1026));
  INV_X1    g601(.A(new_n991), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n999), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n583), .A2(new_n584), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n583), .B2(new_n584), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G305), .A2(G1981), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n583), .A2(new_n584), .A3(new_n1031), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1029), .A2(new_n1034), .A3(new_n1037), .A4(G8), .ZN(new_n1038));
  INV_X1    g613(.A(G288), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G1976), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1029), .A2(G8), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n994), .A2(new_n995), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n988), .B1(new_n1046), .B2(new_n999), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1045), .B1(new_n1047), .B2(new_n1040), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1012), .A2(new_n1024), .A3(new_n1028), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT63), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n1051), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1029), .A2(G8), .A3(new_n1040), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1043), .B(new_n1038), .C1(new_n1056), .C2(new_n1045), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT115), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1028), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(new_n1051), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G164), .A2(G1384), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n999), .B1(new_n1062), .B2(new_n1003), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT50), .B1(new_n994), .B2(new_n995), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1063), .A2(new_n1064), .A3(G2084), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n972), .B1(new_n1062), .B2(KEYINPUT45), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n994), .A2(new_n995), .A3(new_n968), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1966), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1061), .A2(G286), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1058), .A2(new_n1060), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1054), .A2(new_n1055), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1038), .A2(new_n1041), .A3(new_n1039), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1036), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1047), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1074), .B2(KEYINPUT116), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1058), .A2(new_n1059), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1012), .A2(new_n1028), .A3(new_n1049), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1009), .ZN(new_n1080));
  INV_X1    g655(.A(G2078), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n999), .A4(new_n1007), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n752), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1083), .A2(G2078), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1066), .A2(new_n1067), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(new_n571), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n969), .A2(new_n999), .A3(new_n1007), .A4(new_n1086), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1084), .A2(new_n1085), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT124), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1084), .A2(new_n1085), .A3(new_n1095), .A4(new_n1092), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(G171), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1079), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G168), .A2(new_n988), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1069), .A2(KEYINPUT122), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n988), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1099), .B(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1100), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1101), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1099), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1088), .A2(new_n571), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1084), .A2(new_n1085), .A3(G301), .A4(new_n1092), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1115), .B2(new_n1090), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1098), .B(new_n1111), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1348), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1029), .B2(G2067), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1046), .A2(KEYINPUT118), .A3(new_n978), .A4(new_n999), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n619), .ZN(new_n1125));
  XNOR2_X1  g700(.A(G299), .B(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1004), .A2(new_n999), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(G1956), .B1(new_n1128), .B2(new_n996), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  AND4_X1   g705(.A1(new_n999), .A2(new_n1080), .A3(new_n1007), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1126), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  INV_X1    g709(.A(new_n996), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(new_n1127), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G299), .B(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1080), .A2(new_n999), .A3(new_n1007), .A4(new_n1130), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1133), .A2(new_n1140), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1132), .A2(new_n1140), .A3(KEYINPUT61), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT119), .B(G1996), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1008), .A2(new_n1009), .A3(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(G1341), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1046), .B2(new_n999), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n550), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT59), .B(new_n550), .C1(new_n1144), .C2(new_n1147), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1120), .A2(new_n1122), .A3(KEYINPUT60), .A4(new_n1123), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1150), .B(new_n1151), .C1(new_n1152), .C2(new_n619), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT61), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1142), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1124), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(new_n619), .A3(new_n1152), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1141), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1072), .B(new_n1078), .C1(new_n1118), .C2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1111), .B2(KEYINPUT62), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  AOI211_X1 g738(.A(KEYINPUT125), .B(new_n1163), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1109), .A2(new_n1163), .A3(new_n1110), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1079), .A2(new_n1113), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1162), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n986), .B1(new_n1160), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT46), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n784), .B(new_n979), .C1(new_n1170), .C2(G1996), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n975), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n974), .B2(G1996), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1173), .A2(KEYINPUT126), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(KEYINPUT126), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT47), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n974), .A2(G1986), .A3(G290), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1178), .A2(KEYINPUT48), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(KEYINPUT48), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(new_n983), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n980), .A2(new_n866), .A3(new_n723), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(G2067), .B2(new_n794), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n975), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1177), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1169), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g761(.A1(new_n654), .A2(G319), .A3(new_n672), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n1188), .B1(new_n695), .B2(new_n696), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1190));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n1188), .B(new_n1191), .C1(new_n695), .C2(new_n696), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1193), .B1(new_n884), .B2(new_n885), .ZN(new_n1194));
  NOR2_X1   g768(.A1(new_n1194), .A2(new_n964), .ZN(G308));
  NAND2_X1  g769(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n963), .A2(new_n956), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g772(.A1(new_n889), .A2(new_n883), .A3(new_n882), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n1198), .A2(new_n1199), .A3(new_n1193), .ZN(G225));
endmodule


